VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO output_terminal
  CLASS BLOCK ;
  FOREIGN output_terminal ;
  ORIGIN 6.000 6.000 ;
  SIZE 774.000 BY 771.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 756.300 771.300 758.700 ;
        RECT 762.300 686.700 771.300 756.300 ;
        RECT 0.600 684.300 771.300 686.700 ;
        RECT 762.300 614.700 771.300 684.300 ;
        RECT 0.600 612.300 771.300 614.700 ;
        RECT 762.300 542.700 771.300 612.300 ;
        RECT 0.600 540.300 771.300 542.700 ;
        RECT 762.300 470.700 771.300 540.300 ;
        RECT 0.600 468.300 771.300 470.700 ;
        RECT 762.300 398.700 771.300 468.300 ;
        RECT 0.600 396.300 771.300 398.700 ;
        RECT 762.300 326.700 771.300 396.300 ;
        RECT 0.600 324.300 771.300 326.700 ;
        RECT 762.300 254.700 771.300 324.300 ;
        RECT 0.600 252.300 771.300 254.700 ;
        RECT 762.300 182.700 771.300 252.300 ;
        RECT 0.600 180.300 771.300 182.700 ;
        RECT 762.300 110.700 771.300 180.300 ;
        RECT 0.600 108.300 771.300 110.700 ;
        RECT 762.300 38.700 771.300 108.300 ;
        RECT 0.600 36.300 771.300 38.700 ;
        RECT 762.300 0.300 771.300 36.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.300 722.700 -0.300 758.700 ;
        RECT -9.300 720.300 761.400 722.700 ;
        RECT -9.300 650.700 -0.300 720.300 ;
        RECT -9.300 648.300 761.400 650.700 ;
        RECT -9.300 578.700 -0.300 648.300 ;
        RECT -9.300 576.300 761.400 578.700 ;
        RECT -9.300 506.700 -0.300 576.300 ;
        RECT -9.300 504.300 761.400 506.700 ;
        RECT -9.300 434.700 -0.300 504.300 ;
        RECT -9.300 432.300 761.400 434.700 ;
        RECT -9.300 362.700 -0.300 432.300 ;
        RECT -9.300 360.300 761.400 362.700 ;
        RECT -9.300 290.700 -0.300 360.300 ;
        RECT -9.300 288.300 761.400 290.700 ;
        RECT -9.300 218.700 -0.300 288.300 ;
        RECT -9.300 216.300 761.400 218.700 ;
        RECT -9.300 146.700 -0.300 216.300 ;
        RECT -9.300 144.300 761.400 146.700 ;
        RECT -9.300 74.700 -0.300 144.300 ;
        RECT -9.300 72.300 761.400 74.700 ;
        RECT -9.300 2.700 -0.300 72.300 ;
        RECT -9.300 0.300 761.400 2.700 ;
    END
  END vdd
  PIN Dout[11]
    PORT
      LAYER metal2 ;
        RECT 662.400 757.050 663.450 765.450 ;
        RECT 661.950 754.950 664.050 757.050 ;
        RECT 676.950 754.950 679.050 757.050 ;
        RECT 677.400 745.050 678.450 754.950 ;
        RECT 676.950 742.950 679.050 745.050 ;
      LAYER metal3 ;
        RECT 661.950 756.600 664.050 757.050 ;
        RECT 676.950 756.600 679.050 757.050 ;
        RECT 661.950 755.400 679.050 756.600 ;
        RECT 661.950 754.950 664.050 755.400 ;
        RECT 676.950 754.950 679.050 755.400 ;
    END
  END Dout[11]
  PIN Dout[10]
    PORT
      LAYER metal2 ;
        RECT 671.400 699.450 672.450 765.450 ;
        RECT 673.950 699.450 676.050 700.050 ;
        RECT 671.400 698.400 676.050 699.450 ;
        RECT 673.950 697.950 676.050 698.400 ;
    END
  END Dout[10]
  PIN Dout[9]
    PORT
      LAYER metal2 ;
        RECT 707.400 757.050 708.450 765.450 ;
        RECT 706.950 754.950 709.050 757.050 ;
        RECT 721.950 754.950 724.050 757.050 ;
        RECT 722.400 745.050 723.450 754.950 ;
        RECT 721.950 742.950 724.050 745.050 ;
      LAYER metal3 ;
        RECT 706.950 756.600 709.050 757.050 ;
        RECT 721.950 756.600 724.050 757.050 ;
        RECT 706.950 755.400 724.050 756.600 ;
        RECT 706.950 754.950 709.050 755.400 ;
        RECT 721.950 754.950 724.050 755.400 ;
    END
  END Dout[9]
  PIN Dout[8]
    PORT
      LAYER metal2 ;
        RECT 713.400 699.450 714.450 765.450 ;
        RECT 715.950 699.450 718.050 700.050 ;
        RECT 713.400 698.400 718.050 699.450 ;
        RECT 715.950 697.950 718.050 698.400 ;
    END
  END Dout[8]
  PIN Dout[7]
    PORT
      LAYER metal2 ;
        RECT 755.400 709.050 756.450 765.450 ;
        RECT 754.950 706.950 757.050 709.050 ;
        RECT 754.950 697.950 757.050 700.050 ;
        RECT 755.400 673.050 756.450 697.950 ;
        RECT 754.950 670.950 757.050 673.050 ;
      LAYER metal3 ;
        RECT 754.950 706.950 757.050 709.050 ;
        RECT 755.400 700.050 756.600 706.950 ;
        RECT 754.950 697.950 757.050 700.050 ;
    END
  END Dout[7]
  PIN Dout[6]
    PORT
      LAYER metal2 ;
        RECT 748.950 625.950 751.050 628.050 ;
      LAYER metal3 ;
        RECT 748.950 627.600 751.050 628.050 ;
        RECT 767.400 627.600 768.600 630.600 ;
        RECT 748.950 626.400 768.600 627.600 ;
        RECT 748.950 625.950 751.050 626.400 ;
    END
  END Dout[6]
  PIN Dout[5]
    PORT
      LAYER metal2 ;
        RECT 727.950 600.450 730.050 601.050 ;
        RECT 727.950 599.400 732.450 600.450 ;
        RECT 727.950 598.950 730.050 599.400 ;
        RECT 731.400 595.050 732.450 599.400 ;
        RECT 730.950 592.950 733.050 595.050 ;
      LAYER metal3 ;
        RECT 730.950 594.600 733.050 595.050 ;
        RECT 730.950 593.400 768.600 594.600 ;
        RECT 730.950 592.950 733.050 593.400 ;
    END
  END Dout[5]
  PIN Dout[4]
    PORT
      LAYER metal2 ;
        RECT 748.950 553.950 751.050 556.050 ;
      LAYER metal3 ;
        RECT 748.950 555.600 751.050 556.050 ;
        RECT 767.400 555.600 768.600 558.600 ;
        RECT 748.950 554.400 768.600 555.600 ;
        RECT 748.950 553.950 751.050 554.400 ;
    END
  END Dout[4]
  PIN Dout[3]
    PORT
      LAYER metal2 ;
        RECT 748.950 528.450 751.050 529.050 ;
        RECT 746.400 527.400 751.050 528.450 ;
        RECT 746.400 523.050 747.450 527.400 ;
        RECT 748.950 526.950 751.050 527.400 ;
        RECT 745.950 520.950 748.050 523.050 ;
      LAYER metal3 ;
        RECT 745.950 522.600 748.050 523.050 ;
        RECT 745.950 521.400 768.600 522.600 ;
        RECT 745.950 520.950 748.050 521.400 ;
    END
  END Dout[3]
  PIN Dout[2]
    PORT
      LAYER metal2 ;
        RECT 706.950 493.950 709.050 496.050 ;
        RECT 703.950 483.450 706.050 484.050 ;
        RECT 707.400 483.450 708.450 493.950 ;
        RECT 703.950 482.400 708.450 483.450 ;
        RECT 703.950 481.950 706.050 482.400 ;
      LAYER metal3 ;
        RECT 706.950 495.600 709.050 496.050 ;
        RECT 706.950 494.400 768.600 495.600 ;
        RECT 706.950 493.950 709.050 494.400 ;
    END
  END Dout[2]
  PIN Dout[1]
    PORT
      LAYER metal2 ;
        RECT 736.950 487.950 739.050 490.050 ;
        RECT 733.950 411.450 736.050 412.050 ;
        RECT 737.400 411.450 738.450 487.950 ;
        RECT 733.950 410.400 738.450 411.450 ;
        RECT 733.950 409.950 736.050 410.400 ;
      LAYER metal3 ;
        RECT 736.950 489.600 739.050 490.050 ;
        RECT 736.950 488.400 768.600 489.600 ;
        RECT 736.950 487.950 739.050 488.400 ;
    END
  END Dout[1]
  PIN Dout[0]
    PORT
      LAYER metal2 ;
        RECT 745.950 481.950 748.050 484.050 ;
      LAYER metal3 ;
        RECT 745.950 483.600 748.050 484.050 ;
        RECT 745.950 482.400 768.600 483.600 ;
        RECT 745.950 481.950 748.050 482.400 ;
    END
  END Dout[0]
  PIN ISin
    PORT
      LAYER metal2 ;
        RECT 28.950 736.950 31.050 739.050 ;
      LAYER metal3 ;
        RECT 28.950 738.600 31.050 739.050 ;
        RECT -3.600 737.400 31.050 738.600 ;
        RECT 28.950 736.950 31.050 737.400 ;
    END
  END ISin
  PIN Rdy
    PORT
      LAYER metal2 ;
        RECT 10.950 457.950 13.050 460.050 ;
        RECT 11.400 339.450 12.450 457.950 ;
        RECT 13.950 339.450 16.050 340.050 ;
        RECT 11.400 338.400 16.050 339.450 ;
        RECT 13.950 337.950 16.050 338.400 ;
      LAYER metal3 ;
        RECT 10.950 459.600 13.050 460.050 ;
        RECT -3.600 458.400 13.050 459.600 ;
        RECT 10.950 457.950 13.050 458.400 ;
    END
  END Rdy
  PIN Vld
    PORT
      LAYER metal2 ;
        RECT 521.400 764.400 525.450 765.450 ;
        RECT 524.400 745.050 525.450 764.400 ;
        RECT 523.950 742.950 526.050 745.050 ;
    END
  END Vld
  PIN Xin[1]
    PORT
      LAYER metal2 ;
        RECT 478.950 99.450 481.050 100.050 ;
        RECT 476.400 98.400 481.050 99.450 ;
        RECT 476.400 88.050 477.450 98.400 ;
        RECT 478.950 97.950 481.050 98.400 ;
        RECT 601.950 88.950 604.050 91.050 ;
        RECT 602.400 88.050 603.450 88.950 ;
        RECT 475.950 85.950 478.050 88.050 ;
        RECT 601.950 85.950 604.050 88.050 ;
        RECT 469.950 16.950 472.050 19.050 ;
        RECT 470.400 13.050 471.450 16.950 ;
        RECT 476.400 13.050 477.450 85.950 ;
        RECT 556.950 16.950 559.050 19.050 ;
        RECT 557.400 13.050 558.450 16.950 ;
        RECT 454.950 10.950 457.050 13.050 ;
        RECT 469.950 10.950 472.050 13.050 ;
        RECT 475.950 10.950 478.050 13.050 ;
        RECT 556.950 10.950 559.050 13.050 ;
        RECT 455.400 -3.600 456.450 10.950 ;
      LAYER metal3 ;
        RECT 475.950 87.600 478.050 88.050 ;
        RECT 601.950 87.600 604.050 88.050 ;
        RECT 475.950 86.400 604.050 87.600 ;
        RECT 475.950 85.950 478.050 86.400 ;
        RECT 601.950 85.950 604.050 86.400 ;
        RECT 454.950 12.600 457.050 13.050 ;
        RECT 469.950 12.600 472.050 13.050 ;
        RECT 475.950 12.600 478.050 13.050 ;
        RECT 556.950 12.600 559.050 13.050 ;
        RECT 454.950 11.400 559.050 12.600 ;
        RECT 454.950 10.950 457.050 11.400 ;
        RECT 469.950 10.950 472.050 11.400 ;
        RECT 475.950 10.950 478.050 11.400 ;
        RECT 556.950 10.950 559.050 11.400 ;
    END
  END Xin[1]
  PIN Xin[0]
    PORT
      LAYER metal2 ;
        RECT 193.950 169.950 196.050 172.050 ;
        RECT 220.950 169.950 223.050 172.050 ;
        RECT 221.400 16.050 222.450 169.950 ;
        RECT 535.950 160.950 538.050 163.050 ;
        RECT 265.950 16.950 268.050 19.050 ;
        RECT 385.950 16.950 388.050 19.050 ;
        RECT 266.400 16.050 267.450 16.950 ;
        RECT 386.400 16.050 387.450 16.950 ;
        RECT 536.400 16.050 537.450 160.950 ;
        RECT 220.950 13.950 223.050 16.050 ;
        RECT 265.950 13.950 268.050 16.050 ;
        RECT 385.950 13.950 388.050 16.050 ;
        RECT 460.950 13.950 463.050 16.050 ;
        RECT 535.950 13.950 538.050 16.050 ;
        RECT 461.400 -3.600 462.450 13.950 ;
      LAYER metal3 ;
        RECT 193.950 171.600 196.050 172.050 ;
        RECT 220.950 171.600 223.050 172.050 ;
        RECT 193.950 170.400 223.050 171.600 ;
        RECT 193.950 169.950 196.050 170.400 ;
        RECT 220.950 169.950 223.050 170.400 ;
        RECT 220.950 15.600 223.050 16.050 ;
        RECT 265.950 15.600 268.050 16.050 ;
        RECT 385.950 15.600 388.050 16.050 ;
        RECT 460.950 15.600 463.050 16.050 ;
        RECT 535.950 15.600 538.050 16.050 ;
        RECT 220.950 14.400 538.050 15.600 ;
        RECT 220.950 13.950 223.050 14.400 ;
        RECT 265.950 13.950 268.050 14.400 ;
        RECT 385.950 13.950 388.050 14.400 ;
        RECT 460.950 13.950 463.050 14.400 ;
        RECT 535.950 13.950 538.050 14.400 ;
    END
  END Xin[0]
  PIN Yin[1]
    PORT
      LAYER metal2 ;
        RECT 250.950 448.950 253.050 451.050 ;
        RECT 251.400 445.050 252.450 448.950 ;
        RECT 124.950 442.950 127.050 445.050 ;
        RECT 250.950 442.950 253.050 445.050 ;
        RECT 265.950 442.950 268.050 445.050 ;
        RECT 125.400 388.050 126.450 442.950 ;
        RECT 124.950 385.950 127.050 388.050 ;
        RECT 266.400 277.050 267.450 442.950 ;
        RECT 265.950 274.950 268.050 277.050 ;
        RECT 328.950 274.950 331.050 277.050 ;
        RECT 391.950 274.950 394.050 277.050 ;
        RECT 329.400 274.050 330.450 274.950 ;
        RECT 328.950 271.950 331.050 274.050 ;
        RECT 392.400 61.050 393.450 274.950 ;
        RECT 391.950 58.950 394.050 61.050 ;
        RECT 532.950 58.950 535.050 61.050 ;
        RECT 556.950 58.950 559.050 61.050 ;
        RECT 533.400 -3.600 534.450 58.950 ;
        RECT 557.400 58.050 558.450 58.950 ;
        RECT 556.950 55.950 559.050 58.050 ;
      LAYER metal3 ;
        RECT 124.950 444.600 127.050 445.050 ;
        RECT 250.950 444.600 253.050 445.050 ;
        RECT 265.950 444.600 268.050 445.050 ;
        RECT 124.950 443.400 268.050 444.600 ;
        RECT 124.950 442.950 127.050 443.400 ;
        RECT 250.950 442.950 253.050 443.400 ;
        RECT 265.950 442.950 268.050 443.400 ;
        RECT 265.950 276.600 268.050 277.050 ;
        RECT 328.950 276.600 331.050 277.050 ;
        RECT 391.950 276.600 394.050 277.050 ;
        RECT 265.950 275.400 394.050 276.600 ;
        RECT 265.950 274.950 268.050 275.400 ;
        RECT 328.950 274.950 331.050 275.400 ;
        RECT 391.950 274.950 394.050 275.400 ;
        RECT 391.950 60.600 394.050 61.050 ;
        RECT 532.950 60.600 535.050 61.050 ;
        RECT 556.950 60.600 559.050 61.050 ;
        RECT 391.950 59.400 559.050 60.600 ;
        RECT 391.950 58.950 394.050 59.400 ;
        RECT 532.950 58.950 535.050 59.400 ;
        RECT 556.950 58.950 559.050 59.400 ;
    END
  END Yin[1]
  PIN Yin[0]
    PORT
      LAYER metal2 ;
        RECT 97.950 459.450 100.050 460.050 ;
        RECT 97.950 458.400 102.450 459.450 ;
        RECT 97.950 457.950 100.050 458.400 ;
        RECT 101.400 451.050 102.450 458.400 ;
        RECT 100.950 448.950 103.050 451.050 ;
        RECT 136.950 448.950 139.050 451.050 ;
        RECT 412.950 448.950 415.050 451.050 ;
        RECT 137.400 442.050 138.450 448.950 ;
        RECT 413.400 442.050 414.450 448.950 ;
        RECT 136.950 439.950 139.050 442.050 ;
        RECT 412.950 439.950 415.050 442.050 ;
        RECT 532.950 439.950 535.050 442.050 ;
        RECT 529.950 306.450 532.050 307.050 ;
        RECT 533.400 306.450 534.450 439.950 ;
        RECT 529.950 305.400 534.450 306.450 ;
        RECT 529.950 304.950 532.050 305.400 ;
        RECT 530.400 276.450 531.450 304.950 ;
        RECT 527.400 275.400 531.450 276.450 ;
        RECT 527.400 7.050 528.450 275.400 ;
        RECT 526.950 4.950 529.050 7.050 ;
        RECT 538.950 4.950 541.050 7.050 ;
        RECT 539.400 -3.600 540.450 4.950 ;
      LAYER metal3 ;
        RECT 100.950 450.600 103.050 451.050 ;
        RECT 136.950 450.600 139.050 451.050 ;
        RECT 100.950 449.400 139.050 450.600 ;
        RECT 100.950 448.950 103.050 449.400 ;
        RECT 136.950 448.950 139.050 449.400 ;
        RECT 136.950 441.600 139.050 442.050 ;
        RECT 412.950 441.600 415.050 442.050 ;
        RECT 532.950 441.600 535.050 442.050 ;
        RECT 136.950 440.400 535.050 441.600 ;
        RECT 136.950 439.950 139.050 440.400 ;
        RECT 412.950 439.950 415.050 440.400 ;
        RECT 532.950 439.950 535.050 440.400 ;
        RECT 526.950 6.600 529.050 7.050 ;
        RECT 538.950 6.600 541.050 7.050 ;
        RECT 526.950 5.400 541.050 6.600 ;
        RECT 526.950 4.950 529.050 5.400 ;
        RECT 538.950 4.950 541.050 5.400 ;
    END
  END Yin[0]
  PIN clk
    PORT
      LAYER metal2 ;
        RECT 583.950 523.950 586.050 526.050 ;
        RECT 584.400 520.050 585.450 523.950 ;
        RECT 562.950 517.950 565.050 520.050 ;
        RECT 583.950 517.950 586.050 520.050 ;
        RECT 563.400 499.050 564.450 517.950 ;
        RECT 37.950 496.950 40.050 499.050 ;
        RECT 394.950 496.950 397.050 499.050 ;
        RECT 562.950 496.950 565.050 499.050 ;
        RECT 34.950 453.450 37.050 454.050 ;
        RECT 38.400 453.450 39.450 496.950 ;
        RECT 395.400 487.050 396.450 496.950 ;
        RECT 394.950 484.950 397.050 487.050 ;
        RECT 34.950 452.400 39.450 453.450 ;
        RECT 34.950 451.950 37.050 452.400 ;
        RECT 38.400 406.050 39.450 452.400 ;
        RECT 37.950 403.950 40.050 406.050 ;
        RECT 55.950 403.950 58.050 406.050 ;
        RECT 56.400 199.050 57.450 403.950 ;
        RECT 563.400 400.050 564.450 496.950 ;
        RECT 562.950 397.950 565.050 400.050 ;
        RECT 568.950 397.950 571.050 400.050 ;
        RECT 569.400 343.050 570.450 397.950 ;
        RECT 568.950 340.950 571.050 343.050 ;
        RECT 616.950 340.950 619.050 343.050 ;
        RECT 55.950 196.950 58.050 199.050 ;
        RECT 91.950 196.950 94.050 199.050 ;
        RECT 92.400 127.050 93.450 196.950 ;
        RECT 91.950 124.950 94.050 127.050 ;
        RECT 617.400 94.050 618.450 340.950 ;
        RECT 616.950 91.950 619.050 94.050 ;
        RECT 643.950 91.950 646.050 94.050 ;
      LAYER metal3 ;
        RECT 562.950 519.600 565.050 520.050 ;
        RECT 583.950 519.600 586.050 520.050 ;
        RECT 562.950 518.400 586.050 519.600 ;
        RECT 562.950 517.950 565.050 518.400 ;
        RECT 583.950 517.950 586.050 518.400 ;
        RECT 37.950 498.600 40.050 499.050 ;
        RECT 394.950 498.600 397.050 499.050 ;
        RECT 562.950 498.600 565.050 499.050 ;
        RECT 37.950 497.400 565.050 498.600 ;
        RECT 37.950 496.950 40.050 497.400 ;
        RECT 394.950 496.950 397.050 497.400 ;
        RECT 562.950 496.950 565.050 497.400 ;
        RECT 34.950 453.600 37.050 454.050 ;
        RECT -3.600 452.400 37.050 453.600 ;
        RECT 34.950 451.950 37.050 452.400 ;
        RECT 37.950 405.600 40.050 406.050 ;
        RECT 55.950 405.600 58.050 406.050 ;
        RECT 37.950 404.400 58.050 405.600 ;
        RECT 37.950 403.950 40.050 404.400 ;
        RECT 55.950 403.950 58.050 404.400 ;
        RECT 562.950 399.600 565.050 400.050 ;
        RECT 568.950 399.600 571.050 400.050 ;
        RECT 562.950 398.400 571.050 399.600 ;
        RECT 562.950 397.950 565.050 398.400 ;
        RECT 568.950 397.950 571.050 398.400 ;
        RECT 568.950 342.600 571.050 343.050 ;
        RECT 616.950 342.600 619.050 343.050 ;
        RECT 568.950 341.400 619.050 342.600 ;
        RECT 568.950 340.950 571.050 341.400 ;
        RECT 616.950 340.950 619.050 341.400 ;
        RECT 55.950 198.600 58.050 199.050 ;
        RECT 91.950 198.600 94.050 199.050 ;
        RECT 55.950 197.400 94.050 198.600 ;
        RECT 55.950 196.950 58.050 197.400 ;
        RECT 91.950 196.950 94.050 197.400 ;
        RECT 616.950 93.600 619.050 94.050 ;
        RECT 643.950 93.600 646.050 94.050 ;
        RECT 616.950 92.400 646.050 93.600 ;
        RECT 616.950 91.950 619.050 92.400 ;
        RECT 643.950 91.950 646.050 92.400 ;
    END
  END clk
  PIN selSign
    PORT
      LAYER metal2 ;
        RECT 748.950 88.950 751.050 91.050 ;
        RECT 749.400 48.450 750.450 88.950 ;
        RECT 751.950 48.450 754.050 49.050 ;
        RECT 749.400 47.400 754.050 48.450 ;
        RECT 751.950 46.950 754.050 47.400 ;
        RECT 752.400 37.050 753.450 46.950 ;
        RECT 742.950 34.950 745.050 37.050 ;
        RECT 751.950 34.950 754.050 37.050 ;
        RECT 743.400 4.050 744.450 34.950 ;
        RECT 748.950 16.950 751.050 19.050 ;
        RECT 749.400 4.050 750.450 16.950 ;
        RECT 742.950 1.950 745.050 4.050 ;
        RECT 748.950 1.950 751.050 4.050 ;
        RECT 743.400 -3.600 744.450 1.950 ;
      LAYER metal3 ;
        RECT 742.950 36.600 745.050 37.050 ;
        RECT 751.950 36.600 754.050 37.050 ;
        RECT 742.950 35.400 754.050 36.600 ;
        RECT 742.950 34.950 745.050 35.400 ;
        RECT 751.950 34.950 754.050 35.400 ;
        RECT 742.950 3.600 745.050 4.050 ;
        RECT 748.950 3.600 751.050 4.050 ;
        RECT 742.950 2.400 751.050 3.600 ;
        RECT 742.950 1.950 745.050 2.400 ;
        RECT 748.950 1.950 751.050 2.400 ;
    END
  END selSign
  PIN selXY
    PORT
      LAYER metal2 ;
        RECT 691.950 625.950 694.050 628.050 ;
        RECT 700.950 625.950 703.050 628.050 ;
        RECT 688.950 600.450 691.050 601.050 ;
        RECT 692.400 600.450 693.450 625.950 ;
        RECT 688.950 599.400 693.450 600.450 ;
        RECT 688.950 598.950 691.050 599.400 ;
        RECT 692.400 556.050 693.450 599.400 ;
        RECT 691.950 553.950 694.050 556.050 ;
        RECT 694.950 553.950 697.050 556.050 ;
        RECT 700.950 553.950 703.050 556.050 ;
        RECT 691.950 411.450 694.050 412.050 ;
        RECT 695.400 411.450 696.450 553.950 ;
        RECT 691.950 410.400 696.450 411.450 ;
        RECT 691.950 409.950 694.050 410.400 ;
        RECT 695.400 387.450 696.450 410.400 ;
        RECT 695.400 386.400 699.450 387.450 ;
        RECT 698.400 276.450 699.450 386.400 ;
        RECT 695.400 275.400 699.450 276.450 ;
        RECT 695.400 -3.600 696.450 275.400 ;
      LAYER metal3 ;
        RECT 691.950 627.600 694.050 628.050 ;
        RECT 700.950 627.600 703.050 628.050 ;
        RECT 691.950 626.400 703.050 627.600 ;
        RECT 691.950 625.950 694.050 626.400 ;
        RECT 700.950 625.950 703.050 626.400 ;
        RECT 691.950 555.600 694.050 556.050 ;
        RECT 694.950 555.600 697.050 556.050 ;
        RECT 700.950 555.600 703.050 556.050 ;
        RECT 691.950 554.400 703.050 555.600 ;
        RECT 691.950 553.950 694.050 554.400 ;
        RECT 694.950 553.950 697.050 554.400 ;
        RECT 700.950 553.950 703.050 554.400 ;
    END
  END selXY
  OBS
      LAYER metal1 ;
        RECT 29.850 749.400 31.650 755.250 ;
        RECT 34.350 748.200 36.150 755.250 ;
        RECT 73.650 749.400 75.450 755.250 ;
        RECT 32.550 747.300 36.150 748.200 ;
        RECT 74.250 747.300 75.450 749.400 ;
        RECT 76.650 750.300 78.450 755.250 ;
        RECT 79.650 751.200 81.450 755.250 ;
        RECT 82.650 750.300 84.450 755.250 ;
        RECT 76.650 748.950 84.450 750.300 ;
        RECT 87.150 749.400 88.950 755.250 ;
        RECT 90.150 752.400 91.950 755.250 ;
        RECT 94.950 753.300 96.750 755.250 ;
        RECT 93.000 752.400 96.750 753.300 ;
        RECT 99.450 752.400 101.250 755.250 ;
        RECT 102.750 752.400 104.550 755.250 ;
        RECT 106.650 752.400 108.450 755.250 ;
        RECT 110.850 752.400 112.650 755.250 ;
        RECT 115.350 752.400 117.150 755.250 ;
        RECT 93.000 751.500 94.050 752.400 ;
        RECT 91.950 749.400 94.050 751.500 ;
        RECT 102.750 750.600 103.800 752.400 ;
        RECT 29.100 741.150 30.900 742.950 ;
        RECT 28.950 739.050 31.050 741.150 ;
        RECT 32.550 739.950 33.750 747.300 ;
        RECT 74.250 746.250 78.000 747.300 ;
        RECT 76.950 742.950 78.150 746.250 ;
        RECT 80.100 744.150 81.900 745.950 ;
        RECT 35.100 741.150 36.900 742.950 ;
        RECT 31.950 737.850 34.050 739.950 ;
        RECT 34.950 739.050 37.050 741.150 ;
        RECT 76.950 740.850 79.050 742.950 ;
        RECT 79.950 742.050 82.050 744.150 ;
        RECT 82.950 740.850 85.050 742.950 ;
        RECT 73.950 737.850 76.050 739.950 ;
        RECT 32.550 729.600 33.750 737.850 ;
        RECT 74.250 736.050 76.050 737.850 ;
        RECT 77.850 735.600 79.050 740.850 ;
        RECT 83.100 739.050 84.900 740.850 ;
        RECT 87.150 736.800 88.050 749.400 ;
        RECT 95.550 748.800 97.350 750.600 ;
        RECT 98.850 749.550 103.800 750.600 ;
        RECT 111.300 751.500 112.350 752.400 ;
        RECT 111.300 750.300 115.050 751.500 ;
        RECT 98.850 748.800 100.650 749.550 ;
        RECT 95.850 747.900 96.900 748.800 ;
        RECT 106.050 748.200 107.850 750.000 ;
        RECT 112.950 749.400 115.050 750.300 ;
        RECT 118.650 749.400 120.450 755.250 ;
        RECT 151.650 749.400 153.450 755.250 ;
        RECT 106.050 747.900 106.950 748.200 ;
        RECT 95.850 747.000 106.950 747.900 ;
        RECT 119.250 747.150 120.450 749.400 ;
        RECT 95.850 745.800 96.900 747.000 ;
        RECT 90.000 744.600 96.900 745.800 ;
        RECT 90.000 743.850 90.900 744.600 ;
        RECT 95.100 744.000 96.900 744.600 ;
        RECT 89.100 742.050 90.900 743.850 ;
        RECT 92.100 742.950 93.900 743.700 ;
        RECT 106.050 742.950 106.950 747.000 ;
        RECT 115.950 745.050 120.450 747.150 ;
        RECT 152.250 747.300 153.450 749.400 ;
        RECT 154.650 750.300 156.450 755.250 ;
        RECT 157.650 751.200 159.450 755.250 ;
        RECT 160.650 750.300 162.450 755.250 ;
        RECT 154.650 748.950 162.450 750.300 ;
        RECT 165.150 749.400 166.950 755.250 ;
        RECT 168.150 752.400 169.950 755.250 ;
        RECT 172.950 753.300 174.750 755.250 ;
        RECT 171.000 752.400 174.750 753.300 ;
        RECT 177.450 752.400 179.250 755.250 ;
        RECT 180.750 752.400 182.550 755.250 ;
        RECT 184.650 752.400 186.450 755.250 ;
        RECT 188.850 752.400 190.650 755.250 ;
        RECT 193.350 752.400 195.150 755.250 ;
        RECT 171.000 751.500 172.050 752.400 ;
        RECT 169.950 749.400 172.050 751.500 ;
        RECT 180.750 750.600 181.800 752.400 ;
        RECT 152.250 746.250 156.000 747.300 ;
        RECT 114.150 743.250 118.050 745.050 ;
        RECT 115.950 742.950 118.050 743.250 ;
        RECT 92.100 741.900 100.050 742.950 ;
        RECT 97.950 740.850 100.050 741.900 ;
        RECT 103.950 740.850 106.950 742.950 ;
        RECT 96.450 737.100 98.250 737.400 ;
        RECT 96.450 736.800 104.850 737.100 ;
        RECT 87.150 736.200 104.850 736.800 ;
        RECT 87.150 735.600 98.250 736.200 ;
        RECT 29.550 723.750 31.350 729.600 ;
        RECT 32.550 723.750 34.350 729.600 ;
        RECT 35.550 723.750 37.350 729.600 ;
        RECT 74.400 723.750 76.200 729.600 ;
        RECT 77.700 723.750 79.500 735.600 ;
        RECT 81.900 723.750 83.700 735.600 ;
        RECT 87.150 723.750 88.950 735.600 ;
        RECT 101.250 734.700 103.050 735.300 ;
        RECT 95.550 733.500 103.050 734.700 ;
        RECT 103.950 734.100 104.850 736.200 ;
        RECT 106.050 736.200 106.950 740.850 ;
        RECT 116.250 737.400 118.050 739.200 ;
        RECT 112.950 736.200 117.150 737.400 ;
        RECT 106.050 735.300 112.050 736.200 ;
        RECT 112.950 735.300 115.050 736.200 ;
        RECT 119.250 735.600 120.450 745.050 ;
        RECT 154.950 742.950 156.150 746.250 ;
        RECT 158.100 744.150 159.900 745.950 ;
        RECT 154.950 740.850 157.050 742.950 ;
        RECT 157.950 742.050 160.050 744.150 ;
        RECT 160.950 740.850 163.050 742.950 ;
        RECT 151.950 737.850 154.050 739.950 ;
        RECT 152.250 736.050 154.050 737.850 ;
        RECT 155.850 735.600 157.050 740.850 ;
        RECT 161.100 739.050 162.900 740.850 ;
        RECT 165.150 736.800 166.050 749.400 ;
        RECT 173.550 748.800 175.350 750.600 ;
        RECT 176.850 749.550 181.800 750.600 ;
        RECT 189.300 751.500 190.350 752.400 ;
        RECT 189.300 750.300 193.050 751.500 ;
        RECT 176.850 748.800 178.650 749.550 ;
        RECT 173.850 747.900 174.900 748.800 ;
        RECT 184.050 748.200 185.850 750.000 ;
        RECT 190.950 749.400 193.050 750.300 ;
        RECT 196.650 749.400 198.450 755.250 ;
        RECT 230.550 752.400 232.350 755.250 ;
        RECT 233.550 752.400 235.350 755.250 ;
        RECT 269.550 752.400 271.350 755.250 ;
        RECT 272.550 752.400 274.350 755.250 ;
        RECT 275.550 752.400 277.350 755.250 ;
        RECT 184.050 747.900 184.950 748.200 ;
        RECT 173.850 747.000 184.950 747.900 ;
        RECT 197.250 747.150 198.450 749.400 ;
        RECT 173.850 745.800 174.900 747.000 ;
        RECT 168.000 744.600 174.900 745.800 ;
        RECT 168.000 743.850 168.900 744.600 ;
        RECT 173.100 744.000 174.900 744.600 ;
        RECT 167.100 742.050 168.900 743.850 ;
        RECT 170.100 742.950 171.900 743.700 ;
        RECT 184.050 742.950 184.950 747.000 ;
        RECT 193.950 745.050 198.450 747.150 ;
        RECT 192.150 743.250 196.050 745.050 ;
        RECT 193.950 742.950 196.050 743.250 ;
        RECT 170.100 741.900 178.050 742.950 ;
        RECT 175.950 740.850 178.050 741.900 ;
        RECT 181.950 740.850 184.950 742.950 ;
        RECT 174.450 737.100 176.250 737.400 ;
        RECT 174.450 736.800 182.850 737.100 ;
        RECT 165.150 736.200 182.850 736.800 ;
        RECT 165.150 735.600 176.250 736.200 ;
        RECT 111.150 734.400 112.050 735.300 ;
        RECT 108.450 734.100 110.250 734.400 ;
        RECT 95.550 732.600 96.750 733.500 ;
        RECT 103.950 733.200 110.250 734.100 ;
        RECT 108.450 732.600 110.250 733.200 ;
        RECT 111.150 732.600 113.850 734.400 ;
        RECT 91.950 730.500 96.750 732.600 ;
        RECT 99.150 730.500 106.050 732.300 ;
        RECT 95.550 729.600 96.750 730.500 ;
        RECT 90.150 723.750 91.950 729.600 ;
        RECT 95.250 723.750 97.050 729.600 ;
        RECT 100.050 723.750 101.850 729.600 ;
        RECT 103.050 723.750 104.850 730.500 ;
        RECT 111.150 729.600 115.050 731.700 ;
        RECT 106.950 723.750 108.750 729.600 ;
        RECT 111.150 723.750 112.950 729.600 ;
        RECT 115.650 723.750 117.450 726.600 ;
        RECT 118.650 723.750 120.450 735.600 ;
        RECT 152.400 723.750 154.200 729.600 ;
        RECT 155.700 723.750 157.500 735.600 ;
        RECT 159.900 723.750 161.700 735.600 ;
        RECT 165.150 723.750 166.950 735.600 ;
        RECT 179.250 734.700 181.050 735.300 ;
        RECT 173.550 733.500 181.050 734.700 ;
        RECT 181.950 734.100 182.850 736.200 ;
        RECT 184.050 736.200 184.950 740.850 ;
        RECT 194.250 737.400 196.050 739.200 ;
        RECT 190.950 736.200 195.150 737.400 ;
        RECT 184.050 735.300 190.050 736.200 ;
        RECT 190.950 735.300 193.050 736.200 ;
        RECT 197.250 735.600 198.450 745.050 ;
        RECT 229.950 743.850 232.050 745.950 ;
        RECT 233.400 744.150 234.600 752.400 ;
        RECT 273.450 748.200 274.350 752.400 ;
        RECT 278.550 749.400 280.350 755.250 ;
        RECT 314.850 749.400 316.650 755.250 ;
        RECT 273.450 747.300 276.750 748.200 ;
        RECT 274.950 746.400 276.750 747.300 ;
        RECT 230.100 742.050 231.900 743.850 ;
        RECT 232.950 742.050 235.050 744.150 ;
        RECT 268.950 743.850 271.050 745.950 ;
        RECT 269.100 742.050 270.900 743.850 ;
        RECT 189.150 734.400 190.050 735.300 ;
        RECT 186.450 734.100 188.250 734.400 ;
        RECT 173.550 732.600 174.750 733.500 ;
        RECT 181.950 733.200 188.250 734.100 ;
        RECT 186.450 732.600 188.250 733.200 ;
        RECT 189.150 732.600 191.850 734.400 ;
        RECT 169.950 730.500 174.750 732.600 ;
        RECT 177.150 730.500 184.050 732.300 ;
        RECT 173.550 729.600 174.750 730.500 ;
        RECT 168.150 723.750 169.950 729.600 ;
        RECT 173.250 723.750 175.050 729.600 ;
        RECT 178.050 723.750 179.850 729.600 ;
        RECT 181.050 723.750 182.850 730.500 ;
        RECT 189.150 729.600 193.050 731.700 ;
        RECT 184.950 723.750 186.750 729.600 ;
        RECT 189.150 723.750 190.950 729.600 ;
        RECT 193.650 723.750 195.450 726.600 ;
        RECT 196.650 723.750 198.450 735.600 ;
        RECT 233.400 729.600 234.600 742.050 ;
        RECT 271.950 740.850 274.050 742.950 ;
        RECT 272.100 739.050 273.900 740.850 ;
        RECT 275.700 738.150 276.600 746.400 ;
        RECT 279.000 744.150 280.050 749.400 ;
        RECT 319.350 748.200 321.150 755.250 ;
        RECT 356.850 749.400 358.650 755.250 ;
        RECT 361.350 748.200 363.150 755.250 ;
        RECT 398.550 750.300 400.350 755.250 ;
        RECT 401.550 751.200 403.350 755.250 ;
        RECT 404.550 750.300 406.350 755.250 ;
        RECT 398.550 748.950 406.350 750.300 ;
        RECT 407.550 749.400 409.350 755.250 ;
        RECT 440.850 749.400 442.650 755.250 ;
        RECT 277.950 742.050 280.050 744.150 ;
        RECT 317.550 747.300 321.150 748.200 ;
        RECT 359.550 747.300 363.150 748.200 ;
        RECT 407.550 747.300 408.750 749.400 ;
        RECT 445.350 748.200 447.150 755.250 ;
        RECT 274.950 738.000 276.750 738.150 ;
        RECT 269.550 736.800 276.750 738.000 ;
        RECT 269.550 735.600 270.750 736.800 ;
        RECT 274.950 736.350 276.750 736.800 ;
        RECT 230.550 723.750 232.350 729.600 ;
        RECT 233.550 723.750 235.350 729.600 ;
        RECT 269.550 723.750 271.350 735.600 ;
        RECT 278.100 735.450 279.450 742.050 ;
        RECT 314.100 741.150 315.900 742.950 ;
        RECT 313.950 739.050 316.050 741.150 ;
        RECT 317.550 739.950 318.750 747.300 ;
        RECT 320.100 741.150 321.900 742.950 ;
        RECT 356.100 741.150 357.900 742.950 ;
        RECT 316.950 737.850 319.050 739.950 ;
        RECT 319.950 739.050 322.050 741.150 ;
        RECT 355.950 739.050 358.050 741.150 ;
        RECT 359.550 739.950 360.750 747.300 ;
        RECT 405.000 746.250 408.750 747.300 ;
        RECT 443.550 747.300 447.150 748.200 ;
        RECT 453.150 749.400 454.950 755.250 ;
        RECT 456.150 752.400 457.950 755.250 ;
        RECT 460.950 753.300 462.750 755.250 ;
        RECT 459.000 752.400 462.750 753.300 ;
        RECT 465.450 752.400 467.250 755.250 ;
        RECT 468.750 752.400 470.550 755.250 ;
        RECT 472.650 752.400 474.450 755.250 ;
        RECT 476.850 752.400 478.650 755.250 ;
        RECT 481.350 752.400 483.150 755.250 ;
        RECT 459.000 751.500 460.050 752.400 ;
        RECT 457.950 749.400 460.050 751.500 ;
        RECT 468.750 750.600 469.800 752.400 ;
        RECT 401.100 744.150 402.900 745.950 ;
        RECT 362.100 741.150 363.900 742.950 ;
        RECT 358.950 737.850 361.050 739.950 ;
        RECT 361.950 739.050 364.050 741.150 ;
        RECT 397.950 740.850 400.050 742.950 ;
        RECT 400.950 742.050 403.050 744.150 ;
        RECT 404.850 742.950 406.050 746.250 ;
        RECT 403.950 740.850 406.050 742.950 ;
        RECT 440.100 741.150 441.900 742.950 ;
        RECT 398.100 739.050 399.900 740.850 ;
        RECT 274.050 723.750 275.850 735.450 ;
        RECT 277.050 734.100 279.450 735.450 ;
        RECT 277.050 723.750 278.850 734.100 ;
        RECT 317.550 729.600 318.750 737.850 ;
        RECT 359.550 729.600 360.750 737.850 ;
        RECT 403.950 735.600 405.150 740.850 ;
        RECT 406.950 737.850 409.050 739.950 ;
        RECT 439.950 739.050 442.050 741.150 ;
        RECT 443.550 739.950 444.750 747.300 ;
        RECT 446.100 741.150 447.900 742.950 ;
        RECT 442.950 737.850 445.050 739.950 ;
        RECT 445.950 739.050 448.050 741.150 ;
        RECT 406.950 736.050 408.750 737.850 ;
        RECT 314.550 723.750 316.350 729.600 ;
        RECT 317.550 723.750 319.350 729.600 ;
        RECT 320.550 723.750 322.350 729.600 ;
        RECT 356.550 723.750 358.350 729.600 ;
        RECT 359.550 723.750 361.350 729.600 ;
        RECT 362.550 723.750 364.350 729.600 ;
        RECT 399.300 723.750 401.100 735.600 ;
        RECT 403.500 723.750 405.300 735.600 ;
        RECT 443.550 729.600 444.750 737.850 ;
        RECT 453.150 736.800 454.050 749.400 ;
        RECT 461.550 748.800 463.350 750.600 ;
        RECT 464.850 749.550 469.800 750.600 ;
        RECT 477.300 751.500 478.350 752.400 ;
        RECT 477.300 750.300 481.050 751.500 ;
        RECT 464.850 748.800 466.650 749.550 ;
        RECT 461.850 747.900 462.900 748.800 ;
        RECT 472.050 748.200 473.850 750.000 ;
        RECT 478.950 749.400 481.050 750.300 ;
        RECT 484.650 749.400 486.450 755.250 ;
        RECT 518.550 752.400 520.350 755.250 ;
        RECT 472.050 747.900 472.950 748.200 ;
        RECT 461.850 747.000 472.950 747.900 ;
        RECT 485.250 747.150 486.450 749.400 ;
        RECT 519.150 748.500 520.350 752.400 ;
        RECT 521.850 749.400 523.650 755.250 ;
        RECT 524.850 749.400 526.650 755.250 ;
        RECT 531.150 749.400 532.950 755.250 ;
        RECT 534.150 752.400 535.950 755.250 ;
        RECT 538.950 753.300 540.750 755.250 ;
        RECT 537.000 752.400 540.750 753.300 ;
        RECT 543.450 752.400 545.250 755.250 ;
        RECT 546.750 752.400 548.550 755.250 ;
        RECT 550.650 752.400 552.450 755.250 ;
        RECT 554.850 752.400 556.650 755.250 ;
        RECT 559.350 752.400 561.150 755.250 ;
        RECT 537.000 751.500 538.050 752.400 ;
        RECT 535.950 749.400 538.050 751.500 ;
        RECT 546.750 750.600 547.800 752.400 ;
        RECT 519.150 747.600 524.250 748.500 ;
        RECT 461.850 745.800 462.900 747.000 ;
        RECT 456.000 744.600 462.900 745.800 ;
        RECT 456.000 743.850 456.900 744.600 ;
        RECT 461.100 744.000 462.900 744.600 ;
        RECT 455.100 742.050 456.900 743.850 ;
        RECT 458.100 742.950 459.900 743.700 ;
        RECT 472.050 742.950 472.950 747.000 ;
        RECT 481.950 745.050 486.450 747.150 ;
        RECT 480.150 743.250 484.050 745.050 ;
        RECT 481.950 742.950 484.050 743.250 ;
        RECT 458.100 741.900 466.050 742.950 ;
        RECT 463.950 740.850 466.050 741.900 ;
        RECT 469.950 740.850 472.950 742.950 ;
        RECT 462.450 737.100 464.250 737.400 ;
        RECT 462.450 736.800 470.850 737.100 ;
        RECT 453.150 736.200 470.850 736.800 ;
        RECT 453.150 735.600 464.250 736.200 ;
        RECT 406.800 723.750 408.600 729.600 ;
        RECT 440.550 723.750 442.350 729.600 ;
        RECT 443.550 723.750 445.350 729.600 ;
        RECT 446.550 723.750 448.350 729.600 ;
        RECT 453.150 723.750 454.950 735.600 ;
        RECT 467.250 734.700 469.050 735.300 ;
        RECT 461.550 733.500 469.050 734.700 ;
        RECT 469.950 734.100 470.850 736.200 ;
        RECT 472.050 736.200 472.950 740.850 ;
        RECT 482.250 737.400 484.050 739.200 ;
        RECT 478.950 736.200 483.150 737.400 ;
        RECT 472.050 735.300 478.050 736.200 ;
        RECT 478.950 735.300 481.050 736.200 ;
        RECT 485.250 735.600 486.450 745.050 ;
        RECT 522.000 746.700 524.250 747.600 ;
        RECT 517.950 740.850 520.050 742.950 ;
        RECT 518.100 739.050 519.900 740.850 ;
        RECT 522.000 738.300 523.050 746.700 ;
        RECT 525.150 742.950 526.350 749.400 ;
        RECT 523.950 740.850 526.350 742.950 ;
        RECT 522.000 737.400 524.250 738.300 ;
        RECT 477.150 734.400 478.050 735.300 ;
        RECT 474.450 734.100 476.250 734.400 ;
        RECT 461.550 732.600 462.750 733.500 ;
        RECT 469.950 733.200 476.250 734.100 ;
        RECT 474.450 732.600 476.250 733.200 ;
        RECT 477.150 732.600 479.850 734.400 ;
        RECT 457.950 730.500 462.750 732.600 ;
        RECT 465.150 730.500 472.050 732.300 ;
        RECT 461.550 729.600 462.750 730.500 ;
        RECT 456.150 723.750 457.950 729.600 ;
        RECT 461.250 723.750 463.050 729.600 ;
        RECT 466.050 723.750 467.850 729.600 ;
        RECT 469.050 723.750 470.850 730.500 ;
        RECT 477.150 729.600 481.050 731.700 ;
        RECT 472.950 723.750 474.750 729.600 ;
        RECT 477.150 723.750 478.950 729.600 ;
        RECT 481.650 723.750 483.450 726.600 ;
        RECT 484.650 723.750 486.450 735.600 ;
        RECT 518.550 736.500 524.250 737.400 ;
        RECT 518.550 729.600 519.750 736.500 ;
        RECT 525.150 735.600 526.350 740.850 ;
        RECT 531.150 736.800 532.050 749.400 ;
        RECT 539.550 748.800 541.350 750.600 ;
        RECT 542.850 749.550 547.800 750.600 ;
        RECT 555.300 751.500 556.350 752.400 ;
        RECT 555.300 750.300 559.050 751.500 ;
        RECT 542.850 748.800 544.650 749.550 ;
        RECT 539.850 747.900 540.900 748.800 ;
        RECT 550.050 748.200 551.850 750.000 ;
        RECT 556.950 749.400 559.050 750.300 ;
        RECT 562.650 749.400 564.450 755.250 ;
        RECT 596.550 752.400 598.350 755.250 ;
        RECT 599.550 752.400 601.350 755.250 ;
        RECT 635.550 752.400 637.350 755.250 ;
        RECT 638.550 752.400 640.350 755.250 ;
        RECT 550.050 747.900 550.950 748.200 ;
        RECT 539.850 747.000 550.950 747.900 ;
        RECT 563.250 747.150 564.450 749.400 ;
        RECT 539.850 745.800 540.900 747.000 ;
        RECT 534.000 744.600 540.900 745.800 ;
        RECT 534.000 743.850 534.900 744.600 ;
        RECT 539.100 744.000 540.900 744.600 ;
        RECT 533.100 742.050 534.900 743.850 ;
        RECT 536.100 742.950 537.900 743.700 ;
        RECT 550.050 742.950 550.950 747.000 ;
        RECT 559.950 745.050 564.450 747.150 ;
        RECT 558.150 743.250 562.050 745.050 ;
        RECT 559.950 742.950 562.050 743.250 ;
        RECT 536.100 741.900 544.050 742.950 ;
        RECT 541.950 740.850 544.050 741.900 ;
        RECT 547.950 740.850 550.950 742.950 ;
        RECT 540.450 737.100 542.250 737.400 ;
        RECT 540.450 736.800 548.850 737.100 ;
        RECT 531.150 736.200 548.850 736.800 ;
        RECT 531.150 735.600 542.250 736.200 ;
        RECT 518.550 723.750 520.350 729.600 ;
        RECT 521.850 723.750 523.650 735.600 ;
        RECT 524.850 723.750 526.650 735.600 ;
        RECT 531.150 723.750 532.950 735.600 ;
        RECT 545.250 734.700 547.050 735.300 ;
        RECT 539.550 733.500 547.050 734.700 ;
        RECT 547.950 734.100 548.850 736.200 ;
        RECT 550.050 736.200 550.950 740.850 ;
        RECT 560.250 737.400 562.050 739.200 ;
        RECT 556.950 736.200 561.150 737.400 ;
        RECT 550.050 735.300 556.050 736.200 ;
        RECT 556.950 735.300 559.050 736.200 ;
        RECT 563.250 735.600 564.450 745.050 ;
        RECT 595.950 743.850 598.050 745.950 ;
        RECT 599.400 744.150 600.600 752.400 ;
        RECT 596.100 742.050 597.900 743.850 ;
        RECT 598.950 742.050 601.050 744.150 ;
        RECT 634.950 743.850 637.050 745.950 ;
        RECT 638.400 744.150 639.600 752.400 ;
        RECT 676.350 749.400 678.150 755.250 ;
        RECT 679.350 749.400 681.150 755.250 ;
        RECT 682.650 752.400 684.450 755.250 ;
        RECT 716.550 752.400 718.350 755.250 ;
        RECT 635.100 742.050 636.900 743.850 ;
        RECT 637.950 742.050 640.050 744.150 ;
        RECT 676.650 742.950 677.850 749.400 ;
        RECT 682.650 748.500 683.850 752.400 ;
        RECT 678.750 747.600 683.850 748.500 ;
        RECT 717.150 748.500 718.350 752.400 ;
        RECT 719.850 749.400 721.650 755.250 ;
        RECT 722.850 749.400 724.650 755.250 ;
        RECT 717.150 747.600 722.250 748.500 ;
        RECT 678.750 746.700 681.000 747.600 ;
        RECT 555.150 734.400 556.050 735.300 ;
        RECT 552.450 734.100 554.250 734.400 ;
        RECT 539.550 732.600 540.750 733.500 ;
        RECT 547.950 733.200 554.250 734.100 ;
        RECT 552.450 732.600 554.250 733.200 ;
        RECT 555.150 732.600 557.850 734.400 ;
        RECT 535.950 730.500 540.750 732.600 ;
        RECT 543.150 730.500 550.050 732.300 ;
        RECT 539.550 729.600 540.750 730.500 ;
        RECT 534.150 723.750 535.950 729.600 ;
        RECT 539.250 723.750 541.050 729.600 ;
        RECT 544.050 723.750 545.850 729.600 ;
        RECT 547.050 723.750 548.850 730.500 ;
        RECT 555.150 729.600 559.050 731.700 ;
        RECT 550.950 723.750 552.750 729.600 ;
        RECT 555.150 723.750 556.950 729.600 ;
        RECT 559.650 723.750 561.450 726.600 ;
        RECT 562.650 723.750 564.450 735.600 ;
        RECT 599.400 729.600 600.600 742.050 ;
        RECT 638.400 729.600 639.600 742.050 ;
        RECT 676.650 740.850 679.050 742.950 ;
        RECT 676.650 735.600 677.850 740.850 ;
        RECT 679.950 738.300 681.000 746.700 ;
        RECT 720.000 746.700 722.250 747.600 ;
        RECT 682.950 740.850 685.050 742.950 ;
        RECT 715.950 740.850 718.050 742.950 ;
        RECT 683.100 739.050 684.900 740.850 ;
        RECT 716.100 739.050 717.900 740.850 ;
        RECT 678.750 737.400 681.000 738.300 ;
        RECT 720.000 738.300 721.050 746.700 ;
        RECT 723.150 742.950 724.350 749.400 ;
        RECT 721.950 740.850 724.350 742.950 ;
        RECT 720.000 737.400 722.250 738.300 ;
        RECT 678.750 736.500 684.450 737.400 ;
        RECT 596.550 723.750 598.350 729.600 ;
        RECT 599.550 723.750 601.350 729.600 ;
        RECT 635.550 723.750 637.350 729.600 ;
        RECT 638.550 723.750 640.350 729.600 ;
        RECT 676.350 723.750 678.150 735.600 ;
        RECT 679.350 723.750 681.150 735.600 ;
        RECT 683.250 729.600 684.450 736.500 ;
        RECT 682.650 723.750 684.450 729.600 ;
        RECT 716.550 736.500 722.250 737.400 ;
        RECT 716.550 729.600 717.750 736.500 ;
        RECT 723.150 735.600 724.350 740.850 ;
        RECT 716.550 723.750 718.350 729.600 ;
        RECT 719.850 723.750 721.650 735.600 ;
        RECT 722.850 723.750 724.650 735.600 ;
        RECT 34.650 707.400 36.450 719.250 ;
        RECT 37.650 707.400 39.450 719.250 ;
        RECT 40.650 707.400 42.450 719.250 ;
        RECT 76.650 713.400 78.450 719.250 ;
        RECT 79.650 714.000 81.450 719.250 ;
        RECT 77.250 713.100 78.450 713.400 ;
        RECT 82.650 713.400 84.450 719.250 ;
        RECT 85.650 713.400 87.450 719.250 ;
        RECT 119.550 713.400 121.350 719.250 ;
        RECT 122.550 713.400 124.350 719.250 ;
        RECT 125.550 714.000 127.350 719.250 ;
        RECT 82.650 713.100 84.300 713.400 ;
        RECT 77.250 712.200 84.300 713.100 ;
        RECT 122.700 713.100 124.350 713.400 ;
        RECT 128.550 713.400 130.350 719.250 ;
        RECT 128.550 713.100 129.750 713.400 ;
        RECT 122.700 712.200 129.750 713.100 ;
        RECT 37.800 700.950 39.150 707.400 ;
        RECT 77.250 703.950 78.300 712.200 ;
        RECT 83.100 708.150 84.900 709.950 ;
        RECT 122.100 708.150 123.900 709.950 ;
        RECT 79.950 705.150 81.750 706.950 ;
        RECT 82.950 706.050 85.050 708.150 ;
        RECT 86.100 705.150 87.900 706.950 ;
        RECT 119.100 705.150 120.900 706.950 ;
        RECT 121.950 706.050 124.050 708.150 ;
        RECT 125.250 705.150 127.050 706.950 ;
        RECT 76.950 701.850 79.050 703.950 ;
        RECT 79.950 703.050 82.050 705.150 ;
        RECT 85.950 703.050 88.050 705.150 ;
        RECT 118.950 703.050 121.050 705.150 ;
        RECT 124.950 703.050 127.050 705.150 ;
        RECT 128.700 703.950 129.750 712.200 ;
        RECT 166.350 707.400 168.150 719.250 ;
        RECT 169.350 707.400 171.150 719.250 ;
        RECT 172.650 713.400 174.450 719.250 ;
        RECT 208.650 713.400 210.450 719.250 ;
        RECT 211.650 713.400 213.450 719.250 ;
        RECT 245.550 713.400 247.350 719.250 ;
        RECT 248.550 713.400 250.350 719.250 ;
        RECT 287.400 713.400 289.200 719.250 ;
        RECT 127.950 701.850 130.050 703.950 ;
        RECT 166.650 702.150 167.850 707.400 ;
        RECT 173.250 706.500 174.450 713.400 ;
        RECT 168.750 705.600 174.450 706.500 ;
        RECT 168.750 704.700 171.000 705.600 ;
        RECT 34.950 698.850 39.150 700.950 ;
        RECT 40.950 698.850 43.050 700.950 ;
        RECT 37.800 693.600 39.150 698.850 ;
        RECT 41.100 697.050 42.900 698.850 ;
        RECT 77.400 697.650 78.600 701.850 ;
        RECT 128.400 697.650 129.600 701.850 ;
        RECT 77.400 696.000 81.900 697.650 ;
        RECT 34.650 687.750 36.450 693.600 ;
        RECT 37.650 687.750 39.450 693.600 ;
        RECT 40.650 687.750 42.450 693.600 ;
        RECT 80.100 687.750 81.900 696.000 ;
        RECT 85.500 687.750 87.300 696.600 ;
        RECT 119.700 687.750 121.500 696.600 ;
        RECT 125.100 696.000 129.600 697.650 ;
        RECT 166.650 700.050 169.050 702.150 ;
        RECT 125.100 687.750 126.900 696.000 ;
        RECT 166.650 693.600 167.850 700.050 ;
        RECT 169.950 696.300 171.000 704.700 ;
        RECT 173.100 702.150 174.900 703.950 ;
        RECT 172.950 700.050 175.050 702.150 ;
        RECT 209.400 700.950 210.600 713.400 ;
        RECT 248.400 700.950 249.600 713.400 ;
        RECT 290.700 707.400 292.500 719.250 ;
        RECT 294.900 707.400 296.700 719.250 ;
        RECT 326.550 707.400 328.350 719.250 ;
        RECT 331.050 707.550 332.850 719.250 ;
        RECT 334.050 708.900 335.850 719.250 ;
        RECT 334.050 707.550 336.450 708.900 ;
        RECT 287.250 705.150 289.050 706.950 ;
        RECT 286.950 703.050 289.050 705.150 ;
        RECT 290.850 702.150 292.050 707.400 ;
        RECT 326.550 706.200 327.750 707.400 ;
        RECT 331.950 706.200 333.750 706.650 ;
        RECT 326.550 705.000 333.750 706.200 ;
        RECT 331.950 704.850 333.750 705.000 ;
        RECT 296.100 702.150 297.900 703.950 ;
        RECT 329.100 702.150 330.900 703.950 ;
        RECT 208.950 698.850 211.050 700.950 ;
        RECT 212.100 699.150 213.900 700.950 ;
        RECT 245.100 699.150 246.900 700.950 ;
        RECT 168.750 695.400 171.000 696.300 ;
        RECT 168.750 694.500 173.850 695.400 ;
        RECT 166.350 687.750 168.150 693.600 ;
        RECT 169.350 687.750 171.150 693.600 ;
        RECT 172.650 690.600 173.850 694.500 ;
        RECT 209.400 690.600 210.600 698.850 ;
        RECT 211.950 697.050 214.050 699.150 ;
        RECT 244.950 697.050 247.050 699.150 ;
        RECT 247.950 698.850 250.050 700.950 ;
        RECT 289.950 700.050 292.050 702.150 ;
        RECT 248.400 690.600 249.600 698.850 ;
        RECT 289.950 696.750 291.150 700.050 ;
        RECT 292.950 698.850 295.050 700.950 ;
        RECT 295.950 700.050 298.050 702.150 ;
        RECT 326.100 699.150 327.900 700.950 ;
        RECT 328.950 700.050 331.050 702.150 ;
        RECT 293.100 697.050 294.900 698.850 ;
        RECT 325.950 697.050 328.050 699.150 ;
        RECT 287.250 695.700 291.000 696.750 ;
        RECT 332.700 696.600 333.600 704.850 ;
        RECT 335.100 700.950 336.450 707.550 ;
        RECT 371.550 708.300 373.350 719.250 ;
        RECT 374.550 709.200 376.350 719.250 ;
        RECT 377.550 708.300 379.350 719.250 ;
        RECT 371.550 707.400 379.350 708.300 ;
        RECT 380.550 707.400 382.350 719.250 ;
        RECT 418.650 718.500 426.450 719.250 ;
        RECT 418.650 707.400 420.450 718.500 ;
        RECT 421.650 707.400 423.450 717.600 ;
        RECT 424.650 708.600 426.450 718.500 ;
        RECT 427.650 709.500 429.450 719.250 ;
        RECT 430.650 708.600 432.450 719.250 ;
        RECT 424.650 707.700 432.450 708.600 ;
        RECT 435.150 707.400 436.950 719.250 ;
        RECT 438.150 713.400 439.950 719.250 ;
        RECT 443.250 713.400 445.050 719.250 ;
        RECT 448.050 713.400 449.850 719.250 ;
        RECT 443.550 712.500 444.750 713.400 ;
        RECT 451.050 712.500 452.850 719.250 ;
        RECT 454.950 713.400 456.750 719.250 ;
        RECT 459.150 713.400 460.950 719.250 ;
        RECT 463.650 716.400 465.450 719.250 ;
        RECT 439.950 710.400 444.750 712.500 ;
        RECT 447.150 710.700 454.050 712.500 ;
        RECT 459.150 711.300 463.050 713.400 ;
        RECT 443.550 709.500 444.750 710.400 ;
        RECT 456.450 709.800 458.250 710.400 ;
        RECT 443.550 708.300 451.050 709.500 ;
        RECT 449.250 707.700 451.050 708.300 ;
        RECT 451.950 708.900 458.250 709.800 ;
        RECT 380.700 702.150 381.900 707.400 ;
        RECT 421.800 706.500 423.600 707.400 ;
        RECT 435.150 706.800 446.250 707.400 ;
        RECT 451.950 706.800 452.850 708.900 ;
        RECT 456.450 708.600 458.250 708.900 ;
        RECT 459.150 708.600 461.850 710.400 ;
        RECT 459.150 707.700 460.050 708.600 ;
        RECT 421.800 705.600 425.850 706.500 ;
        RECT 419.100 702.150 420.900 703.950 ;
        RECT 424.950 702.150 425.850 705.600 ;
        RECT 435.150 706.200 452.850 706.800 ;
        RECT 430.950 702.150 432.750 703.950 ;
        RECT 334.950 698.850 337.050 700.950 ;
        RECT 370.950 698.850 373.050 700.950 ;
        RECT 374.100 699.150 375.900 700.950 ;
        RECT 331.950 695.700 333.750 696.600 ;
        RECT 287.250 693.600 288.450 695.700 ;
        RECT 330.450 694.800 333.750 695.700 ;
        RECT 172.650 687.750 174.450 690.600 ;
        RECT 208.650 687.750 210.450 690.600 ;
        RECT 211.650 687.750 213.450 690.600 ;
        RECT 245.550 687.750 247.350 690.600 ;
        RECT 248.550 687.750 250.350 690.600 ;
        RECT 286.650 687.750 288.450 693.600 ;
        RECT 289.650 692.700 297.450 694.050 ;
        RECT 289.650 687.750 291.450 692.700 ;
        RECT 292.650 687.750 294.450 691.800 ;
        RECT 295.650 687.750 297.450 692.700 ;
        RECT 330.450 690.600 331.350 694.800 ;
        RECT 336.000 693.600 337.050 698.850 ;
        RECT 371.100 697.050 372.900 698.850 ;
        RECT 373.950 697.050 376.050 699.150 ;
        RECT 376.950 698.850 379.050 700.950 ;
        RECT 379.950 700.050 382.050 702.150 ;
        RECT 418.950 700.050 421.050 702.150 ;
        RECT 377.100 697.050 378.900 698.850 ;
        RECT 380.700 693.600 381.900 700.050 ;
        RECT 421.950 698.850 424.050 700.950 ;
        RECT 424.950 700.050 427.050 702.150 ;
        RECT 422.250 697.050 424.050 698.850 ;
        RECT 426.000 693.600 427.050 700.050 ;
        RECT 427.950 698.850 430.050 700.950 ;
        RECT 430.950 700.050 433.050 702.150 ;
        RECT 427.950 697.050 429.750 698.850 ;
        RECT 435.150 693.600 436.050 706.200 ;
        RECT 444.450 705.900 452.850 706.200 ;
        RECT 454.050 706.800 460.050 707.700 ;
        RECT 460.950 706.800 463.050 707.700 ;
        RECT 466.650 707.400 468.450 719.250 ;
        RECT 500.550 713.400 502.350 719.250 ;
        RECT 503.550 713.400 505.350 719.250 ;
        RECT 539.400 713.400 541.200 719.250 ;
        RECT 444.450 705.600 446.250 705.900 ;
        RECT 454.050 702.150 454.950 706.800 ;
        RECT 460.950 705.600 465.150 706.800 ;
        RECT 464.250 703.800 466.050 705.600 ;
        RECT 445.950 701.100 448.050 702.150 ;
        RECT 437.100 699.150 438.900 700.950 ;
        RECT 440.100 700.050 448.050 701.100 ;
        RECT 451.950 700.050 454.950 702.150 ;
        RECT 440.100 699.300 441.900 700.050 ;
        RECT 438.000 698.400 438.900 699.150 ;
        RECT 443.100 698.400 444.900 699.000 ;
        RECT 438.000 697.200 444.900 698.400 ;
        RECT 443.850 696.000 444.900 697.200 ;
        RECT 454.050 696.000 454.950 700.050 ;
        RECT 463.950 699.750 466.050 700.050 ;
        RECT 462.150 697.950 466.050 699.750 ;
        RECT 467.250 697.950 468.450 707.400 ;
        RECT 503.400 700.950 504.600 713.400 ;
        RECT 538.950 711.450 541.050 712.050 ;
        RECT 536.550 710.550 541.050 711.450 ;
        RECT 500.100 699.150 501.900 700.950 ;
        RECT 443.850 695.100 454.950 696.000 ;
        RECT 463.950 695.850 468.450 697.950 ;
        RECT 499.950 697.050 502.050 699.150 ;
        RECT 502.950 698.850 505.050 700.950 ;
        RECT 536.550 699.450 537.450 710.550 ;
        RECT 538.950 709.950 541.050 710.550 ;
        RECT 542.700 707.400 544.500 719.250 ;
        RECT 546.900 707.400 548.700 719.250 ;
        RECT 584.400 713.400 586.200 719.250 ;
        RECT 587.700 707.400 589.500 719.250 ;
        RECT 591.900 707.400 593.700 719.250 ;
        RECT 626.400 713.400 628.200 719.250 ;
        RECT 629.700 707.400 631.500 719.250 ;
        RECT 633.900 707.400 635.700 719.250 ;
        RECT 668.550 713.400 670.350 719.250 ;
        RECT 539.250 705.150 541.050 706.950 ;
        RECT 538.950 703.050 541.050 705.150 ;
        RECT 542.850 702.150 544.050 707.400 ;
        RECT 584.250 705.150 586.050 706.950 ;
        RECT 548.100 702.150 549.900 703.950 ;
        RECT 583.950 703.050 586.050 705.150 ;
        RECT 587.850 702.150 589.050 707.400 ;
        RECT 626.250 705.150 628.050 706.950 ;
        RECT 593.100 702.150 594.900 703.950 ;
        RECT 625.950 703.050 628.050 705.150 ;
        RECT 629.850 702.150 631.050 707.400 ;
        RECT 668.550 706.500 669.750 713.400 ;
        RECT 671.850 707.400 673.650 719.250 ;
        RECT 674.850 707.400 676.650 719.250 ;
        RECT 710.550 713.400 712.350 719.250 ;
        RECT 668.550 705.600 674.250 706.500 ;
        RECT 672.000 704.700 674.250 705.600 ;
        RECT 635.100 702.150 636.900 703.950 ;
        RECT 668.100 702.150 669.900 703.950 ;
        RECT 541.950 700.050 544.050 702.150 ;
        RECT 538.950 699.450 541.050 700.050 ;
        RECT 443.850 694.200 444.900 695.100 ;
        RECT 454.050 694.800 454.950 695.100 ;
        RECT 326.550 687.750 328.350 690.600 ;
        RECT 329.550 687.750 331.350 690.600 ;
        RECT 332.550 687.750 334.350 690.600 ;
        RECT 335.550 687.750 337.350 693.600 ;
        RECT 372.000 687.750 373.800 693.600 ;
        RECT 376.200 691.950 381.900 693.600 ;
        RECT 376.200 687.750 378.000 691.950 ;
        RECT 379.500 687.750 381.300 690.600 ;
        RECT 421.800 687.750 423.600 693.600 ;
        RECT 426.000 687.750 427.800 693.600 ;
        RECT 430.200 687.750 432.000 693.600 ;
        RECT 435.150 687.750 436.950 693.600 ;
        RECT 439.950 691.500 442.050 693.600 ;
        RECT 443.550 692.400 445.350 694.200 ;
        RECT 446.850 693.450 448.650 694.200 ;
        RECT 446.850 692.400 451.800 693.450 ;
        RECT 454.050 693.000 455.850 694.800 ;
        RECT 467.250 693.600 468.450 695.850 ;
        RECT 460.950 692.700 463.050 693.600 ;
        RECT 441.000 690.600 442.050 691.500 ;
        RECT 450.750 690.600 451.800 692.400 ;
        RECT 459.300 691.500 463.050 692.700 ;
        RECT 459.300 690.600 460.350 691.500 ;
        RECT 438.150 687.750 439.950 690.600 ;
        RECT 441.000 689.700 444.750 690.600 ;
        RECT 442.950 687.750 444.750 689.700 ;
        RECT 447.450 687.750 449.250 690.600 ;
        RECT 450.750 687.750 452.550 690.600 ;
        RECT 454.650 687.750 456.450 690.600 ;
        RECT 458.850 687.750 460.650 690.600 ;
        RECT 463.350 687.750 465.150 690.600 ;
        RECT 466.650 687.750 468.450 693.600 ;
        RECT 503.400 690.600 504.600 698.850 ;
        RECT 536.550 698.550 541.050 699.450 ;
        RECT 538.950 697.950 541.050 698.550 ;
        RECT 541.950 696.750 543.150 700.050 ;
        RECT 544.950 698.850 547.050 700.950 ;
        RECT 547.950 700.050 550.050 702.150 ;
        RECT 586.950 700.050 589.050 702.150 ;
        RECT 545.100 697.050 546.900 698.850 ;
        RECT 586.950 696.750 588.150 700.050 ;
        RECT 589.950 698.850 592.050 700.950 ;
        RECT 592.950 700.050 595.050 702.150 ;
        RECT 628.950 700.050 631.050 702.150 ;
        RECT 590.100 697.050 591.900 698.850 ;
        RECT 628.950 696.750 630.150 700.050 ;
        RECT 631.950 698.850 634.050 700.950 ;
        RECT 634.950 700.050 637.050 702.150 ;
        RECT 667.950 700.050 670.050 702.150 ;
        RECT 632.100 697.050 633.900 698.850 ;
        RECT 539.250 695.700 543.000 696.750 ;
        RECT 584.250 695.700 588.000 696.750 ;
        RECT 626.250 695.700 630.000 696.750 ;
        RECT 672.000 696.300 673.050 704.700 ;
        RECT 675.150 702.150 676.350 707.400 ;
        RECT 710.550 706.500 711.750 713.400 ;
        RECT 713.850 707.400 715.650 719.250 ;
        RECT 716.850 707.400 718.650 719.250 ;
        RECT 749.550 713.400 751.350 719.250 ;
        RECT 752.550 713.400 754.350 719.250 ;
        RECT 755.550 713.400 757.350 719.250 ;
        RECT 710.550 705.600 716.250 706.500 ;
        RECT 714.000 704.700 716.250 705.600 ;
        RECT 710.100 702.150 711.900 703.950 ;
        RECT 673.950 700.050 676.350 702.150 ;
        RECT 709.950 700.050 712.050 702.150 ;
        RECT 539.250 693.600 540.450 695.700 ;
        RECT 500.550 687.750 502.350 690.600 ;
        RECT 503.550 687.750 505.350 690.600 ;
        RECT 538.650 687.750 540.450 693.600 ;
        RECT 541.650 692.700 549.450 694.050 ;
        RECT 584.250 693.600 585.450 695.700 ;
        RECT 541.650 687.750 543.450 692.700 ;
        RECT 544.650 687.750 546.450 691.800 ;
        RECT 547.650 687.750 549.450 692.700 ;
        RECT 583.650 687.750 585.450 693.600 ;
        RECT 586.650 692.700 594.450 694.050 ;
        RECT 626.250 693.600 627.450 695.700 ;
        RECT 672.000 695.400 674.250 696.300 ;
        RECT 669.150 694.500 674.250 695.400 ;
        RECT 586.650 687.750 588.450 692.700 ;
        RECT 589.650 687.750 591.450 691.800 ;
        RECT 592.650 687.750 594.450 692.700 ;
        RECT 625.650 687.750 627.450 693.600 ;
        RECT 628.650 692.700 636.450 694.050 ;
        RECT 628.650 687.750 630.450 692.700 ;
        RECT 631.650 687.750 633.450 691.800 ;
        RECT 634.650 687.750 636.450 692.700 ;
        RECT 669.150 690.600 670.350 694.500 ;
        RECT 675.150 693.600 676.350 700.050 ;
        RECT 714.000 696.300 715.050 704.700 ;
        RECT 717.150 702.150 718.350 707.400 ;
        RECT 752.550 705.150 753.750 713.400 ;
        RECT 715.950 700.050 718.350 702.150 ;
        RECT 748.950 701.850 751.050 703.950 ;
        RECT 751.950 703.050 754.050 705.150 ;
        RECT 749.100 700.050 750.900 701.850 ;
        RECT 714.000 695.400 716.250 696.300 ;
        RECT 711.150 694.500 716.250 695.400 ;
        RECT 668.550 687.750 670.350 690.600 ;
        RECT 671.850 687.750 673.650 693.600 ;
        RECT 674.850 687.750 676.650 693.600 ;
        RECT 711.150 690.600 712.350 694.500 ;
        RECT 717.150 693.600 718.350 700.050 ;
        RECT 752.550 695.700 753.750 703.050 ;
        RECT 754.950 701.850 757.050 703.950 ;
        RECT 755.100 700.050 756.900 701.850 ;
        RECT 752.550 694.800 756.150 695.700 ;
        RECT 710.550 687.750 712.350 690.600 ;
        RECT 713.850 687.750 715.650 693.600 ;
        RECT 716.850 687.750 718.650 693.600 ;
        RECT 749.850 687.750 751.650 693.600 ;
        RECT 754.350 687.750 756.150 694.800 ;
        RECT 34.650 680.400 36.450 683.250 ;
        RECT 37.650 680.400 39.450 683.250 ;
        RECT 35.400 672.150 36.600 680.400 ;
        RECT 71.700 674.400 73.500 683.250 ;
        RECT 77.100 675.000 78.900 683.250 ;
        RECT 119.850 676.200 121.650 683.250 ;
        RECT 124.350 677.400 126.150 683.250 ;
        RECT 119.850 675.300 123.450 676.200 ;
        RECT 34.950 670.050 37.050 672.150 ;
        RECT 37.950 671.850 40.050 673.950 ;
        RECT 77.100 673.350 81.600 675.000 ;
        RECT 38.100 670.050 39.900 671.850 ;
        RECT 35.400 657.600 36.600 670.050 ;
        RECT 80.400 669.150 81.600 673.350 ;
        RECT 119.100 669.150 120.900 670.950 ;
        RECT 70.950 665.850 73.050 667.950 ;
        RECT 76.950 665.850 79.050 667.950 ;
        RECT 79.950 667.050 82.050 669.150 ;
        RECT 118.950 667.050 121.050 669.150 ;
        RECT 122.250 667.950 123.450 675.300 ;
        RECT 158.700 674.400 160.500 683.250 ;
        RECT 164.100 675.000 165.900 683.250 ;
        RECT 205.350 677.400 207.150 683.250 ;
        RECT 208.350 677.400 210.150 683.250 ;
        RECT 211.650 680.400 213.450 683.250 ;
        RECT 164.100 673.350 168.600 675.000 ;
        RECT 125.100 669.150 126.900 670.950 ;
        RECT 167.400 669.150 168.600 673.350 ;
        RECT 205.650 670.950 206.850 677.400 ;
        RECT 211.650 676.500 212.850 680.400 ;
        RECT 245.550 678.300 247.350 683.250 ;
        RECT 248.550 679.200 250.350 683.250 ;
        RECT 251.550 678.300 253.350 683.250 ;
        RECT 245.550 676.950 253.350 678.300 ;
        RECT 254.550 677.400 256.350 683.250 ;
        RECT 290.550 680.400 292.350 683.250 ;
        RECT 207.750 675.600 212.850 676.500 ;
        RECT 207.750 674.700 210.000 675.600 ;
        RECT 71.100 664.050 72.900 665.850 ;
        RECT 73.950 662.850 76.050 664.950 ;
        RECT 77.250 664.050 79.050 665.850 ;
        RECT 74.100 661.050 75.900 662.850 ;
        RECT 80.700 658.800 81.750 667.050 ;
        RECT 121.950 665.850 124.050 667.950 ;
        RECT 124.950 667.050 127.050 669.150 ;
        RECT 157.950 665.850 160.050 667.950 ;
        RECT 163.950 665.850 166.050 667.950 ;
        RECT 166.950 667.050 169.050 669.150 ;
        RECT 205.650 668.850 208.050 670.950 ;
        RECT 74.700 657.900 81.750 658.800 ;
        RECT 74.700 657.600 76.350 657.900 ;
        RECT 34.650 651.750 36.450 657.600 ;
        RECT 37.650 651.750 39.450 657.600 ;
        RECT 71.550 651.750 73.350 657.600 ;
        RECT 74.550 651.750 76.350 657.600 ;
        RECT 80.550 657.600 81.750 657.900 ;
        RECT 122.250 657.600 123.450 665.850 ;
        RECT 158.100 664.050 159.900 665.850 ;
        RECT 160.950 662.850 163.050 664.950 ;
        RECT 164.250 664.050 166.050 665.850 ;
        RECT 161.100 661.050 162.900 662.850 ;
        RECT 167.700 658.800 168.750 667.050 ;
        RECT 205.650 663.600 206.850 668.850 ;
        RECT 208.950 666.300 210.000 674.700 ;
        RECT 238.950 675.450 241.050 676.050 ;
        RECT 244.950 675.450 247.050 676.050 ;
        RECT 238.950 674.550 247.050 675.450 ;
        RECT 254.550 675.300 255.750 677.400 ;
        RECT 291.150 676.500 292.350 680.400 ;
        RECT 293.850 677.400 295.650 683.250 ;
        RECT 296.850 677.400 298.650 683.250 ;
        RECT 291.150 675.600 296.250 676.500 ;
        RECT 238.950 673.950 241.050 674.550 ;
        RECT 244.950 673.950 247.050 674.550 ;
        RECT 252.000 674.250 255.750 675.300 ;
        RECT 294.000 674.700 296.250 675.600 ;
        RECT 248.100 672.150 249.900 673.950 ;
        RECT 211.950 668.850 214.050 670.950 ;
        RECT 244.950 668.850 247.050 670.950 ;
        RECT 247.950 670.050 250.050 672.150 ;
        RECT 251.850 670.950 253.050 674.250 ;
        RECT 250.950 668.850 253.050 670.950 ;
        RECT 289.950 668.850 292.050 670.950 ;
        RECT 212.100 667.050 213.900 668.850 ;
        RECT 245.100 667.050 246.900 668.850 ;
        RECT 207.750 665.400 210.000 666.300 ;
        RECT 207.750 664.500 213.450 665.400 ;
        RECT 161.700 657.900 168.750 658.800 ;
        RECT 161.700 657.600 163.350 657.900 ;
        RECT 77.550 651.750 79.350 657.000 ;
        RECT 80.550 651.750 82.350 657.600 ;
        RECT 118.650 651.750 120.450 657.600 ;
        RECT 121.650 651.750 123.450 657.600 ;
        RECT 124.650 651.750 126.450 657.600 ;
        RECT 158.550 651.750 160.350 657.600 ;
        RECT 161.550 651.750 163.350 657.600 ;
        RECT 167.550 657.600 168.750 657.900 ;
        RECT 164.550 651.750 166.350 657.000 ;
        RECT 167.550 651.750 169.350 657.600 ;
        RECT 205.350 651.750 207.150 663.600 ;
        RECT 208.350 651.750 210.150 663.600 ;
        RECT 212.250 657.600 213.450 664.500 ;
        RECT 250.950 663.600 252.150 668.850 ;
        RECT 253.950 665.850 256.050 667.950 ;
        RECT 290.100 667.050 291.900 668.850 ;
        RECT 294.000 666.300 295.050 674.700 ;
        RECT 297.150 670.950 298.350 677.400 ;
        RECT 332.700 674.400 334.500 683.250 ;
        RECT 338.100 675.000 339.900 683.250 ;
        RECT 338.100 673.350 342.600 675.000 ;
        RECT 377.700 674.400 379.500 683.250 ;
        RECT 383.100 675.000 384.900 683.250 ;
        RECT 428.100 675.000 429.900 683.250 ;
        RECT 383.100 673.350 387.600 675.000 ;
        RECT 310.950 672.450 313.050 673.050 ;
        RECT 334.950 672.450 337.050 673.050 ;
        RECT 310.950 671.550 337.050 672.450 ;
        RECT 310.950 670.950 313.050 671.550 ;
        RECT 334.950 670.950 337.050 671.550 ;
        RECT 295.950 668.850 298.350 670.950 ;
        RECT 341.400 669.150 342.600 673.350 ;
        RECT 386.400 669.150 387.600 673.350 ;
        RECT 425.400 673.350 429.900 675.000 ;
        RECT 433.500 674.400 435.300 683.250 ;
        RECT 464.550 680.400 466.350 683.250 ;
        RECT 465.150 676.500 466.350 680.400 ;
        RECT 467.850 677.400 469.650 683.250 ;
        RECT 470.850 677.400 472.650 683.250 ;
        RECT 505.650 677.400 507.450 683.250 ;
        RECT 465.150 675.600 470.250 676.500 ;
        RECT 468.000 674.700 470.250 675.600 ;
        RECT 425.400 669.150 426.600 673.350 ;
        RECT 253.950 664.050 255.750 665.850 ;
        RECT 294.000 665.400 296.250 666.300 ;
        RECT 290.550 664.500 296.250 665.400 ;
        RECT 211.650 651.750 213.450 657.600 ;
        RECT 246.300 651.750 248.100 663.600 ;
        RECT 250.500 651.750 252.300 663.600 ;
        RECT 290.550 657.600 291.750 664.500 ;
        RECT 297.150 663.600 298.350 668.850 ;
        RECT 331.950 665.850 334.050 667.950 ;
        RECT 337.950 665.850 340.050 667.950 ;
        RECT 340.950 667.050 343.050 669.150 ;
        RECT 332.100 664.050 333.900 665.850 ;
        RECT 253.800 651.750 255.600 657.600 ;
        RECT 290.550 651.750 292.350 657.600 ;
        RECT 293.850 651.750 295.650 663.600 ;
        RECT 296.850 651.750 298.650 663.600 ;
        RECT 334.950 662.850 337.050 664.950 ;
        RECT 338.250 664.050 340.050 665.850 ;
        RECT 335.100 661.050 336.900 662.850 ;
        RECT 341.700 658.800 342.750 667.050 ;
        RECT 376.950 665.850 379.050 667.950 ;
        RECT 382.950 665.850 385.050 667.950 ;
        RECT 385.950 667.050 388.050 669.150 ;
        RECT 424.950 667.050 427.050 669.150 ;
        RECT 463.950 668.850 466.050 670.950 ;
        RECT 377.100 664.050 378.900 665.850 ;
        RECT 379.950 662.850 382.050 664.950 ;
        RECT 383.250 664.050 385.050 665.850 ;
        RECT 380.100 661.050 381.900 662.850 ;
        RECT 386.700 658.800 387.750 667.050 ;
        RECT 335.700 657.900 342.750 658.800 ;
        RECT 335.700 657.600 337.350 657.900 ;
        RECT 332.550 651.750 334.350 657.600 ;
        RECT 335.550 651.750 337.350 657.600 ;
        RECT 341.550 657.600 342.750 657.900 ;
        RECT 380.700 657.900 387.750 658.800 ;
        RECT 380.700 657.600 382.350 657.900 ;
        RECT 338.550 651.750 340.350 657.000 ;
        RECT 341.550 651.750 343.350 657.600 ;
        RECT 377.550 651.750 379.350 657.600 ;
        RECT 380.550 651.750 382.350 657.600 ;
        RECT 386.550 657.600 387.750 657.900 ;
        RECT 425.250 658.800 426.300 667.050 ;
        RECT 427.950 665.850 430.050 667.950 ;
        RECT 433.950 665.850 436.050 667.950 ;
        RECT 464.100 667.050 465.900 668.850 ;
        RECT 468.000 666.300 469.050 674.700 ;
        RECT 471.150 670.950 472.350 677.400 ;
        RECT 506.250 675.300 507.450 677.400 ;
        RECT 508.650 678.300 510.450 683.250 ;
        RECT 511.650 679.200 513.450 683.250 ;
        RECT 514.650 678.300 516.450 683.250 ;
        RECT 508.650 676.950 516.450 678.300 ;
        RECT 519.150 677.400 520.950 683.250 ;
        RECT 522.150 680.400 523.950 683.250 ;
        RECT 526.950 681.300 528.750 683.250 ;
        RECT 525.000 680.400 528.750 681.300 ;
        RECT 531.450 680.400 533.250 683.250 ;
        RECT 534.750 680.400 536.550 683.250 ;
        RECT 538.650 680.400 540.450 683.250 ;
        RECT 542.850 680.400 544.650 683.250 ;
        RECT 547.350 680.400 549.150 683.250 ;
        RECT 525.000 679.500 526.050 680.400 ;
        RECT 523.950 677.400 526.050 679.500 ;
        RECT 534.750 678.600 535.800 680.400 ;
        RECT 506.250 674.250 510.000 675.300 ;
        RECT 469.950 668.850 472.350 670.950 ;
        RECT 508.950 670.950 510.150 674.250 ;
        RECT 512.100 672.150 513.900 673.950 ;
        RECT 508.950 668.850 511.050 670.950 ;
        RECT 511.950 670.050 514.050 672.150 ;
        RECT 514.950 668.850 517.050 670.950 ;
        RECT 427.950 664.050 429.750 665.850 ;
        RECT 430.950 662.850 433.050 664.950 ;
        RECT 434.100 664.050 435.900 665.850 ;
        RECT 468.000 665.400 470.250 666.300 ;
        RECT 464.550 664.500 470.250 665.400 ;
        RECT 431.100 661.050 432.900 662.850 ;
        RECT 425.250 657.900 432.300 658.800 ;
        RECT 425.250 657.600 426.450 657.900 ;
        RECT 383.550 651.750 385.350 657.000 ;
        RECT 386.550 651.750 388.350 657.600 ;
        RECT 424.650 651.750 426.450 657.600 ;
        RECT 430.650 657.600 432.300 657.900 ;
        RECT 464.550 657.600 465.750 664.500 ;
        RECT 471.150 663.600 472.350 668.850 ;
        RECT 505.950 665.850 508.050 667.950 ;
        RECT 506.250 664.050 508.050 665.850 ;
        RECT 509.850 663.600 511.050 668.850 ;
        RECT 515.100 667.050 516.900 668.850 ;
        RECT 519.150 664.800 520.050 677.400 ;
        RECT 527.550 676.800 529.350 678.600 ;
        RECT 530.850 677.550 535.800 678.600 ;
        RECT 543.300 679.500 544.350 680.400 ;
        RECT 543.300 678.300 547.050 679.500 ;
        RECT 530.850 676.800 532.650 677.550 ;
        RECT 527.850 675.900 528.900 676.800 ;
        RECT 538.050 676.200 539.850 678.000 ;
        RECT 544.950 677.400 547.050 678.300 ;
        RECT 550.650 677.400 552.450 683.250 ;
        RECT 581.550 680.400 583.350 683.250 ;
        RECT 584.550 680.400 586.350 683.250 ;
        RECT 538.050 675.900 538.950 676.200 ;
        RECT 527.850 675.000 538.950 675.900 ;
        RECT 551.250 675.150 552.450 677.400 ;
        RECT 527.850 673.800 528.900 675.000 ;
        RECT 522.000 672.600 528.900 673.800 ;
        RECT 522.000 671.850 522.900 672.600 ;
        RECT 527.100 672.000 528.900 672.600 ;
        RECT 521.100 670.050 522.900 671.850 ;
        RECT 524.100 670.950 525.900 671.700 ;
        RECT 538.050 670.950 538.950 675.000 ;
        RECT 547.950 673.050 552.450 675.150 ;
        RECT 546.150 671.250 550.050 673.050 ;
        RECT 547.950 670.950 550.050 671.250 ;
        RECT 524.100 669.900 532.050 670.950 ;
        RECT 529.950 668.850 532.050 669.900 ;
        RECT 535.950 668.850 538.950 670.950 ;
        RECT 528.450 665.100 530.250 665.400 ;
        RECT 528.450 664.800 536.850 665.100 ;
        RECT 519.150 664.200 536.850 664.800 ;
        RECT 519.150 663.600 530.250 664.200 ;
        RECT 427.650 651.750 429.450 657.000 ;
        RECT 430.650 651.750 432.450 657.600 ;
        RECT 433.650 651.750 435.450 657.600 ;
        RECT 464.550 651.750 466.350 657.600 ;
        RECT 467.850 651.750 469.650 663.600 ;
        RECT 470.850 651.750 472.650 663.600 ;
        RECT 506.400 651.750 508.200 657.600 ;
        RECT 509.700 651.750 511.500 663.600 ;
        RECT 513.900 651.750 515.700 663.600 ;
        RECT 519.150 651.750 520.950 663.600 ;
        RECT 533.250 662.700 535.050 663.300 ;
        RECT 527.550 661.500 535.050 662.700 ;
        RECT 535.950 662.100 536.850 664.200 ;
        RECT 538.050 664.200 538.950 668.850 ;
        RECT 548.250 665.400 550.050 667.200 ;
        RECT 544.950 664.200 549.150 665.400 ;
        RECT 538.050 663.300 544.050 664.200 ;
        RECT 544.950 663.300 547.050 664.200 ;
        RECT 551.250 663.600 552.450 673.050 ;
        RECT 580.950 671.850 583.050 673.950 ;
        RECT 584.400 672.150 585.600 680.400 ;
        RECT 623.850 676.200 625.650 683.250 ;
        RECT 628.350 677.400 630.150 683.250 ;
        RECT 664.650 677.400 666.450 683.250 ;
        RECT 623.850 675.300 627.450 676.200 ;
        RECT 581.100 670.050 582.900 671.850 ;
        RECT 583.950 670.050 586.050 672.150 ;
        RECT 543.150 662.400 544.050 663.300 ;
        RECT 540.450 662.100 542.250 662.400 ;
        RECT 527.550 660.600 528.750 661.500 ;
        RECT 535.950 661.200 542.250 662.100 ;
        RECT 540.450 660.600 542.250 661.200 ;
        RECT 543.150 660.600 545.850 662.400 ;
        RECT 523.950 658.500 528.750 660.600 ;
        RECT 531.150 658.500 538.050 660.300 ;
        RECT 527.550 657.600 528.750 658.500 ;
        RECT 522.150 651.750 523.950 657.600 ;
        RECT 527.250 651.750 529.050 657.600 ;
        RECT 532.050 651.750 533.850 657.600 ;
        RECT 535.050 651.750 536.850 658.500 ;
        RECT 543.150 657.600 547.050 659.700 ;
        RECT 538.950 651.750 540.750 657.600 ;
        RECT 543.150 651.750 544.950 657.600 ;
        RECT 547.650 651.750 549.450 654.600 ;
        RECT 550.650 651.750 552.450 663.600 ;
        RECT 584.400 657.600 585.600 670.050 ;
        RECT 623.100 669.150 624.900 670.950 ;
        RECT 622.950 667.050 625.050 669.150 ;
        RECT 626.250 667.950 627.450 675.300 ;
        RECT 665.250 675.300 666.450 677.400 ;
        RECT 667.650 678.300 669.450 683.250 ;
        RECT 670.650 679.200 672.450 683.250 ;
        RECT 673.650 678.300 675.450 683.250 ;
        RECT 667.650 676.950 675.450 678.300 ;
        RECT 707.550 678.300 709.350 683.250 ;
        RECT 710.550 679.200 712.350 683.250 ;
        RECT 713.550 678.300 715.350 683.250 ;
        RECT 707.550 676.950 715.350 678.300 ;
        RECT 716.550 677.400 718.350 683.250 ;
        RECT 749.550 680.400 751.350 683.250 ;
        RECT 716.550 675.300 717.750 677.400 ;
        RECT 750.150 676.500 751.350 680.400 ;
        RECT 752.850 677.400 754.650 683.250 ;
        RECT 755.850 677.400 757.650 683.250 ;
        RECT 750.150 675.600 755.250 676.500 ;
        RECT 665.250 674.250 669.000 675.300 ;
        RECT 714.000 674.250 717.750 675.300 ;
        RECT 753.000 674.700 755.250 675.600 ;
        RECT 667.950 670.950 669.150 674.250 ;
        RECT 671.100 672.150 672.900 673.950 ;
        RECT 710.100 672.150 711.900 673.950 ;
        RECT 629.100 669.150 630.900 670.950 ;
        RECT 625.950 665.850 628.050 667.950 ;
        RECT 628.950 667.050 631.050 669.150 ;
        RECT 667.950 668.850 670.050 670.950 ;
        RECT 670.950 670.050 673.050 672.150 ;
        RECT 673.950 668.850 676.050 670.950 ;
        RECT 706.950 668.850 709.050 670.950 ;
        RECT 709.950 670.050 712.050 672.150 ;
        RECT 713.850 670.950 715.050 674.250 ;
        RECT 712.950 668.850 715.050 670.950 ;
        RECT 748.950 668.850 751.050 670.950 ;
        RECT 664.950 665.850 667.050 667.950 ;
        RECT 626.250 657.600 627.450 665.850 ;
        RECT 665.250 664.050 667.050 665.850 ;
        RECT 668.850 663.600 670.050 668.850 ;
        RECT 674.100 667.050 675.900 668.850 ;
        RECT 707.100 667.050 708.900 668.850 ;
        RECT 712.950 663.600 714.150 668.850 ;
        RECT 715.950 665.850 718.050 667.950 ;
        RECT 749.100 667.050 750.900 668.850 ;
        RECT 753.000 666.300 754.050 674.700 ;
        RECT 756.150 670.950 757.350 677.400 ;
        RECT 754.950 668.850 757.350 670.950 ;
        RECT 715.950 664.050 717.750 665.850 ;
        RECT 753.000 665.400 755.250 666.300 ;
        RECT 749.550 664.500 755.250 665.400 ;
        RECT 581.550 651.750 583.350 657.600 ;
        RECT 584.550 651.750 586.350 657.600 ;
        RECT 622.650 651.750 624.450 657.600 ;
        RECT 625.650 651.750 627.450 657.600 ;
        RECT 628.650 651.750 630.450 657.600 ;
        RECT 665.400 651.750 667.200 657.600 ;
        RECT 668.700 651.750 670.500 663.600 ;
        RECT 672.900 651.750 674.700 663.600 ;
        RECT 708.300 651.750 710.100 663.600 ;
        RECT 712.500 651.750 714.300 663.600 ;
        RECT 749.550 657.600 750.750 664.500 ;
        RECT 756.150 663.600 757.350 668.850 ;
        RECT 715.800 651.750 717.600 657.600 ;
        RECT 749.550 651.750 751.350 657.600 ;
        RECT 752.850 651.750 754.650 663.600 ;
        RECT 755.850 651.750 757.650 663.600 ;
        RECT 31.650 641.400 33.450 647.250 ;
        RECT 34.650 641.400 36.450 647.250 ;
        RECT 37.650 641.400 39.450 647.250 ;
        RECT 73.650 641.400 75.450 647.250 ;
        RECT 76.650 641.400 78.450 647.250 ;
        RECT 79.650 641.400 81.450 647.250 ;
        RECT 113.550 641.400 115.350 647.250 ;
        RECT 116.550 641.400 118.350 647.250 ;
        RECT 119.550 642.000 121.350 647.250 ;
        RECT 35.250 633.150 36.450 641.400 ;
        RECT 77.250 633.150 78.450 641.400 ;
        RECT 116.700 641.100 118.350 641.400 ;
        RECT 122.550 641.400 124.350 647.250 ;
        RECT 160.650 641.400 162.450 647.250 ;
        RECT 163.650 641.400 165.450 647.250 ;
        RECT 166.650 641.400 168.450 647.250 ;
        RECT 202.650 641.400 204.450 647.250 ;
        RECT 205.650 641.400 207.450 647.250 ;
        RECT 208.650 641.400 210.450 647.250 ;
        RECT 242.400 641.400 244.200 647.250 ;
        RECT 122.550 641.100 123.750 641.400 ;
        RECT 116.700 640.200 123.750 641.100 ;
        RECT 116.100 636.150 117.900 637.950 ;
        RECT 113.100 633.150 114.900 634.950 ;
        RECT 115.950 634.050 118.050 636.150 ;
        RECT 119.250 633.150 121.050 634.950 ;
        RECT 31.950 629.850 34.050 631.950 ;
        RECT 34.950 631.050 37.050 633.150 ;
        RECT 32.100 628.050 33.900 629.850 ;
        RECT 35.250 623.700 36.450 631.050 ;
        RECT 37.950 629.850 40.050 631.950 ;
        RECT 73.950 629.850 76.050 631.950 ;
        RECT 76.950 631.050 79.050 633.150 ;
        RECT 38.100 628.050 39.900 629.850 ;
        RECT 74.100 628.050 75.900 629.850 ;
        RECT 77.250 623.700 78.450 631.050 ;
        RECT 79.950 629.850 82.050 631.950 ;
        RECT 112.950 631.050 115.050 633.150 ;
        RECT 118.950 631.050 121.050 633.150 ;
        RECT 122.700 631.950 123.750 640.200 ;
        RECT 164.250 633.150 165.450 641.400 ;
        RECT 206.250 633.150 207.450 641.400 ;
        RECT 245.700 635.400 247.500 647.250 ;
        RECT 249.900 635.400 251.700 647.250 ;
        RECT 286.650 641.400 288.450 647.250 ;
        RECT 289.650 641.400 291.450 647.250 ;
        RECT 292.650 641.400 294.450 647.250 ;
        RECT 323.550 641.400 325.350 647.250 ;
        RECT 326.550 641.400 328.350 647.250 ;
        RECT 329.550 641.400 331.350 647.250 ;
        RECT 367.650 641.400 369.450 647.250 ;
        RECT 370.650 641.400 372.450 647.250 ;
        RECT 373.650 641.400 375.450 647.250 ;
        RECT 409.650 641.400 411.450 647.250 ;
        RECT 412.650 642.000 414.450 647.250 ;
        RECT 242.250 633.150 244.050 634.950 ;
        RECT 121.950 629.850 124.050 631.950 ;
        RECT 160.950 629.850 163.050 631.950 ;
        RECT 163.950 631.050 166.050 633.150 ;
        RECT 80.100 628.050 81.900 629.850 ;
        RECT 122.400 625.650 123.600 629.850 ;
        RECT 161.100 628.050 162.900 629.850 ;
        RECT 32.850 622.800 36.450 623.700 ;
        RECT 74.850 622.800 78.450 623.700 ;
        RECT 32.850 615.750 34.650 622.800 ;
        RECT 37.350 615.750 39.150 621.600 ;
        RECT 74.850 615.750 76.650 622.800 ;
        RECT 79.350 615.750 81.150 621.600 ;
        RECT 113.700 615.750 115.500 624.600 ;
        RECT 119.100 624.000 123.600 625.650 ;
        RECT 119.100 615.750 120.900 624.000 ;
        RECT 164.250 623.700 165.450 631.050 ;
        RECT 166.950 629.850 169.050 631.950 ;
        RECT 202.950 629.850 205.050 631.950 ;
        RECT 205.950 631.050 208.050 633.150 ;
        RECT 167.100 628.050 168.900 629.850 ;
        RECT 203.100 628.050 204.900 629.850 ;
        RECT 206.250 623.700 207.450 631.050 ;
        RECT 208.950 629.850 211.050 631.950 ;
        RECT 241.950 631.050 244.050 633.150 ;
        RECT 245.850 630.150 247.050 635.400 ;
        RECT 290.250 633.150 291.450 641.400 ;
        RECT 326.550 633.150 327.750 641.400 ;
        RECT 371.250 633.150 372.450 641.400 ;
        RECT 410.250 641.100 411.450 641.400 ;
        RECT 415.650 641.400 417.450 647.250 ;
        RECT 418.650 641.400 420.450 647.250 ;
        RECT 454.650 641.400 456.450 647.250 ;
        RECT 457.650 641.400 459.450 647.250 ;
        RECT 490.650 641.400 492.450 647.250 ;
        RECT 493.650 641.400 495.450 647.250 ;
        RECT 496.650 641.400 498.450 647.250 ;
        RECT 530.550 641.400 532.350 647.250 ;
        RECT 533.550 641.400 535.350 647.250 ;
        RECT 536.550 642.000 538.350 647.250 ;
        RECT 415.650 641.100 417.300 641.400 ;
        RECT 410.250 640.200 417.300 641.100 ;
        RECT 251.100 630.150 252.900 631.950 ;
        RECT 209.100 628.050 210.900 629.850 ;
        RECT 244.950 628.050 247.050 630.150 ;
        RECT 244.950 624.750 246.150 628.050 ;
        RECT 247.950 626.850 250.050 628.950 ;
        RECT 250.950 628.050 253.050 630.150 ;
        RECT 286.950 629.850 289.050 631.950 ;
        RECT 289.950 631.050 292.050 633.150 ;
        RECT 287.100 628.050 288.900 629.850 ;
        RECT 248.100 625.050 249.900 626.850 ;
        RECT 161.850 622.800 165.450 623.700 ;
        RECT 203.850 622.800 207.450 623.700 ;
        RECT 242.250 623.700 246.000 624.750 ;
        RECT 290.250 623.700 291.450 631.050 ;
        RECT 292.950 629.850 295.050 631.950 ;
        RECT 322.950 629.850 325.050 631.950 ;
        RECT 325.950 631.050 328.050 633.150 ;
        RECT 293.100 628.050 294.900 629.850 ;
        RECT 323.100 628.050 324.900 629.850 ;
        RECT 161.850 615.750 163.650 622.800 ;
        RECT 166.350 615.750 168.150 621.600 ;
        RECT 203.850 615.750 205.650 622.800 ;
        RECT 242.250 621.600 243.450 623.700 ;
        RECT 287.850 622.800 291.450 623.700 ;
        RECT 326.550 623.700 327.750 631.050 ;
        RECT 328.950 629.850 331.050 631.950 ;
        RECT 367.950 629.850 370.050 631.950 ;
        RECT 370.950 631.050 373.050 633.150 ;
        RECT 410.250 631.950 411.300 640.200 ;
        RECT 416.100 636.150 417.900 637.950 ;
        RECT 412.950 633.150 414.750 634.950 ;
        RECT 415.950 634.050 418.050 636.150 ;
        RECT 419.100 633.150 420.900 634.950 ;
        RECT 329.100 628.050 330.900 629.850 ;
        RECT 368.100 628.050 369.900 629.850 ;
        RECT 371.250 623.700 372.450 631.050 ;
        RECT 373.950 629.850 376.050 631.950 ;
        RECT 409.950 629.850 412.050 631.950 ;
        RECT 412.950 631.050 415.050 633.150 ;
        RECT 418.950 631.050 421.050 633.150 ;
        RECT 374.100 628.050 375.900 629.850 ;
        RECT 410.400 625.650 411.600 629.850 ;
        RECT 455.400 628.950 456.600 641.400 ;
        RECT 494.250 633.150 495.450 641.400 ;
        RECT 533.700 641.100 535.350 641.400 ;
        RECT 539.550 641.400 541.350 647.250 ;
        RECT 577.650 641.400 579.450 647.250 ;
        RECT 580.650 641.400 582.450 647.250 ;
        RECT 583.650 641.400 585.450 647.250 ;
        RECT 616.650 641.400 618.450 647.250 ;
        RECT 619.650 641.400 621.450 647.250 ;
        RECT 622.650 641.400 624.450 647.250 ;
        RECT 659.400 641.400 661.200 647.250 ;
        RECT 539.550 641.100 540.750 641.400 ;
        RECT 533.700 640.200 540.750 641.100 ;
        RECT 533.100 636.150 534.900 637.950 ;
        RECT 530.100 633.150 531.900 634.950 ;
        RECT 532.950 634.050 535.050 636.150 ;
        RECT 536.250 633.150 538.050 634.950 ;
        RECT 490.950 629.850 493.050 631.950 ;
        RECT 493.950 631.050 496.050 633.150 ;
        RECT 454.950 626.850 457.050 628.950 ;
        RECT 458.100 627.150 459.900 628.950 ;
        RECT 491.100 628.050 492.900 629.850 ;
        RECT 410.400 624.000 414.900 625.650 ;
        RECT 326.550 622.800 330.150 623.700 ;
        RECT 208.350 615.750 210.150 621.600 ;
        RECT 241.650 615.750 243.450 621.600 ;
        RECT 244.650 620.700 252.450 622.050 ;
        RECT 244.650 615.750 246.450 620.700 ;
        RECT 247.650 615.750 249.450 619.800 ;
        RECT 250.650 615.750 252.450 620.700 ;
        RECT 287.850 615.750 289.650 622.800 ;
        RECT 292.350 615.750 294.150 621.600 ;
        RECT 323.850 615.750 325.650 621.600 ;
        RECT 328.350 615.750 330.150 622.800 ;
        RECT 368.850 622.800 372.450 623.700 ;
        RECT 368.850 615.750 370.650 622.800 ;
        RECT 373.350 615.750 375.150 621.600 ;
        RECT 413.100 615.750 414.900 624.000 ;
        RECT 418.500 615.750 420.300 624.600 ;
        RECT 455.400 618.600 456.600 626.850 ;
        RECT 457.950 625.050 460.050 627.150 ;
        RECT 494.250 623.700 495.450 631.050 ;
        RECT 496.950 629.850 499.050 631.950 ;
        RECT 529.950 631.050 532.050 633.150 ;
        RECT 535.950 631.050 538.050 633.150 ;
        RECT 539.700 631.950 540.750 640.200 ;
        RECT 581.250 633.150 582.450 641.400 ;
        RECT 620.250 633.150 621.450 641.400 ;
        RECT 662.700 635.400 664.500 647.250 ;
        RECT 666.900 635.400 668.700 647.250 ;
        RECT 701.550 641.400 703.350 647.250 ;
        RECT 659.250 633.150 661.050 634.950 ;
        RECT 538.950 629.850 541.050 631.950 ;
        RECT 577.950 629.850 580.050 631.950 ;
        RECT 580.950 631.050 583.050 633.150 ;
        RECT 497.100 628.050 498.900 629.850 ;
        RECT 508.950 627.450 511.050 628.050 ;
        RECT 532.950 627.450 535.050 628.050 ;
        RECT 508.950 626.550 535.050 627.450 ;
        RECT 508.950 625.950 511.050 626.550 ;
        RECT 532.950 625.950 535.050 626.550 ;
        RECT 539.400 625.650 540.600 629.850 ;
        RECT 578.100 628.050 579.900 629.850 ;
        RECT 491.850 622.800 495.450 623.700 ;
        RECT 454.650 615.750 456.450 618.600 ;
        RECT 457.650 615.750 459.450 618.600 ;
        RECT 491.850 615.750 493.650 622.800 ;
        RECT 496.350 615.750 498.150 621.600 ;
        RECT 530.700 615.750 532.500 624.600 ;
        RECT 536.100 624.000 540.600 625.650 ;
        RECT 536.100 615.750 537.900 624.000 ;
        RECT 581.250 623.700 582.450 631.050 ;
        RECT 583.950 629.850 586.050 631.950 ;
        RECT 616.950 629.850 619.050 631.950 ;
        RECT 619.950 631.050 622.050 633.150 ;
        RECT 584.100 628.050 585.900 629.850 ;
        RECT 617.100 628.050 618.900 629.850 ;
        RECT 620.250 623.700 621.450 631.050 ;
        RECT 622.950 629.850 625.050 631.950 ;
        RECT 658.950 631.050 661.050 633.150 ;
        RECT 662.850 630.150 664.050 635.400 ;
        RECT 701.550 634.500 702.750 641.400 ;
        RECT 704.850 635.400 706.650 647.250 ;
        RECT 707.850 635.400 709.650 647.250 ;
        RECT 743.550 641.400 745.350 647.250 ;
        RECT 701.550 633.600 707.250 634.500 ;
        RECT 705.000 632.700 707.250 633.600 ;
        RECT 668.100 630.150 669.900 631.950 ;
        RECT 701.100 630.150 702.900 631.950 ;
        RECT 623.100 628.050 624.900 629.850 ;
        RECT 661.950 628.050 664.050 630.150 ;
        RECT 661.950 624.750 663.150 628.050 ;
        RECT 664.950 626.850 667.050 628.950 ;
        RECT 667.950 628.050 670.050 630.150 ;
        RECT 700.950 628.050 703.050 630.150 ;
        RECT 665.100 625.050 666.900 626.850 ;
        RECT 578.850 622.800 582.450 623.700 ;
        RECT 617.850 622.800 621.450 623.700 ;
        RECT 659.250 623.700 663.000 624.750 ;
        RECT 705.000 624.300 706.050 632.700 ;
        RECT 708.150 630.150 709.350 635.400 ;
        RECT 743.550 634.500 744.750 641.400 ;
        RECT 746.850 635.400 748.650 647.250 ;
        RECT 749.850 635.400 751.650 647.250 ;
        RECT 743.550 633.600 749.250 634.500 ;
        RECT 747.000 632.700 749.250 633.600 ;
        RECT 743.100 630.150 744.900 631.950 ;
        RECT 706.950 628.050 709.350 630.150 ;
        RECT 742.950 628.050 745.050 630.150 ;
        RECT 578.850 615.750 580.650 622.800 ;
        RECT 583.350 615.750 585.150 621.600 ;
        RECT 617.850 615.750 619.650 622.800 ;
        RECT 659.250 621.600 660.450 623.700 ;
        RECT 705.000 623.400 707.250 624.300 ;
        RECT 702.150 622.500 707.250 623.400 ;
        RECT 622.350 615.750 624.150 621.600 ;
        RECT 658.650 615.750 660.450 621.600 ;
        RECT 661.650 620.700 669.450 622.050 ;
        RECT 661.650 615.750 663.450 620.700 ;
        RECT 664.650 615.750 666.450 619.800 ;
        RECT 667.650 615.750 669.450 620.700 ;
        RECT 702.150 618.600 703.350 622.500 ;
        RECT 708.150 621.600 709.350 628.050 ;
        RECT 747.000 624.300 748.050 632.700 ;
        RECT 750.150 630.150 751.350 635.400 ;
        RECT 748.950 628.050 751.350 630.150 ;
        RECT 747.000 623.400 749.250 624.300 ;
        RECT 744.150 622.500 749.250 623.400 ;
        RECT 701.550 615.750 703.350 618.600 ;
        RECT 704.850 615.750 706.650 621.600 ;
        RECT 707.850 615.750 709.650 621.600 ;
        RECT 744.150 618.600 745.350 622.500 ;
        RECT 750.150 621.600 751.350 628.050 ;
        RECT 743.550 615.750 745.350 618.600 ;
        RECT 746.850 615.750 748.650 621.600 ;
        RECT 749.850 615.750 751.650 621.600 ;
        RECT 34.650 608.400 36.450 611.250 ;
        RECT 37.650 608.400 39.450 611.250 ;
        RECT 40.650 608.400 42.450 611.250 ;
        RECT 73.650 608.400 75.450 611.250 ;
        RECT 76.650 608.400 78.450 611.250 ;
        RECT 37.950 601.950 39.000 608.400 ;
        RECT 37.950 599.850 40.050 601.950 ;
        RECT 74.400 600.150 75.600 608.400 ;
        RECT 81.150 605.400 82.950 611.250 ;
        RECT 84.150 608.400 85.950 611.250 ;
        RECT 88.950 609.300 90.750 611.250 ;
        RECT 87.000 608.400 90.750 609.300 ;
        RECT 93.450 608.400 95.250 611.250 ;
        RECT 96.750 608.400 98.550 611.250 ;
        RECT 100.650 608.400 102.450 611.250 ;
        RECT 104.850 608.400 106.650 611.250 ;
        RECT 109.350 608.400 111.150 611.250 ;
        RECT 87.000 607.500 88.050 608.400 ;
        RECT 85.950 605.400 88.050 607.500 ;
        RECT 96.750 606.600 97.800 608.400 ;
        RECT 34.950 596.850 37.050 598.950 ;
        RECT 35.100 595.050 36.900 596.850 ;
        RECT 37.950 592.650 39.000 599.850 ;
        RECT 40.950 596.850 43.050 598.950 ;
        RECT 73.950 598.050 76.050 600.150 ;
        RECT 76.950 599.850 79.050 601.950 ;
        RECT 77.100 598.050 78.900 599.850 ;
        RECT 41.100 595.050 42.900 596.850 ;
        RECT 36.450 591.600 39.000 592.650 ;
        RECT 36.450 579.750 38.250 591.600 ;
        RECT 40.650 579.750 42.450 591.600 ;
        RECT 74.400 585.600 75.600 598.050 ;
        RECT 81.150 592.800 82.050 605.400 ;
        RECT 89.550 604.800 91.350 606.600 ;
        RECT 92.850 605.550 97.800 606.600 ;
        RECT 105.300 607.500 106.350 608.400 ;
        RECT 105.300 606.300 109.050 607.500 ;
        RECT 92.850 604.800 94.650 605.550 ;
        RECT 89.850 603.900 90.900 604.800 ;
        RECT 100.050 604.200 101.850 606.000 ;
        RECT 106.950 605.400 109.050 606.300 ;
        RECT 112.650 605.400 114.450 611.250 ;
        RECT 100.050 603.900 100.950 604.200 ;
        RECT 89.850 603.000 100.950 603.900 ;
        RECT 113.250 603.150 114.450 605.400 ;
        RECT 89.850 601.800 90.900 603.000 ;
        RECT 84.000 600.600 90.900 601.800 ;
        RECT 84.000 599.850 84.900 600.600 ;
        RECT 89.100 600.000 90.900 600.600 ;
        RECT 83.100 598.050 84.900 599.850 ;
        RECT 86.100 598.950 87.900 599.700 ;
        RECT 100.050 598.950 100.950 603.000 ;
        RECT 109.950 601.050 114.450 603.150 ;
        RECT 146.700 602.400 148.500 611.250 ;
        RECT 152.100 603.000 153.900 611.250 ;
        RECT 188.550 603.900 190.350 611.250 ;
        RECT 193.050 605.400 194.850 611.250 ;
        RECT 196.050 606.900 197.850 611.250 ;
        RECT 233.550 608.400 235.350 611.250 ;
        RECT 236.550 608.400 238.350 611.250 ;
        RECT 239.550 608.400 241.350 611.250 ;
        RECT 196.050 605.400 199.350 606.900 ;
        RECT 194.250 603.900 196.050 604.500 ;
        RECT 152.100 601.350 156.600 603.000 ;
        RECT 188.550 602.700 196.050 603.900 ;
        RECT 108.150 599.250 112.050 601.050 ;
        RECT 109.950 598.950 112.050 599.250 ;
        RECT 86.100 597.900 94.050 598.950 ;
        RECT 91.950 596.850 94.050 597.900 ;
        RECT 97.950 596.850 100.950 598.950 ;
        RECT 90.450 593.100 92.250 593.400 ;
        RECT 90.450 592.800 98.850 593.100 ;
        RECT 81.150 592.200 98.850 592.800 ;
        RECT 81.150 591.600 92.250 592.200 ;
        RECT 73.650 579.750 75.450 585.600 ;
        RECT 76.650 579.750 78.450 585.600 ;
        RECT 81.150 579.750 82.950 591.600 ;
        RECT 95.250 590.700 97.050 591.300 ;
        RECT 89.550 589.500 97.050 590.700 ;
        RECT 97.950 590.100 98.850 592.200 ;
        RECT 100.050 592.200 100.950 596.850 ;
        RECT 110.250 593.400 112.050 595.200 ;
        RECT 106.950 592.200 111.150 593.400 ;
        RECT 100.050 591.300 106.050 592.200 ;
        RECT 106.950 591.300 109.050 592.200 ;
        RECT 113.250 591.600 114.450 601.050 ;
        RECT 155.400 597.150 156.600 601.350 ;
        RECT 145.950 593.850 148.050 595.950 ;
        RECT 151.950 593.850 154.050 595.950 ;
        RECT 154.950 595.050 157.050 597.150 ;
        RECT 187.950 596.850 190.050 598.950 ;
        RECT 188.100 595.050 189.900 596.850 ;
        RECT 146.100 592.050 147.900 593.850 ;
        RECT 105.150 590.400 106.050 591.300 ;
        RECT 102.450 590.100 104.250 590.400 ;
        RECT 89.550 588.600 90.750 589.500 ;
        RECT 97.950 589.200 104.250 590.100 ;
        RECT 102.450 588.600 104.250 589.200 ;
        RECT 105.150 588.600 107.850 590.400 ;
        RECT 85.950 586.500 90.750 588.600 ;
        RECT 93.150 586.500 100.050 588.300 ;
        RECT 89.550 585.600 90.750 586.500 ;
        RECT 84.150 579.750 85.950 585.600 ;
        RECT 89.250 579.750 91.050 585.600 ;
        RECT 94.050 579.750 95.850 585.600 ;
        RECT 97.050 579.750 98.850 586.500 ;
        RECT 105.150 585.600 109.050 587.700 ;
        RECT 100.950 579.750 102.750 585.600 ;
        RECT 105.150 579.750 106.950 585.600 ;
        RECT 109.650 579.750 111.450 582.600 ;
        RECT 112.650 579.750 114.450 591.600 ;
        RECT 148.950 590.850 151.050 592.950 ;
        RECT 152.250 592.050 154.050 593.850 ;
        RECT 149.100 589.050 150.900 590.850 ;
        RECT 155.700 586.800 156.750 595.050 ;
        RECT 149.700 585.900 156.750 586.800 ;
        RECT 149.700 585.600 151.350 585.900 ;
        RECT 146.550 579.750 148.350 585.600 ;
        RECT 149.550 579.750 151.350 585.600 ;
        RECT 155.550 585.600 156.750 585.900 ;
        RECT 191.700 585.600 192.900 602.700 ;
        RECT 198.150 598.950 199.350 605.400 ;
        RECT 237.000 601.950 238.050 608.400 ;
        RECT 275.700 602.400 277.500 611.250 ;
        RECT 281.100 603.000 282.900 611.250 ;
        RECT 320.850 605.400 322.650 611.250 ;
        RECT 325.350 604.200 327.150 611.250 ;
        RECT 361.650 608.400 363.450 611.250 ;
        RECT 364.650 608.400 366.450 611.250 ;
        RECT 323.550 603.300 327.150 604.200 ;
        RECT 235.950 599.850 238.050 601.950 ;
        RECT 281.100 601.350 285.600 603.000 ;
        RECT 194.100 597.150 195.900 598.950 ;
        RECT 193.950 595.050 196.050 597.150 ;
        RECT 196.950 596.850 199.350 598.950 ;
        RECT 232.950 596.850 235.050 598.950 ;
        RECT 198.150 591.600 199.350 596.850 ;
        RECT 233.100 595.050 234.900 596.850 ;
        RECT 237.000 592.650 238.050 599.850 ;
        RECT 238.950 596.850 241.050 598.950 ;
        RECT 284.400 597.150 285.600 601.350 ;
        RECT 320.100 597.150 321.900 598.950 ;
        RECT 239.100 595.050 240.900 596.850 ;
        RECT 274.950 593.850 277.050 595.950 ;
        RECT 280.950 593.850 283.050 595.950 ;
        RECT 283.950 595.050 286.050 597.150 ;
        RECT 319.950 595.050 322.050 597.150 ;
        RECT 323.550 595.950 324.750 603.300 ;
        RECT 362.400 600.150 363.600 608.400 ;
        RECT 395.550 606.300 397.350 611.250 ;
        RECT 398.550 607.200 400.350 611.250 ;
        RECT 401.550 606.300 403.350 611.250 ;
        RECT 395.550 604.950 403.350 606.300 ;
        RECT 404.550 605.400 406.350 611.250 ;
        RECT 404.550 603.300 405.750 605.400 ;
        RECT 443.850 604.200 445.650 611.250 ;
        RECT 448.350 605.400 450.150 611.250 ;
        RECT 453.150 605.400 454.950 611.250 ;
        RECT 456.150 608.400 457.950 611.250 ;
        RECT 460.950 609.300 462.750 611.250 ;
        RECT 459.000 608.400 462.750 609.300 ;
        RECT 465.450 608.400 467.250 611.250 ;
        RECT 468.750 608.400 470.550 611.250 ;
        RECT 472.650 608.400 474.450 611.250 ;
        RECT 476.850 608.400 478.650 611.250 ;
        RECT 481.350 608.400 483.150 611.250 ;
        RECT 459.000 607.500 460.050 608.400 ;
        RECT 457.950 605.400 460.050 607.500 ;
        RECT 468.750 606.600 469.800 608.400 ;
        RECT 443.850 603.300 447.450 604.200 ;
        RECT 402.000 602.250 405.750 603.300 ;
        RECT 326.100 597.150 327.900 598.950 ;
        RECT 361.950 598.050 364.050 600.150 ;
        RECT 364.950 599.850 367.050 601.950 ;
        RECT 398.100 600.150 399.900 601.950 ;
        RECT 365.100 598.050 366.900 599.850 ;
        RECT 237.000 591.600 239.550 592.650 ;
        RECT 275.100 592.050 276.900 593.850 ;
        RECT 152.550 579.750 154.350 585.000 ;
        RECT 155.550 579.750 157.350 585.600 ;
        RECT 188.550 579.750 190.350 585.600 ;
        RECT 191.550 579.750 193.350 585.600 ;
        RECT 195.150 579.750 196.950 591.600 ;
        RECT 198.150 579.750 199.950 591.600 ;
        RECT 233.550 579.750 235.350 591.600 ;
        RECT 237.750 579.750 239.550 591.600 ;
        RECT 277.950 590.850 280.050 592.950 ;
        RECT 281.250 592.050 283.050 593.850 ;
        RECT 278.100 589.050 279.900 590.850 ;
        RECT 284.700 586.800 285.750 595.050 ;
        RECT 322.950 593.850 325.050 595.950 ;
        RECT 325.950 595.050 328.050 597.150 ;
        RECT 278.700 585.900 285.750 586.800 ;
        RECT 278.700 585.600 280.350 585.900 ;
        RECT 275.550 579.750 277.350 585.600 ;
        RECT 278.550 579.750 280.350 585.600 ;
        RECT 284.550 585.600 285.750 585.900 ;
        RECT 323.550 585.600 324.750 593.850 ;
        RECT 362.400 585.600 363.600 598.050 ;
        RECT 394.950 596.850 397.050 598.950 ;
        RECT 397.950 598.050 400.050 600.150 ;
        RECT 401.850 598.950 403.050 602.250 ;
        RECT 400.950 596.850 403.050 598.950 ;
        RECT 443.100 597.150 444.900 598.950 ;
        RECT 395.100 595.050 396.900 596.850 ;
        RECT 400.950 591.600 402.150 596.850 ;
        RECT 403.950 593.850 406.050 595.950 ;
        RECT 442.950 595.050 445.050 597.150 ;
        RECT 446.250 595.950 447.450 603.300 ;
        RECT 449.100 597.150 450.900 598.950 ;
        RECT 445.950 593.850 448.050 595.950 ;
        RECT 448.950 595.050 451.050 597.150 ;
        RECT 403.950 592.050 405.750 593.850 ;
        RECT 281.550 579.750 283.350 585.000 ;
        RECT 284.550 579.750 286.350 585.600 ;
        RECT 320.550 579.750 322.350 585.600 ;
        RECT 323.550 579.750 325.350 585.600 ;
        RECT 326.550 579.750 328.350 585.600 ;
        RECT 361.650 579.750 363.450 585.600 ;
        RECT 364.650 579.750 366.450 585.600 ;
        RECT 396.300 579.750 398.100 591.600 ;
        RECT 400.500 579.750 402.300 591.600 ;
        RECT 446.250 585.600 447.450 593.850 ;
        RECT 453.150 592.800 454.050 605.400 ;
        RECT 461.550 604.800 463.350 606.600 ;
        RECT 464.850 605.550 469.800 606.600 ;
        RECT 477.300 607.500 478.350 608.400 ;
        RECT 477.300 606.300 481.050 607.500 ;
        RECT 464.850 604.800 466.650 605.550 ;
        RECT 461.850 603.900 462.900 604.800 ;
        RECT 472.050 604.200 473.850 606.000 ;
        RECT 478.950 605.400 481.050 606.300 ;
        RECT 484.650 605.400 486.450 611.250 ;
        RECT 472.050 603.900 472.950 604.200 ;
        RECT 461.850 603.000 472.950 603.900 ;
        RECT 485.250 603.150 486.450 605.400 ;
        RECT 521.850 604.200 523.650 611.250 ;
        RECT 526.350 605.400 528.150 611.250 ;
        RECT 530.550 605.400 532.350 611.250 ;
        RECT 533.850 608.400 535.650 611.250 ;
        RECT 538.350 608.400 540.150 611.250 ;
        RECT 542.550 608.400 544.350 611.250 ;
        RECT 546.450 608.400 548.250 611.250 ;
        RECT 549.750 608.400 551.550 611.250 ;
        RECT 554.250 609.300 556.050 611.250 ;
        RECT 554.250 608.400 558.000 609.300 ;
        RECT 559.050 608.400 560.850 611.250 ;
        RECT 538.650 607.500 539.700 608.400 ;
        RECT 535.950 606.300 539.700 607.500 ;
        RECT 547.200 606.600 548.250 608.400 ;
        RECT 556.950 607.500 558.000 608.400 ;
        RECT 535.950 605.400 538.050 606.300 ;
        RECT 521.850 603.300 525.450 604.200 ;
        RECT 461.850 601.800 462.900 603.000 ;
        RECT 456.000 600.600 462.900 601.800 ;
        RECT 456.000 599.850 456.900 600.600 ;
        RECT 461.100 600.000 462.900 600.600 ;
        RECT 455.100 598.050 456.900 599.850 ;
        RECT 458.100 598.950 459.900 599.700 ;
        RECT 472.050 598.950 472.950 603.000 ;
        RECT 481.950 601.050 486.450 603.150 ;
        RECT 480.150 599.250 484.050 601.050 ;
        RECT 481.950 598.950 484.050 599.250 ;
        RECT 458.100 597.900 466.050 598.950 ;
        RECT 463.950 596.850 466.050 597.900 ;
        RECT 469.950 596.850 472.950 598.950 ;
        RECT 462.450 593.100 464.250 593.400 ;
        RECT 462.450 592.800 470.850 593.100 ;
        RECT 453.150 592.200 470.850 592.800 ;
        RECT 453.150 591.600 464.250 592.200 ;
        RECT 403.800 579.750 405.600 585.600 ;
        RECT 442.650 579.750 444.450 585.600 ;
        RECT 445.650 579.750 447.450 585.600 ;
        RECT 448.650 579.750 450.450 585.600 ;
        RECT 453.150 579.750 454.950 591.600 ;
        RECT 467.250 590.700 469.050 591.300 ;
        RECT 461.550 589.500 469.050 590.700 ;
        RECT 469.950 590.100 470.850 592.200 ;
        RECT 472.050 592.200 472.950 596.850 ;
        RECT 482.250 593.400 484.050 595.200 ;
        RECT 478.950 592.200 483.150 593.400 ;
        RECT 472.050 591.300 478.050 592.200 ;
        RECT 478.950 591.300 481.050 592.200 ;
        RECT 485.250 591.600 486.450 601.050 ;
        RECT 521.100 597.150 522.900 598.950 ;
        RECT 520.950 595.050 523.050 597.150 ;
        RECT 524.250 595.950 525.450 603.300 ;
        RECT 530.550 603.150 531.750 605.400 ;
        RECT 543.150 604.200 544.950 606.000 ;
        RECT 547.200 605.550 552.150 606.600 ;
        RECT 550.350 604.800 552.150 605.550 ;
        RECT 553.650 604.800 555.450 606.600 ;
        RECT 556.950 605.400 559.050 607.500 ;
        RECT 562.050 605.400 563.850 611.250 ;
        RECT 596.550 608.400 598.350 611.250 ;
        RECT 599.550 608.400 601.350 611.250 ;
        RECT 544.050 603.900 544.950 604.200 ;
        RECT 554.100 603.900 555.150 604.800 ;
        RECT 530.550 601.050 535.050 603.150 ;
        RECT 544.050 603.000 555.150 603.900 ;
        RECT 527.100 597.150 528.900 598.950 ;
        RECT 523.950 593.850 526.050 595.950 ;
        RECT 526.950 595.050 529.050 597.150 ;
        RECT 477.150 590.400 478.050 591.300 ;
        RECT 474.450 590.100 476.250 590.400 ;
        RECT 461.550 588.600 462.750 589.500 ;
        RECT 469.950 589.200 476.250 590.100 ;
        RECT 474.450 588.600 476.250 589.200 ;
        RECT 477.150 588.600 479.850 590.400 ;
        RECT 457.950 586.500 462.750 588.600 ;
        RECT 465.150 586.500 472.050 588.300 ;
        RECT 461.550 585.600 462.750 586.500 ;
        RECT 456.150 579.750 457.950 585.600 ;
        RECT 461.250 579.750 463.050 585.600 ;
        RECT 466.050 579.750 467.850 585.600 ;
        RECT 469.050 579.750 470.850 586.500 ;
        RECT 477.150 585.600 481.050 587.700 ;
        RECT 472.950 579.750 474.750 585.600 ;
        RECT 477.150 579.750 478.950 585.600 ;
        RECT 481.650 579.750 483.450 582.600 ;
        RECT 484.650 579.750 486.450 591.600 ;
        RECT 524.250 585.600 525.450 593.850 ;
        RECT 530.550 591.600 531.750 601.050 ;
        RECT 532.950 599.250 536.850 601.050 ;
        RECT 532.950 598.950 535.050 599.250 ;
        RECT 544.050 598.950 544.950 603.000 ;
        RECT 554.100 601.800 555.150 603.000 ;
        RECT 554.100 600.600 561.000 601.800 ;
        RECT 554.100 600.000 555.900 600.600 ;
        RECT 560.100 599.850 561.000 600.600 ;
        RECT 557.100 598.950 558.900 599.700 ;
        RECT 544.050 596.850 547.050 598.950 ;
        RECT 550.950 597.900 558.900 598.950 ;
        RECT 560.100 598.050 561.900 599.850 ;
        RECT 550.950 596.850 553.050 597.900 ;
        RECT 532.950 593.400 534.750 595.200 ;
        RECT 533.850 592.200 538.050 593.400 ;
        RECT 544.050 592.200 544.950 596.850 ;
        RECT 552.750 593.100 554.550 593.400 ;
        RECT 520.650 579.750 522.450 585.600 ;
        RECT 523.650 579.750 525.450 585.600 ;
        RECT 526.650 579.750 528.450 585.600 ;
        RECT 530.550 579.750 532.350 591.600 ;
        RECT 535.950 591.300 538.050 592.200 ;
        RECT 538.950 591.300 544.950 592.200 ;
        RECT 546.150 592.800 554.550 593.100 ;
        RECT 562.950 592.800 563.850 605.400 ;
        RECT 595.950 599.850 598.050 601.950 ;
        RECT 599.400 600.150 600.600 608.400 ;
        RECT 635.550 606.300 637.350 611.250 ;
        RECT 638.550 607.200 640.350 611.250 ;
        RECT 641.550 606.300 643.350 611.250 ;
        RECT 635.550 604.950 643.350 606.300 ;
        RECT 644.550 605.400 646.350 611.250 ;
        RECT 682.350 605.400 684.150 611.250 ;
        RECT 685.350 605.400 687.150 611.250 ;
        RECT 688.650 608.400 690.450 611.250 ;
        RECT 722.550 608.400 724.350 611.250 ;
        RECT 644.550 603.300 645.750 605.400 ;
        RECT 642.000 602.250 645.750 603.300 ;
        RECT 638.100 600.150 639.900 601.950 ;
        RECT 596.100 598.050 597.900 599.850 ;
        RECT 598.950 598.050 601.050 600.150 ;
        RECT 546.150 592.200 563.850 592.800 ;
        RECT 538.950 590.400 539.850 591.300 ;
        RECT 537.150 588.600 539.850 590.400 ;
        RECT 540.750 590.100 542.550 590.400 ;
        RECT 546.150 590.100 547.050 592.200 ;
        RECT 552.750 591.600 563.850 592.200 ;
        RECT 540.750 589.200 547.050 590.100 ;
        RECT 547.950 590.700 549.750 591.300 ;
        RECT 547.950 589.500 555.450 590.700 ;
        RECT 540.750 588.600 542.550 589.200 ;
        RECT 554.250 588.600 555.450 589.500 ;
        RECT 535.950 585.600 539.850 587.700 ;
        RECT 544.950 586.500 551.850 588.300 ;
        RECT 554.250 586.500 559.050 588.600 ;
        RECT 533.550 579.750 535.350 582.600 ;
        RECT 538.050 579.750 539.850 585.600 ;
        RECT 542.250 579.750 544.050 585.600 ;
        RECT 546.150 579.750 547.950 586.500 ;
        RECT 554.250 585.600 555.450 586.500 ;
        RECT 549.150 579.750 550.950 585.600 ;
        RECT 553.950 579.750 555.750 585.600 ;
        RECT 559.050 579.750 560.850 585.600 ;
        RECT 562.050 579.750 563.850 591.600 ;
        RECT 599.400 585.600 600.600 598.050 ;
        RECT 634.950 596.850 637.050 598.950 ;
        RECT 637.950 598.050 640.050 600.150 ;
        RECT 641.850 598.950 643.050 602.250 ;
        RECT 640.950 596.850 643.050 598.950 ;
        RECT 682.650 598.950 683.850 605.400 ;
        RECT 688.650 604.500 689.850 608.400 ;
        RECT 684.750 603.600 689.850 604.500 ;
        RECT 723.150 604.500 724.350 608.400 ;
        RECT 725.850 605.400 727.650 611.250 ;
        RECT 728.850 605.400 730.650 611.250 ;
        RECT 723.150 603.600 728.250 604.500 ;
        RECT 684.750 602.700 687.000 603.600 ;
        RECT 682.650 596.850 685.050 598.950 ;
        RECT 635.100 595.050 636.900 596.850 ;
        RECT 640.950 591.600 642.150 596.850 ;
        RECT 643.950 593.850 646.050 595.950 ;
        RECT 643.950 592.050 645.750 593.850 ;
        RECT 682.650 591.600 683.850 596.850 ;
        RECT 685.950 594.300 687.000 602.700 ;
        RECT 726.000 602.700 728.250 603.600 ;
        RECT 688.950 596.850 691.050 598.950 ;
        RECT 721.950 596.850 724.050 598.950 ;
        RECT 689.100 595.050 690.900 596.850 ;
        RECT 722.100 595.050 723.900 596.850 ;
        RECT 684.750 593.400 687.000 594.300 ;
        RECT 726.000 594.300 727.050 602.700 ;
        RECT 729.150 598.950 730.350 605.400 ;
        RECT 727.950 596.850 730.350 598.950 ;
        RECT 726.000 593.400 728.250 594.300 ;
        RECT 684.750 592.500 690.450 593.400 ;
        RECT 596.550 579.750 598.350 585.600 ;
        RECT 599.550 579.750 601.350 585.600 ;
        RECT 636.300 579.750 638.100 591.600 ;
        RECT 640.500 579.750 642.300 591.600 ;
        RECT 643.800 579.750 645.600 585.600 ;
        RECT 682.350 579.750 684.150 591.600 ;
        RECT 685.350 579.750 687.150 591.600 ;
        RECT 689.250 585.600 690.450 592.500 ;
        RECT 688.650 579.750 690.450 585.600 ;
        RECT 722.550 592.500 728.250 593.400 ;
        RECT 722.550 585.600 723.750 592.500 ;
        RECT 729.150 591.600 730.350 596.850 ;
        RECT 722.550 579.750 724.350 585.600 ;
        RECT 725.850 579.750 727.650 591.600 ;
        RECT 728.850 579.750 730.650 591.600 ;
        RECT 35.400 569.400 37.200 575.250 ;
        RECT 38.700 563.400 40.500 575.250 ;
        RECT 42.900 563.400 44.700 575.250 ;
        RECT 77.550 569.400 79.350 575.250 ;
        RECT 80.550 569.400 82.350 575.250 ;
        RECT 83.550 569.400 85.350 575.250 ;
        RECT 35.250 561.150 37.050 562.950 ;
        RECT 34.950 559.050 37.050 561.150 ;
        RECT 38.850 558.150 40.050 563.400 ;
        RECT 80.550 561.150 81.750 569.400 ;
        RECT 120.300 563.400 122.100 575.250 ;
        RECT 124.500 563.400 126.300 575.250 ;
        RECT 127.800 569.400 129.600 575.250 ;
        RECT 161.550 569.400 163.350 575.250 ;
        RECT 164.550 569.400 166.350 575.250 ;
        RECT 167.550 569.400 169.350 575.250 ;
        RECT 44.100 558.150 45.900 559.950 ;
        RECT 37.950 556.050 40.050 558.150 ;
        RECT 37.950 552.750 39.150 556.050 ;
        RECT 40.950 554.850 43.050 556.950 ;
        RECT 43.950 556.050 46.050 558.150 ;
        RECT 76.950 557.850 79.050 559.950 ;
        RECT 79.950 559.050 82.050 561.150 ;
        RECT 77.100 556.050 78.900 557.850 ;
        RECT 41.100 553.050 42.900 554.850 ;
        RECT 35.250 551.700 39.000 552.750 ;
        RECT 80.550 551.700 81.750 559.050 ;
        RECT 82.950 557.850 85.050 559.950 ;
        RECT 119.100 558.150 120.900 559.950 ;
        RECT 124.950 558.150 126.150 563.400 ;
        RECT 127.950 561.150 129.750 562.950 ;
        RECT 164.550 561.150 165.750 569.400 ;
        RECT 203.550 563.400 205.350 575.250 ;
        RECT 207.750 563.400 209.550 575.250 ;
        RECT 245.550 569.400 247.350 575.250 ;
        RECT 248.550 569.400 250.350 575.250 ;
        RECT 207.000 562.350 209.550 563.400 ;
        RECT 127.950 559.050 130.050 561.150 ;
        RECT 83.100 556.050 84.900 557.850 ;
        RECT 118.950 556.050 121.050 558.150 ;
        RECT 121.950 554.850 124.050 556.950 ;
        RECT 124.950 556.050 127.050 558.150 ;
        RECT 160.950 557.850 163.050 559.950 ;
        RECT 163.950 559.050 166.050 561.150 ;
        RECT 161.100 556.050 162.900 557.850 ;
        RECT 122.100 553.050 123.900 554.850 ;
        RECT 125.850 552.750 127.050 556.050 ;
        RECT 126.000 551.700 129.750 552.750 ;
        RECT 35.250 549.600 36.450 551.700 ;
        RECT 80.550 550.800 84.150 551.700 ;
        RECT 34.650 543.750 36.450 549.600 ;
        RECT 37.650 548.700 45.450 550.050 ;
        RECT 37.650 543.750 39.450 548.700 ;
        RECT 40.650 543.750 42.450 547.800 ;
        RECT 43.650 543.750 45.450 548.700 ;
        RECT 77.850 543.750 79.650 549.600 ;
        RECT 82.350 543.750 84.150 550.800 ;
        RECT 119.550 548.700 127.350 550.050 ;
        RECT 119.550 543.750 121.350 548.700 ;
        RECT 122.550 543.750 124.350 547.800 ;
        RECT 125.550 543.750 127.350 548.700 ;
        RECT 128.550 549.600 129.750 551.700 ;
        RECT 164.550 551.700 165.750 559.050 ;
        RECT 166.950 557.850 169.050 559.950 ;
        RECT 203.100 558.150 204.900 559.950 ;
        RECT 167.100 556.050 168.900 557.850 ;
        RECT 202.950 556.050 205.050 558.150 ;
        RECT 207.000 555.150 208.050 562.350 ;
        RECT 209.100 558.150 210.900 559.950 ;
        RECT 208.950 556.050 211.050 558.150 ;
        RECT 248.400 556.950 249.600 569.400 ;
        RECT 285.300 563.400 287.100 575.250 ;
        RECT 289.500 563.400 291.300 575.250 ;
        RECT 292.800 569.400 294.600 575.250 ;
        RECT 329.400 569.400 331.200 575.250 ;
        RECT 332.700 563.400 334.500 575.250 ;
        RECT 336.900 563.400 338.700 575.250 ;
        RECT 371.550 563.400 373.350 575.250 ;
        RECT 376.050 563.550 377.850 575.250 ;
        RECT 379.050 564.900 380.850 575.250 ;
        RECT 379.050 563.550 381.450 564.900 ;
        RECT 284.100 558.150 285.900 559.950 ;
        RECT 289.950 558.150 291.150 563.400 ;
        RECT 292.950 561.150 294.750 562.950 ;
        RECT 329.250 561.150 331.050 562.950 ;
        RECT 292.950 559.050 295.050 561.150 ;
        RECT 328.950 559.050 331.050 561.150 ;
        RECT 332.850 558.150 334.050 563.400 ;
        RECT 371.550 562.200 372.750 563.400 ;
        RECT 376.950 562.200 378.750 562.650 ;
        RECT 371.550 561.000 378.750 562.200 ;
        RECT 376.950 560.850 378.750 561.000 ;
        RECT 338.100 558.150 339.900 559.950 ;
        RECT 374.100 558.150 375.900 559.950 ;
        RECT 245.100 555.150 246.900 556.950 ;
        RECT 205.950 553.050 208.050 555.150 ;
        RECT 244.950 553.050 247.050 555.150 ;
        RECT 247.950 554.850 250.050 556.950 ;
        RECT 283.950 556.050 286.050 558.150 ;
        RECT 286.950 554.850 289.050 556.950 ;
        RECT 289.950 556.050 292.050 558.150 ;
        RECT 164.550 550.800 168.150 551.700 ;
        RECT 128.550 543.750 130.350 549.600 ;
        RECT 161.850 543.750 163.650 549.600 ;
        RECT 166.350 543.750 168.150 550.800 ;
        RECT 207.000 546.600 208.050 553.050 ;
        RECT 248.400 546.600 249.600 554.850 ;
        RECT 287.100 553.050 288.900 554.850 ;
        RECT 290.850 552.750 292.050 556.050 ;
        RECT 331.950 556.050 334.050 558.150 ;
        RECT 331.950 552.750 333.150 556.050 ;
        RECT 334.950 554.850 337.050 556.950 ;
        RECT 337.950 556.050 340.050 558.150 ;
        RECT 371.100 555.150 372.900 556.950 ;
        RECT 373.950 556.050 376.050 558.150 ;
        RECT 335.100 553.050 336.900 554.850 ;
        RECT 370.950 553.050 373.050 555.150 ;
        RECT 291.000 551.700 294.750 552.750 ;
        RECT 284.550 548.700 292.350 550.050 ;
        RECT 203.550 543.750 205.350 546.600 ;
        RECT 206.550 543.750 208.350 546.600 ;
        RECT 209.550 543.750 211.350 546.600 ;
        RECT 245.550 543.750 247.350 546.600 ;
        RECT 248.550 543.750 250.350 546.600 ;
        RECT 284.550 543.750 286.350 548.700 ;
        RECT 287.550 543.750 289.350 547.800 ;
        RECT 290.550 543.750 292.350 548.700 ;
        RECT 293.550 549.600 294.750 551.700 ;
        RECT 329.250 551.700 333.000 552.750 ;
        RECT 377.700 552.600 378.600 560.850 ;
        RECT 380.100 556.950 381.450 563.550 ;
        RECT 416.550 564.300 418.350 575.250 ;
        RECT 419.550 565.200 421.350 575.250 ;
        RECT 422.550 564.300 424.350 575.250 ;
        RECT 416.550 563.400 424.350 564.300 ;
        RECT 425.550 563.400 427.350 575.250 ;
        RECT 460.650 574.500 468.450 575.250 ;
        RECT 460.650 563.400 462.450 574.500 ;
        RECT 463.650 563.400 465.450 573.600 ;
        RECT 466.650 564.600 468.450 574.500 ;
        RECT 469.650 565.500 471.450 575.250 ;
        RECT 472.650 564.600 474.450 575.250 ;
        RECT 466.650 563.700 474.450 564.600 ;
        RECT 477.150 563.400 478.950 575.250 ;
        RECT 480.150 569.400 481.950 575.250 ;
        RECT 485.250 569.400 487.050 575.250 ;
        RECT 490.050 569.400 491.850 575.250 ;
        RECT 485.550 568.500 486.750 569.400 ;
        RECT 493.050 568.500 494.850 575.250 ;
        RECT 496.950 569.400 498.750 575.250 ;
        RECT 501.150 569.400 502.950 575.250 ;
        RECT 505.650 572.400 507.450 575.250 ;
        RECT 481.950 566.400 486.750 568.500 ;
        RECT 489.150 566.700 496.050 568.500 ;
        RECT 501.150 567.300 505.050 569.400 ;
        RECT 485.550 565.500 486.750 566.400 ;
        RECT 498.450 565.800 500.250 566.400 ;
        RECT 485.550 564.300 493.050 565.500 ;
        RECT 491.250 563.700 493.050 564.300 ;
        RECT 493.950 564.900 500.250 565.800 ;
        RECT 425.700 558.150 426.900 563.400 ;
        RECT 463.800 562.500 465.600 563.400 ;
        RECT 477.150 562.800 488.250 563.400 ;
        RECT 493.950 562.800 494.850 564.900 ;
        RECT 498.450 564.600 500.250 564.900 ;
        RECT 501.150 564.600 503.850 566.400 ;
        RECT 501.150 563.700 502.050 564.600 ;
        RECT 463.800 561.600 467.850 562.500 ;
        RECT 461.100 558.150 462.900 559.950 ;
        RECT 466.950 558.150 467.850 561.600 ;
        RECT 477.150 562.200 494.850 562.800 ;
        RECT 472.950 558.150 474.750 559.950 ;
        RECT 379.950 554.850 382.050 556.950 ;
        RECT 415.950 554.850 418.050 556.950 ;
        RECT 419.100 555.150 420.900 556.950 ;
        RECT 376.950 551.700 378.750 552.600 ;
        RECT 329.250 549.600 330.450 551.700 ;
        RECT 375.450 550.800 378.750 551.700 ;
        RECT 293.550 543.750 295.350 549.600 ;
        RECT 328.650 543.750 330.450 549.600 ;
        RECT 331.650 548.700 339.450 550.050 ;
        RECT 331.650 543.750 333.450 548.700 ;
        RECT 334.650 543.750 336.450 547.800 ;
        RECT 337.650 543.750 339.450 548.700 ;
        RECT 375.450 546.600 376.350 550.800 ;
        RECT 381.000 549.600 382.050 554.850 ;
        RECT 416.100 553.050 417.900 554.850 ;
        RECT 418.950 553.050 421.050 555.150 ;
        RECT 421.950 554.850 424.050 556.950 ;
        RECT 424.950 556.050 427.050 558.150 ;
        RECT 460.950 556.050 463.050 558.150 ;
        RECT 422.100 553.050 423.900 554.850 ;
        RECT 425.700 549.600 426.900 556.050 ;
        RECT 463.950 554.850 466.050 556.950 ;
        RECT 466.950 556.050 469.050 558.150 ;
        RECT 464.250 553.050 466.050 554.850 ;
        RECT 468.000 549.600 469.050 556.050 ;
        RECT 469.950 554.850 472.050 556.950 ;
        RECT 472.950 556.050 475.050 558.150 ;
        RECT 469.950 553.050 471.750 554.850 ;
        RECT 477.150 549.600 478.050 562.200 ;
        RECT 486.450 561.900 494.850 562.200 ;
        RECT 496.050 562.800 502.050 563.700 ;
        RECT 502.950 562.800 505.050 563.700 ;
        RECT 508.650 563.400 510.450 575.250 ;
        RECT 539.550 569.400 541.350 575.250 ;
        RECT 542.550 569.400 544.350 575.250 ;
        RECT 580.650 569.400 582.450 575.250 ;
        RECT 583.650 569.400 585.450 575.250 ;
        RECT 586.650 569.400 588.450 575.250 ;
        RECT 486.450 561.600 488.250 561.900 ;
        RECT 496.050 558.150 496.950 562.800 ;
        RECT 502.950 561.600 507.150 562.800 ;
        RECT 506.250 559.800 508.050 561.600 ;
        RECT 487.950 557.100 490.050 558.150 ;
        RECT 479.100 555.150 480.900 556.950 ;
        RECT 482.100 556.050 490.050 557.100 ;
        RECT 493.950 556.050 496.950 558.150 ;
        RECT 482.100 555.300 483.900 556.050 ;
        RECT 480.000 554.400 480.900 555.150 ;
        RECT 485.100 554.400 486.900 555.000 ;
        RECT 480.000 553.200 486.900 554.400 ;
        RECT 485.850 552.000 486.900 553.200 ;
        RECT 496.050 552.000 496.950 556.050 ;
        RECT 505.950 555.750 508.050 556.050 ;
        RECT 504.150 553.950 508.050 555.750 ;
        RECT 509.250 553.950 510.450 563.400 ;
        RECT 542.400 556.950 543.600 569.400 ;
        RECT 584.250 561.150 585.450 569.400 ;
        RECT 621.300 563.400 623.100 575.250 ;
        RECT 625.500 563.400 627.300 575.250 ;
        RECT 628.800 569.400 630.600 575.250 ;
        RECT 662.550 569.400 664.350 575.250 ;
        RECT 665.550 569.400 667.350 575.250 ;
        RECT 668.550 569.400 670.350 575.250 ;
        RECT 701.550 569.400 703.350 575.250 ;
        RECT 580.950 557.850 583.050 559.950 ;
        RECT 583.950 559.050 586.050 561.150 ;
        RECT 539.100 555.150 540.900 556.950 ;
        RECT 485.850 551.100 496.950 552.000 ;
        RECT 505.950 551.850 510.450 553.950 ;
        RECT 538.950 553.050 541.050 555.150 ;
        RECT 541.950 554.850 544.050 556.950 ;
        RECT 581.100 556.050 582.900 557.850 ;
        RECT 485.850 550.200 486.900 551.100 ;
        RECT 496.050 550.800 496.950 551.100 ;
        RECT 371.550 543.750 373.350 546.600 ;
        RECT 374.550 543.750 376.350 546.600 ;
        RECT 377.550 543.750 379.350 546.600 ;
        RECT 380.550 543.750 382.350 549.600 ;
        RECT 417.000 543.750 418.800 549.600 ;
        RECT 421.200 547.950 426.900 549.600 ;
        RECT 421.200 543.750 423.000 547.950 ;
        RECT 424.500 543.750 426.300 546.600 ;
        RECT 463.800 543.750 465.600 549.600 ;
        RECT 468.000 543.750 469.800 549.600 ;
        RECT 472.200 543.750 474.000 549.600 ;
        RECT 477.150 543.750 478.950 549.600 ;
        RECT 481.950 547.500 484.050 549.600 ;
        RECT 485.550 548.400 487.350 550.200 ;
        RECT 488.850 549.450 490.650 550.200 ;
        RECT 488.850 548.400 493.800 549.450 ;
        RECT 496.050 549.000 497.850 550.800 ;
        RECT 509.250 549.600 510.450 551.850 ;
        RECT 502.950 548.700 505.050 549.600 ;
        RECT 483.000 546.600 484.050 547.500 ;
        RECT 492.750 546.600 493.800 548.400 ;
        RECT 501.300 547.500 505.050 548.700 ;
        RECT 501.300 546.600 502.350 547.500 ;
        RECT 480.150 543.750 481.950 546.600 ;
        RECT 483.000 545.700 486.750 546.600 ;
        RECT 484.950 543.750 486.750 545.700 ;
        RECT 489.450 543.750 491.250 546.600 ;
        RECT 492.750 543.750 494.550 546.600 ;
        RECT 496.650 543.750 498.450 546.600 ;
        RECT 500.850 543.750 502.650 546.600 ;
        RECT 505.350 543.750 507.150 546.600 ;
        RECT 508.650 543.750 510.450 549.600 ;
        RECT 542.400 546.600 543.600 554.850 ;
        RECT 584.250 551.700 585.450 559.050 ;
        RECT 586.950 557.850 589.050 559.950 ;
        RECT 620.100 558.150 621.900 559.950 ;
        RECT 625.950 558.150 627.150 563.400 ;
        RECT 628.950 561.150 630.750 562.950 ;
        RECT 665.550 561.150 666.750 569.400 ;
        RECT 701.550 562.500 702.750 569.400 ;
        RECT 704.850 563.400 706.650 575.250 ;
        RECT 707.850 563.400 709.650 575.250 ;
        RECT 743.550 569.400 745.350 575.250 ;
        RECT 701.550 561.600 707.250 562.500 ;
        RECT 628.950 559.050 631.050 561.150 ;
        RECT 587.100 556.050 588.900 557.850 ;
        RECT 619.950 556.050 622.050 558.150 ;
        RECT 622.950 554.850 625.050 556.950 ;
        RECT 625.950 556.050 628.050 558.150 ;
        RECT 661.950 557.850 664.050 559.950 ;
        RECT 664.950 559.050 667.050 561.150 ;
        RECT 705.000 560.700 707.250 561.600 ;
        RECT 662.100 556.050 663.900 557.850 ;
        RECT 623.100 553.050 624.900 554.850 ;
        RECT 626.850 552.750 628.050 556.050 ;
        RECT 627.000 551.700 630.750 552.750 ;
        RECT 581.850 550.800 585.450 551.700 ;
        RECT 539.550 543.750 541.350 546.600 ;
        RECT 542.550 543.750 544.350 546.600 ;
        RECT 581.850 543.750 583.650 550.800 ;
        RECT 586.350 543.750 588.150 549.600 ;
        RECT 620.550 548.700 628.350 550.050 ;
        RECT 620.550 543.750 622.350 548.700 ;
        RECT 623.550 543.750 625.350 547.800 ;
        RECT 626.550 543.750 628.350 548.700 ;
        RECT 629.550 549.600 630.750 551.700 ;
        RECT 665.550 551.700 666.750 559.050 ;
        RECT 667.950 557.850 670.050 559.950 ;
        RECT 701.100 558.150 702.900 559.950 ;
        RECT 668.100 556.050 669.900 557.850 ;
        RECT 700.950 556.050 703.050 558.150 ;
        RECT 705.000 552.300 706.050 560.700 ;
        RECT 708.150 558.150 709.350 563.400 ;
        RECT 743.550 562.500 744.750 569.400 ;
        RECT 746.850 563.400 748.650 575.250 ;
        RECT 749.850 563.400 751.650 575.250 ;
        RECT 743.550 561.600 749.250 562.500 ;
        RECT 747.000 560.700 749.250 561.600 ;
        RECT 743.100 558.150 744.900 559.950 ;
        RECT 706.950 556.050 709.350 558.150 ;
        RECT 742.950 556.050 745.050 558.150 ;
        RECT 665.550 550.800 669.150 551.700 ;
        RECT 705.000 551.400 707.250 552.300 ;
        RECT 629.550 543.750 631.350 549.600 ;
        RECT 662.850 543.750 664.650 549.600 ;
        RECT 667.350 543.750 669.150 550.800 ;
        RECT 702.150 550.500 707.250 551.400 ;
        RECT 702.150 546.600 703.350 550.500 ;
        RECT 708.150 549.600 709.350 556.050 ;
        RECT 747.000 552.300 748.050 560.700 ;
        RECT 750.150 558.150 751.350 563.400 ;
        RECT 748.950 556.050 751.350 558.150 ;
        RECT 747.000 551.400 749.250 552.300 ;
        RECT 744.150 550.500 749.250 551.400 ;
        RECT 701.550 543.750 703.350 546.600 ;
        RECT 704.850 543.750 706.650 549.600 ;
        RECT 707.850 543.750 709.650 549.600 ;
        RECT 744.150 546.600 745.350 550.500 ;
        RECT 750.150 549.600 751.350 556.050 ;
        RECT 743.550 543.750 745.350 546.600 ;
        RECT 746.850 543.750 748.650 549.600 ;
        RECT 749.850 543.750 751.650 549.600 ;
        RECT 3.150 533.400 4.950 539.250 ;
        RECT 6.150 536.400 7.950 539.250 ;
        RECT 10.950 537.300 12.750 539.250 ;
        RECT 9.000 536.400 12.750 537.300 ;
        RECT 15.450 536.400 17.250 539.250 ;
        RECT 18.750 536.400 20.550 539.250 ;
        RECT 22.650 536.400 24.450 539.250 ;
        RECT 26.850 536.400 28.650 539.250 ;
        RECT 31.350 536.400 33.150 539.250 ;
        RECT 9.000 535.500 10.050 536.400 ;
        RECT 7.950 533.400 10.050 535.500 ;
        RECT 18.750 534.600 19.800 536.400 ;
        RECT 3.150 520.800 4.050 533.400 ;
        RECT 11.550 532.800 13.350 534.600 ;
        RECT 14.850 533.550 19.800 534.600 ;
        RECT 27.300 535.500 28.350 536.400 ;
        RECT 27.300 534.300 31.050 535.500 ;
        RECT 14.850 532.800 16.650 533.550 ;
        RECT 11.850 531.900 12.900 532.800 ;
        RECT 22.050 532.200 23.850 534.000 ;
        RECT 28.950 533.400 31.050 534.300 ;
        RECT 34.650 533.400 36.450 539.250 ;
        RECT 68.850 533.400 70.650 539.250 ;
        RECT 22.050 531.900 22.950 532.200 ;
        RECT 11.850 531.000 22.950 531.900 ;
        RECT 35.250 531.150 36.450 533.400 ;
        RECT 73.350 532.200 75.150 539.250 ;
        RECT 11.850 529.800 12.900 531.000 ;
        RECT 6.000 528.600 12.900 529.800 ;
        RECT 6.000 527.850 6.900 528.600 ;
        RECT 11.100 528.000 12.900 528.600 ;
        RECT 5.100 526.050 6.900 527.850 ;
        RECT 8.100 526.950 9.900 527.700 ;
        RECT 22.050 526.950 22.950 531.000 ;
        RECT 31.950 529.050 36.450 531.150 ;
        RECT 30.150 527.250 34.050 529.050 ;
        RECT 31.950 526.950 34.050 527.250 ;
        RECT 8.100 525.900 16.050 526.950 ;
        RECT 13.950 524.850 16.050 525.900 ;
        RECT 19.950 524.850 22.950 526.950 ;
        RECT 12.450 521.100 14.250 521.400 ;
        RECT 12.450 520.800 20.850 521.100 ;
        RECT 3.150 520.200 20.850 520.800 ;
        RECT 3.150 519.600 14.250 520.200 ;
        RECT 3.150 507.750 4.950 519.600 ;
        RECT 17.250 518.700 19.050 519.300 ;
        RECT 11.550 517.500 19.050 518.700 ;
        RECT 19.950 518.100 20.850 520.200 ;
        RECT 22.050 520.200 22.950 524.850 ;
        RECT 32.250 521.400 34.050 523.200 ;
        RECT 28.950 520.200 33.150 521.400 ;
        RECT 22.050 519.300 28.050 520.200 ;
        RECT 28.950 519.300 31.050 520.200 ;
        RECT 35.250 519.600 36.450 529.050 ;
        RECT 71.550 531.300 75.150 532.200 ;
        RECT 81.150 533.400 82.950 539.250 ;
        RECT 84.150 536.400 85.950 539.250 ;
        RECT 88.950 537.300 90.750 539.250 ;
        RECT 87.000 536.400 90.750 537.300 ;
        RECT 93.450 536.400 95.250 539.250 ;
        RECT 96.750 536.400 98.550 539.250 ;
        RECT 100.650 536.400 102.450 539.250 ;
        RECT 104.850 536.400 106.650 539.250 ;
        RECT 109.350 536.400 111.150 539.250 ;
        RECT 87.000 535.500 88.050 536.400 ;
        RECT 85.950 533.400 88.050 535.500 ;
        RECT 96.750 534.600 97.800 536.400 ;
        RECT 68.100 525.150 69.900 526.950 ;
        RECT 67.950 523.050 70.050 525.150 ;
        RECT 71.550 523.950 72.750 531.300 ;
        RECT 74.100 525.150 75.900 526.950 ;
        RECT 70.950 521.850 73.050 523.950 ;
        RECT 73.950 523.050 76.050 525.150 ;
        RECT 27.150 518.400 28.050 519.300 ;
        RECT 24.450 518.100 26.250 518.400 ;
        RECT 11.550 516.600 12.750 517.500 ;
        RECT 19.950 517.200 26.250 518.100 ;
        RECT 24.450 516.600 26.250 517.200 ;
        RECT 27.150 516.600 29.850 518.400 ;
        RECT 7.950 514.500 12.750 516.600 ;
        RECT 15.150 514.500 22.050 516.300 ;
        RECT 11.550 513.600 12.750 514.500 ;
        RECT 6.150 507.750 7.950 513.600 ;
        RECT 11.250 507.750 13.050 513.600 ;
        RECT 16.050 507.750 17.850 513.600 ;
        RECT 19.050 507.750 20.850 514.500 ;
        RECT 27.150 513.600 31.050 515.700 ;
        RECT 22.950 507.750 24.750 513.600 ;
        RECT 27.150 507.750 28.950 513.600 ;
        RECT 31.650 507.750 33.450 510.600 ;
        RECT 34.650 507.750 36.450 519.600 ;
        RECT 71.550 513.600 72.750 521.850 ;
        RECT 81.150 520.800 82.050 533.400 ;
        RECT 89.550 532.800 91.350 534.600 ;
        RECT 92.850 533.550 97.800 534.600 ;
        RECT 105.300 535.500 106.350 536.400 ;
        RECT 105.300 534.300 109.050 535.500 ;
        RECT 92.850 532.800 94.650 533.550 ;
        RECT 89.850 531.900 90.900 532.800 ;
        RECT 100.050 532.200 101.850 534.000 ;
        RECT 106.950 533.400 109.050 534.300 ;
        RECT 112.650 533.400 114.450 539.250 ;
        RECT 148.650 533.400 150.450 539.250 ;
        RECT 100.050 531.900 100.950 532.200 ;
        RECT 89.850 531.000 100.950 531.900 ;
        RECT 113.250 531.150 114.450 533.400 ;
        RECT 89.850 529.800 90.900 531.000 ;
        RECT 84.000 528.600 90.900 529.800 ;
        RECT 84.000 527.850 84.900 528.600 ;
        RECT 89.100 528.000 90.900 528.600 ;
        RECT 83.100 526.050 84.900 527.850 ;
        RECT 86.100 526.950 87.900 527.700 ;
        RECT 100.050 526.950 100.950 531.000 ;
        RECT 109.950 529.050 114.450 531.150 ;
        RECT 149.250 531.300 150.450 533.400 ;
        RECT 151.650 534.300 153.450 539.250 ;
        RECT 154.650 535.200 156.450 539.250 ;
        RECT 157.650 534.300 159.450 539.250 ;
        RECT 151.650 532.950 159.450 534.300 ;
        RECT 162.150 533.400 163.950 539.250 ;
        RECT 165.150 536.400 166.950 539.250 ;
        RECT 169.950 537.300 171.750 539.250 ;
        RECT 168.000 536.400 171.750 537.300 ;
        RECT 174.450 536.400 176.250 539.250 ;
        RECT 177.750 536.400 179.550 539.250 ;
        RECT 181.650 536.400 183.450 539.250 ;
        RECT 185.850 536.400 187.650 539.250 ;
        RECT 190.350 536.400 192.150 539.250 ;
        RECT 168.000 535.500 169.050 536.400 ;
        RECT 166.950 533.400 169.050 535.500 ;
        RECT 177.750 534.600 178.800 536.400 ;
        RECT 149.250 530.250 153.000 531.300 ;
        RECT 108.150 527.250 112.050 529.050 ;
        RECT 109.950 526.950 112.050 527.250 ;
        RECT 86.100 525.900 94.050 526.950 ;
        RECT 91.950 524.850 94.050 525.900 ;
        RECT 97.950 524.850 100.950 526.950 ;
        RECT 90.450 521.100 92.250 521.400 ;
        RECT 90.450 520.800 98.850 521.100 ;
        RECT 81.150 520.200 98.850 520.800 ;
        RECT 81.150 519.600 92.250 520.200 ;
        RECT 68.550 507.750 70.350 513.600 ;
        RECT 71.550 507.750 73.350 513.600 ;
        RECT 74.550 507.750 76.350 513.600 ;
        RECT 81.150 507.750 82.950 519.600 ;
        RECT 95.250 518.700 97.050 519.300 ;
        RECT 89.550 517.500 97.050 518.700 ;
        RECT 97.950 518.100 98.850 520.200 ;
        RECT 100.050 520.200 100.950 524.850 ;
        RECT 110.250 521.400 112.050 523.200 ;
        RECT 106.950 520.200 111.150 521.400 ;
        RECT 100.050 519.300 106.050 520.200 ;
        RECT 106.950 519.300 109.050 520.200 ;
        RECT 113.250 519.600 114.450 529.050 ;
        RECT 151.950 526.950 153.150 530.250 ;
        RECT 155.100 528.150 156.900 529.950 ;
        RECT 151.950 524.850 154.050 526.950 ;
        RECT 154.950 526.050 157.050 528.150 ;
        RECT 157.950 524.850 160.050 526.950 ;
        RECT 148.950 521.850 151.050 523.950 ;
        RECT 149.250 520.050 151.050 521.850 ;
        RECT 152.850 519.600 154.050 524.850 ;
        RECT 158.100 523.050 159.900 524.850 ;
        RECT 162.150 520.800 163.050 533.400 ;
        RECT 170.550 532.800 172.350 534.600 ;
        RECT 173.850 533.550 178.800 534.600 ;
        RECT 186.300 535.500 187.350 536.400 ;
        RECT 186.300 534.300 190.050 535.500 ;
        RECT 173.850 532.800 175.650 533.550 ;
        RECT 170.850 531.900 171.900 532.800 ;
        RECT 181.050 532.200 182.850 534.000 ;
        RECT 187.950 533.400 190.050 534.300 ;
        RECT 193.650 533.400 195.450 539.250 ;
        RECT 229.650 536.400 231.450 539.250 ;
        RECT 232.650 536.400 234.450 539.250 ;
        RECT 181.050 531.900 181.950 532.200 ;
        RECT 170.850 531.000 181.950 531.900 ;
        RECT 194.250 531.150 195.450 533.400 ;
        RECT 170.850 529.800 171.900 531.000 ;
        RECT 165.000 528.600 171.900 529.800 ;
        RECT 165.000 527.850 165.900 528.600 ;
        RECT 170.100 528.000 171.900 528.600 ;
        RECT 164.100 526.050 165.900 527.850 ;
        RECT 167.100 526.950 168.900 527.700 ;
        RECT 181.050 526.950 181.950 531.000 ;
        RECT 190.950 529.050 195.450 531.150 ;
        RECT 189.150 527.250 193.050 529.050 ;
        RECT 190.950 526.950 193.050 527.250 ;
        RECT 167.100 525.900 175.050 526.950 ;
        RECT 172.950 524.850 175.050 525.900 ;
        RECT 178.950 524.850 181.950 526.950 ;
        RECT 171.450 521.100 173.250 521.400 ;
        RECT 171.450 520.800 179.850 521.100 ;
        RECT 162.150 520.200 179.850 520.800 ;
        RECT 162.150 519.600 173.250 520.200 ;
        RECT 105.150 518.400 106.050 519.300 ;
        RECT 102.450 518.100 104.250 518.400 ;
        RECT 89.550 516.600 90.750 517.500 ;
        RECT 97.950 517.200 104.250 518.100 ;
        RECT 102.450 516.600 104.250 517.200 ;
        RECT 105.150 516.600 107.850 518.400 ;
        RECT 85.950 514.500 90.750 516.600 ;
        RECT 93.150 514.500 100.050 516.300 ;
        RECT 89.550 513.600 90.750 514.500 ;
        RECT 84.150 507.750 85.950 513.600 ;
        RECT 89.250 507.750 91.050 513.600 ;
        RECT 94.050 507.750 95.850 513.600 ;
        RECT 97.050 507.750 98.850 514.500 ;
        RECT 105.150 513.600 109.050 515.700 ;
        RECT 100.950 507.750 102.750 513.600 ;
        RECT 105.150 507.750 106.950 513.600 ;
        RECT 109.650 507.750 111.450 510.600 ;
        RECT 112.650 507.750 114.450 519.600 ;
        RECT 149.400 507.750 151.200 513.600 ;
        RECT 152.700 507.750 154.500 519.600 ;
        RECT 156.900 507.750 158.700 519.600 ;
        RECT 162.150 507.750 163.950 519.600 ;
        RECT 176.250 518.700 178.050 519.300 ;
        RECT 170.550 517.500 178.050 518.700 ;
        RECT 178.950 518.100 179.850 520.200 ;
        RECT 181.050 520.200 181.950 524.850 ;
        RECT 191.250 521.400 193.050 523.200 ;
        RECT 187.950 520.200 192.150 521.400 ;
        RECT 181.050 519.300 187.050 520.200 ;
        RECT 187.950 519.300 190.050 520.200 ;
        RECT 194.250 519.600 195.450 529.050 ;
        RECT 230.400 528.150 231.600 536.400 ;
        RECT 269.850 532.200 271.650 539.250 ;
        RECT 274.350 533.400 276.150 539.250 ;
        RECT 310.650 533.400 312.450 539.250 ;
        RECT 313.650 536.400 315.450 539.250 ;
        RECT 316.650 536.400 318.450 539.250 ;
        RECT 319.650 536.400 321.450 539.250 ;
        RECT 269.850 531.300 273.450 532.200 ;
        RECT 229.950 526.050 232.050 528.150 ;
        RECT 232.950 527.850 235.050 529.950 ;
        RECT 233.100 526.050 234.900 527.850 ;
        RECT 186.150 518.400 187.050 519.300 ;
        RECT 183.450 518.100 185.250 518.400 ;
        RECT 170.550 516.600 171.750 517.500 ;
        RECT 178.950 517.200 185.250 518.100 ;
        RECT 183.450 516.600 185.250 517.200 ;
        RECT 186.150 516.600 188.850 518.400 ;
        RECT 166.950 514.500 171.750 516.600 ;
        RECT 174.150 514.500 181.050 516.300 ;
        RECT 170.550 513.600 171.750 514.500 ;
        RECT 165.150 507.750 166.950 513.600 ;
        RECT 170.250 507.750 172.050 513.600 ;
        RECT 175.050 507.750 176.850 513.600 ;
        RECT 178.050 507.750 179.850 514.500 ;
        RECT 186.150 513.600 190.050 515.700 ;
        RECT 181.950 507.750 183.750 513.600 ;
        RECT 186.150 507.750 187.950 513.600 ;
        RECT 190.650 507.750 192.450 510.600 ;
        RECT 193.650 507.750 195.450 519.600 ;
        RECT 230.400 513.600 231.600 526.050 ;
        RECT 269.100 525.150 270.900 526.950 ;
        RECT 268.950 523.050 271.050 525.150 ;
        RECT 272.250 523.950 273.450 531.300 ;
        RECT 310.950 528.150 312.000 533.400 ;
        RECT 316.650 532.200 317.550 536.400 ;
        RECT 314.250 531.300 317.550 532.200 ;
        RECT 314.250 530.400 316.050 531.300 ;
        RECT 353.700 530.400 355.500 539.250 ;
        RECT 359.100 531.000 360.900 539.250 ;
        RECT 400.650 533.400 402.450 539.250 ;
        RECT 401.250 531.300 402.450 533.400 ;
        RECT 403.650 534.300 405.450 539.250 ;
        RECT 406.650 535.200 408.450 539.250 ;
        RECT 409.650 534.300 411.450 539.250 ;
        RECT 443.550 536.400 445.350 539.250 ;
        RECT 403.650 532.950 411.450 534.300 ;
        RECT 444.150 532.500 445.350 536.400 ;
        RECT 446.850 533.400 448.650 539.250 ;
        RECT 449.850 533.400 451.650 539.250 ;
        RECT 456.150 533.400 457.950 539.250 ;
        RECT 459.150 536.400 460.950 539.250 ;
        RECT 463.950 537.300 465.750 539.250 ;
        RECT 462.000 536.400 465.750 537.300 ;
        RECT 468.450 536.400 470.250 539.250 ;
        RECT 471.750 536.400 473.550 539.250 ;
        RECT 475.650 536.400 477.450 539.250 ;
        RECT 479.850 536.400 481.650 539.250 ;
        RECT 484.350 536.400 486.150 539.250 ;
        RECT 462.000 535.500 463.050 536.400 ;
        RECT 460.950 533.400 463.050 535.500 ;
        RECT 471.750 534.600 472.800 536.400 ;
        RECT 444.150 531.600 449.250 532.500 ;
        RECT 275.100 525.150 276.900 526.950 ;
        RECT 310.950 526.050 313.050 528.150 ;
        RECT 271.950 521.850 274.050 523.950 ;
        RECT 274.950 523.050 277.050 525.150 ;
        RECT 272.250 513.600 273.450 521.850 ;
        RECT 311.550 519.450 312.900 526.050 ;
        RECT 314.400 522.150 315.300 530.400 ;
        RECT 319.950 527.850 322.050 529.950 ;
        RECT 359.100 529.350 363.600 531.000 ;
        RECT 401.250 530.250 405.000 531.300 ;
        RECT 447.000 530.700 449.250 531.600 ;
        RECT 316.950 524.850 319.050 526.950 ;
        RECT 320.100 526.050 321.900 527.850 ;
        RECT 362.400 525.150 363.600 529.350 ;
        RECT 403.950 526.950 405.150 530.250 ;
        RECT 407.100 528.150 408.900 529.950 ;
        RECT 317.100 523.050 318.900 524.850 ;
        RECT 314.250 522.000 316.050 522.150 ;
        RECT 314.250 520.800 321.450 522.000 ;
        RECT 352.950 521.850 355.050 523.950 ;
        RECT 358.950 521.850 361.050 523.950 ;
        RECT 361.950 523.050 364.050 525.150 ;
        RECT 403.950 524.850 406.050 526.950 ;
        RECT 406.950 526.050 409.050 528.150 ;
        RECT 409.950 524.850 412.050 526.950 ;
        RECT 442.950 524.850 445.050 526.950 ;
        RECT 314.250 520.350 316.050 520.800 ;
        RECT 320.250 519.600 321.450 520.800 ;
        RECT 353.100 520.050 354.900 521.850 ;
        RECT 311.550 518.100 313.950 519.450 ;
        RECT 229.650 507.750 231.450 513.600 ;
        RECT 232.650 507.750 234.450 513.600 ;
        RECT 268.650 507.750 270.450 513.600 ;
        RECT 271.650 507.750 273.450 513.600 ;
        RECT 274.650 507.750 276.450 513.600 ;
        RECT 312.150 507.750 313.950 518.100 ;
        RECT 315.150 507.750 316.950 519.450 ;
        RECT 319.650 507.750 321.450 519.600 ;
        RECT 355.950 518.850 358.050 520.950 ;
        RECT 359.250 520.050 361.050 521.850 ;
        RECT 356.100 517.050 357.900 518.850 ;
        RECT 362.700 514.800 363.750 523.050 ;
        RECT 400.950 521.850 403.050 523.950 ;
        RECT 401.250 520.050 403.050 521.850 ;
        RECT 404.850 519.600 406.050 524.850 ;
        RECT 410.100 523.050 411.900 524.850 ;
        RECT 443.100 523.050 444.900 524.850 ;
        RECT 447.000 522.300 448.050 530.700 ;
        RECT 450.150 526.950 451.350 533.400 ;
        RECT 448.950 524.850 451.350 526.950 ;
        RECT 447.000 521.400 449.250 522.300 ;
        RECT 443.550 520.500 449.250 521.400 ;
        RECT 356.700 513.900 363.750 514.800 ;
        RECT 356.700 513.600 358.350 513.900 ;
        RECT 353.550 507.750 355.350 513.600 ;
        RECT 356.550 507.750 358.350 513.600 ;
        RECT 362.550 513.600 363.750 513.900 ;
        RECT 359.550 507.750 361.350 513.000 ;
        RECT 362.550 507.750 364.350 513.600 ;
        RECT 401.400 507.750 403.200 513.600 ;
        RECT 404.700 507.750 406.500 519.600 ;
        RECT 408.900 507.750 410.700 519.600 ;
        RECT 443.550 513.600 444.750 520.500 ;
        RECT 450.150 519.600 451.350 524.850 ;
        RECT 456.150 520.800 457.050 533.400 ;
        RECT 464.550 532.800 466.350 534.600 ;
        RECT 467.850 533.550 472.800 534.600 ;
        RECT 480.300 535.500 481.350 536.400 ;
        RECT 480.300 534.300 484.050 535.500 ;
        RECT 467.850 532.800 469.650 533.550 ;
        RECT 464.850 531.900 465.900 532.800 ;
        RECT 475.050 532.200 476.850 534.000 ;
        RECT 481.950 533.400 484.050 534.300 ;
        RECT 487.650 533.400 489.450 539.250 ;
        RECT 521.550 536.400 523.350 539.250 ;
        RECT 524.550 536.400 526.350 539.250 ;
        RECT 475.050 531.900 475.950 532.200 ;
        RECT 464.850 531.000 475.950 531.900 ;
        RECT 488.250 531.150 489.450 533.400 ;
        RECT 464.850 529.800 465.900 531.000 ;
        RECT 459.000 528.600 465.900 529.800 ;
        RECT 459.000 527.850 459.900 528.600 ;
        RECT 464.100 528.000 465.900 528.600 ;
        RECT 458.100 526.050 459.900 527.850 ;
        RECT 461.100 526.950 462.900 527.700 ;
        RECT 475.050 526.950 475.950 531.000 ;
        RECT 484.950 529.050 489.450 531.150 ;
        RECT 483.150 527.250 487.050 529.050 ;
        RECT 484.950 526.950 487.050 527.250 ;
        RECT 461.100 525.900 469.050 526.950 ;
        RECT 466.950 524.850 469.050 525.900 ;
        RECT 472.950 524.850 475.950 526.950 ;
        RECT 465.450 521.100 467.250 521.400 ;
        RECT 465.450 520.800 473.850 521.100 ;
        RECT 456.150 520.200 473.850 520.800 ;
        RECT 456.150 519.600 467.250 520.200 ;
        RECT 443.550 507.750 445.350 513.600 ;
        RECT 446.850 507.750 448.650 519.600 ;
        RECT 449.850 507.750 451.650 519.600 ;
        RECT 456.150 507.750 457.950 519.600 ;
        RECT 470.250 518.700 472.050 519.300 ;
        RECT 464.550 517.500 472.050 518.700 ;
        RECT 472.950 518.100 473.850 520.200 ;
        RECT 475.050 520.200 475.950 524.850 ;
        RECT 485.250 521.400 487.050 523.200 ;
        RECT 481.950 520.200 486.150 521.400 ;
        RECT 475.050 519.300 481.050 520.200 ;
        RECT 481.950 519.300 484.050 520.200 ;
        RECT 488.250 519.600 489.450 529.050 ;
        RECT 520.950 527.850 523.050 529.950 ;
        RECT 524.400 528.150 525.600 536.400 ;
        RECT 562.650 533.400 564.450 539.250 ;
        RECT 565.650 533.400 567.450 539.250 ;
        RECT 568.650 533.400 570.450 539.250 ;
        RECT 571.650 533.400 573.450 539.250 ;
        RECT 574.650 533.400 576.450 539.250 ;
        RECT 565.800 532.500 567.600 533.400 ;
        RECT 571.800 532.500 573.600 533.400 ;
        RECT 577.650 532.500 579.450 539.250 ;
        RECT 580.650 533.400 582.450 539.250 ;
        RECT 583.650 533.400 585.450 539.250 ;
        RECT 586.650 533.400 588.450 539.250 ;
        RECT 583.800 532.500 585.600 533.400 ;
        RECT 564.900 532.350 567.600 532.500 ;
        RECT 564.750 531.300 567.600 532.350 ;
        RECT 569.700 531.300 573.600 532.500 ;
        RECT 575.700 531.300 579.450 532.500 ;
        RECT 581.550 531.300 585.600 532.500 ;
        RECT 623.850 532.200 625.650 539.250 ;
        RECT 628.350 533.400 630.150 539.250 ;
        RECT 662.850 532.200 664.650 539.250 ;
        RECT 667.350 533.400 669.150 539.250 ;
        RECT 701.550 534.300 703.350 539.250 ;
        RECT 704.550 535.200 706.350 539.250 ;
        RECT 707.550 534.300 709.350 539.250 ;
        RECT 701.550 532.950 709.350 534.300 ;
        RECT 710.550 533.400 712.350 539.250 ;
        RECT 743.550 536.400 745.350 539.250 ;
        RECT 623.850 531.300 627.450 532.200 ;
        RECT 662.850 531.300 666.450 532.200 ;
        RECT 710.550 531.300 711.750 533.400 ;
        RECT 744.150 532.500 745.350 536.400 ;
        RECT 746.850 533.400 748.650 539.250 ;
        RECT 749.850 533.400 751.650 539.250 ;
        RECT 744.150 531.600 749.250 532.500 ;
        RECT 564.750 528.150 565.800 531.300 ;
        RECT 569.700 530.400 570.900 531.300 ;
        RECT 575.700 530.400 576.900 531.300 ;
        RECT 581.550 530.400 582.750 531.300 ;
        RECT 566.700 528.600 570.900 530.400 ;
        RECT 572.700 528.600 576.900 530.400 ;
        RECT 578.700 528.600 582.750 530.400 ;
        RECT 521.100 526.050 522.900 527.850 ;
        RECT 523.950 526.050 526.050 528.150 ;
        RECT 562.950 526.050 565.800 528.150 ;
        RECT 480.150 518.400 481.050 519.300 ;
        RECT 477.450 518.100 479.250 518.400 ;
        RECT 464.550 516.600 465.750 517.500 ;
        RECT 472.950 517.200 479.250 518.100 ;
        RECT 477.450 516.600 479.250 517.200 ;
        RECT 480.150 516.600 482.850 518.400 ;
        RECT 460.950 514.500 465.750 516.600 ;
        RECT 468.150 514.500 475.050 516.300 ;
        RECT 464.550 513.600 465.750 514.500 ;
        RECT 459.150 507.750 460.950 513.600 ;
        RECT 464.250 507.750 466.050 513.600 ;
        RECT 469.050 507.750 470.850 513.600 ;
        RECT 472.050 507.750 473.850 514.500 ;
        RECT 480.150 513.600 484.050 515.700 ;
        RECT 475.950 507.750 477.750 513.600 ;
        RECT 480.150 507.750 481.950 513.600 ;
        RECT 484.650 507.750 486.450 510.600 ;
        RECT 487.650 507.750 489.450 519.600 ;
        RECT 524.400 513.600 525.600 526.050 ;
        RECT 564.750 521.700 565.800 526.050 ;
        RECT 569.700 521.700 570.900 528.600 ;
        RECT 575.700 521.700 576.900 528.600 ;
        RECT 581.550 521.700 582.750 528.600 ;
        RECT 584.100 528.150 585.900 529.950 ;
        RECT 583.950 526.050 586.050 528.150 ;
        RECT 623.100 525.150 624.900 526.950 ;
        RECT 622.950 523.050 625.050 525.150 ;
        RECT 626.250 523.950 627.450 531.300 ;
        RECT 629.100 525.150 630.900 526.950 ;
        RECT 662.100 525.150 663.900 526.950 ;
        RECT 625.950 521.850 628.050 523.950 ;
        RECT 628.950 523.050 631.050 525.150 ;
        RECT 661.950 523.050 664.050 525.150 ;
        RECT 665.250 523.950 666.450 531.300 ;
        RECT 708.000 530.250 711.750 531.300 ;
        RECT 747.000 530.700 749.250 531.600 ;
        RECT 704.100 528.150 705.900 529.950 ;
        RECT 668.100 525.150 669.900 526.950 ;
        RECT 664.950 521.850 667.050 523.950 ;
        RECT 667.950 523.050 670.050 525.150 ;
        RECT 700.950 524.850 703.050 526.950 ;
        RECT 703.950 526.050 706.050 528.150 ;
        RECT 707.850 526.950 709.050 530.250 ;
        RECT 706.950 524.850 709.050 526.950 ;
        RECT 742.950 524.850 745.050 526.950 ;
        RECT 701.100 523.050 702.900 524.850 ;
        RECT 564.750 520.500 567.450 521.700 ;
        RECT 569.700 520.500 573.450 521.700 ;
        RECT 575.700 520.500 579.450 521.700 ;
        RECT 581.550 520.500 585.450 521.700 ;
        RECT 521.550 507.750 523.350 513.600 ;
        RECT 524.550 507.750 526.350 513.600 ;
        RECT 562.650 507.750 564.450 519.600 ;
        RECT 565.650 507.750 567.450 520.500 ;
        RECT 568.650 507.750 570.450 519.600 ;
        RECT 571.650 507.750 573.450 520.500 ;
        RECT 574.650 507.750 576.450 519.600 ;
        RECT 577.650 507.750 579.450 520.500 ;
        RECT 580.650 507.750 582.450 519.600 ;
        RECT 583.650 507.750 585.450 520.500 ;
        RECT 586.650 507.750 588.450 519.600 ;
        RECT 626.250 513.600 627.450 521.850 ;
        RECT 665.250 513.600 666.450 521.850 ;
        RECT 706.950 519.600 708.150 524.850 ;
        RECT 709.950 521.850 712.050 523.950 ;
        RECT 743.100 523.050 744.900 524.850 ;
        RECT 747.000 522.300 748.050 530.700 ;
        RECT 750.150 526.950 751.350 533.400 ;
        RECT 748.950 524.850 751.350 526.950 ;
        RECT 709.950 520.050 711.750 521.850 ;
        RECT 747.000 521.400 749.250 522.300 ;
        RECT 743.550 520.500 749.250 521.400 ;
        RECT 622.650 507.750 624.450 513.600 ;
        RECT 625.650 507.750 627.450 513.600 ;
        RECT 628.650 507.750 630.450 513.600 ;
        RECT 661.650 507.750 663.450 513.600 ;
        RECT 664.650 507.750 666.450 513.600 ;
        RECT 667.650 507.750 669.450 513.600 ;
        RECT 702.300 507.750 704.100 519.600 ;
        RECT 706.500 507.750 708.300 519.600 ;
        RECT 743.550 513.600 744.750 520.500 ;
        RECT 750.150 519.600 751.350 524.850 ;
        RECT 709.800 507.750 711.600 513.600 ;
        RECT 743.550 507.750 745.350 513.600 ;
        RECT 746.850 507.750 748.650 519.600 ;
        RECT 749.850 507.750 751.650 519.600 ;
        RECT 3.150 491.400 4.950 503.250 ;
        RECT 6.150 497.400 7.950 503.250 ;
        RECT 11.250 497.400 13.050 503.250 ;
        RECT 16.050 497.400 17.850 503.250 ;
        RECT 11.550 496.500 12.750 497.400 ;
        RECT 19.050 496.500 20.850 503.250 ;
        RECT 22.950 497.400 24.750 503.250 ;
        RECT 27.150 497.400 28.950 503.250 ;
        RECT 31.650 500.400 33.450 503.250 ;
        RECT 7.950 494.400 12.750 496.500 ;
        RECT 15.150 494.700 22.050 496.500 ;
        RECT 27.150 495.300 31.050 497.400 ;
        RECT 11.550 493.500 12.750 494.400 ;
        RECT 24.450 493.800 26.250 494.400 ;
        RECT 11.550 492.300 19.050 493.500 ;
        RECT 17.250 491.700 19.050 492.300 ;
        RECT 19.950 492.900 26.250 493.800 ;
        RECT 3.150 490.800 14.250 491.400 ;
        RECT 19.950 490.800 20.850 492.900 ;
        RECT 24.450 492.600 26.250 492.900 ;
        RECT 27.150 492.600 29.850 494.400 ;
        RECT 27.150 491.700 28.050 492.600 ;
        RECT 3.150 490.200 20.850 490.800 ;
        RECT 3.150 477.600 4.050 490.200 ;
        RECT 12.450 489.900 20.850 490.200 ;
        RECT 22.050 490.800 28.050 491.700 ;
        RECT 28.950 490.800 31.050 491.700 ;
        RECT 34.650 491.400 36.450 503.250 ;
        RECT 66.300 491.400 68.100 503.250 ;
        RECT 70.500 491.400 72.300 503.250 ;
        RECT 73.800 497.400 75.600 503.250 ;
        RECT 108.300 491.400 110.100 503.250 ;
        RECT 112.500 491.400 114.300 503.250 ;
        RECT 115.800 497.400 117.600 503.250 ;
        RECT 154.650 497.400 156.450 503.250 ;
        RECT 157.650 497.400 159.450 503.250 ;
        RECT 160.650 497.400 162.450 503.250 ;
        RECT 12.450 489.600 14.250 489.900 ;
        RECT 22.050 486.150 22.950 490.800 ;
        RECT 28.950 489.600 33.150 490.800 ;
        RECT 32.250 487.800 34.050 489.600 ;
        RECT 13.950 485.100 16.050 486.150 ;
        RECT 5.100 483.150 6.900 484.950 ;
        RECT 8.100 484.050 16.050 485.100 ;
        RECT 19.950 484.050 22.950 486.150 ;
        RECT 8.100 483.300 9.900 484.050 ;
        RECT 6.000 482.400 6.900 483.150 ;
        RECT 11.100 482.400 12.900 483.000 ;
        RECT 6.000 481.200 12.900 482.400 ;
        RECT 11.850 480.000 12.900 481.200 ;
        RECT 22.050 480.000 22.950 484.050 ;
        RECT 31.950 483.750 34.050 484.050 ;
        RECT 30.150 481.950 34.050 483.750 ;
        RECT 35.250 481.950 36.450 491.400 ;
        RECT 65.100 486.150 66.900 487.950 ;
        RECT 70.950 486.150 72.150 491.400 ;
        RECT 73.950 489.150 75.750 490.950 ;
        RECT 73.950 487.050 76.050 489.150 ;
        RECT 107.100 486.150 108.900 487.950 ;
        RECT 112.950 486.150 114.150 491.400 ;
        RECT 115.950 489.150 117.750 490.950 ;
        RECT 158.250 489.150 159.450 497.400 ;
        RECT 165.150 491.400 166.950 503.250 ;
        RECT 168.150 497.400 169.950 503.250 ;
        RECT 173.250 497.400 175.050 503.250 ;
        RECT 178.050 497.400 179.850 503.250 ;
        RECT 173.550 496.500 174.750 497.400 ;
        RECT 181.050 496.500 182.850 503.250 ;
        RECT 184.950 497.400 186.750 503.250 ;
        RECT 189.150 497.400 190.950 503.250 ;
        RECT 193.650 500.400 195.450 503.250 ;
        RECT 169.950 494.400 174.750 496.500 ;
        RECT 177.150 494.700 184.050 496.500 ;
        RECT 189.150 495.300 193.050 497.400 ;
        RECT 173.550 493.500 174.750 494.400 ;
        RECT 186.450 493.800 188.250 494.400 ;
        RECT 173.550 492.300 181.050 493.500 ;
        RECT 179.250 491.700 181.050 492.300 ;
        RECT 181.950 492.900 188.250 493.800 ;
        RECT 165.150 490.800 176.250 491.400 ;
        RECT 181.950 490.800 182.850 492.900 ;
        RECT 186.450 492.600 188.250 492.900 ;
        RECT 189.150 492.600 191.850 494.400 ;
        RECT 189.150 491.700 190.050 492.600 ;
        RECT 165.150 490.200 182.850 490.800 ;
        RECT 115.950 487.050 118.050 489.150 ;
        RECT 64.950 484.050 67.050 486.150 ;
        RECT 67.950 482.850 70.050 484.950 ;
        RECT 70.950 484.050 73.050 486.150 ;
        RECT 106.950 484.050 109.050 486.150 ;
        RECT 11.850 479.100 22.950 480.000 ;
        RECT 31.950 479.850 36.450 481.950 ;
        RECT 68.100 481.050 69.900 482.850 ;
        RECT 71.850 480.750 73.050 484.050 ;
        RECT 109.950 482.850 112.050 484.950 ;
        RECT 112.950 484.050 115.050 486.150 ;
        RECT 154.950 485.850 157.050 487.950 ;
        RECT 157.950 487.050 160.050 489.150 ;
        RECT 155.100 484.050 156.900 485.850 ;
        RECT 110.100 481.050 111.900 482.850 ;
        RECT 113.850 480.750 115.050 484.050 ;
        RECT 11.850 478.200 12.900 479.100 ;
        RECT 22.050 478.800 22.950 479.100 ;
        RECT 3.150 471.750 4.950 477.600 ;
        RECT 7.950 475.500 10.050 477.600 ;
        RECT 11.550 476.400 13.350 478.200 ;
        RECT 14.850 477.450 16.650 478.200 ;
        RECT 14.850 476.400 19.800 477.450 ;
        RECT 22.050 477.000 23.850 478.800 ;
        RECT 35.250 477.600 36.450 479.850 ;
        RECT 72.000 479.700 75.750 480.750 ;
        RECT 114.000 479.700 117.750 480.750 ;
        RECT 158.250 479.700 159.450 487.050 ;
        RECT 160.950 485.850 163.050 487.950 ;
        RECT 161.100 484.050 162.900 485.850 ;
        RECT 28.950 476.700 31.050 477.600 ;
        RECT 9.000 474.600 10.050 475.500 ;
        RECT 18.750 474.600 19.800 476.400 ;
        RECT 27.300 475.500 31.050 476.700 ;
        RECT 27.300 474.600 28.350 475.500 ;
        RECT 6.150 471.750 7.950 474.600 ;
        RECT 9.000 473.700 12.750 474.600 ;
        RECT 10.950 471.750 12.750 473.700 ;
        RECT 15.450 471.750 17.250 474.600 ;
        RECT 18.750 471.750 20.550 474.600 ;
        RECT 22.650 471.750 24.450 474.600 ;
        RECT 26.850 471.750 28.650 474.600 ;
        RECT 31.350 471.750 33.150 474.600 ;
        RECT 34.650 471.750 36.450 477.600 ;
        RECT 65.550 476.700 73.350 478.050 ;
        RECT 65.550 471.750 67.350 476.700 ;
        RECT 68.550 471.750 70.350 475.800 ;
        RECT 71.550 471.750 73.350 476.700 ;
        RECT 74.550 477.600 75.750 479.700 ;
        RECT 74.550 471.750 76.350 477.600 ;
        RECT 107.550 476.700 115.350 478.050 ;
        RECT 107.550 471.750 109.350 476.700 ;
        RECT 110.550 471.750 112.350 475.800 ;
        RECT 113.550 471.750 115.350 476.700 ;
        RECT 116.550 477.600 117.750 479.700 ;
        RECT 155.850 478.800 159.450 479.700 ;
        RECT 116.550 471.750 118.350 477.600 ;
        RECT 155.850 471.750 157.650 478.800 ;
        RECT 165.150 477.600 166.050 490.200 ;
        RECT 174.450 489.900 182.850 490.200 ;
        RECT 184.050 490.800 190.050 491.700 ;
        RECT 190.950 490.800 193.050 491.700 ;
        RECT 196.650 491.400 198.450 503.250 ;
        RECT 228.300 491.400 230.100 503.250 ;
        RECT 232.500 491.400 234.300 503.250 ;
        RECT 235.800 497.400 237.600 503.250 ;
        RECT 269.550 497.400 271.350 503.250 ;
        RECT 272.550 497.400 274.350 503.250 ;
        RECT 174.450 489.600 176.250 489.900 ;
        RECT 184.050 486.150 184.950 490.800 ;
        RECT 190.950 489.600 195.150 490.800 ;
        RECT 194.250 487.800 196.050 489.600 ;
        RECT 175.950 485.100 178.050 486.150 ;
        RECT 167.100 483.150 168.900 484.950 ;
        RECT 170.100 484.050 178.050 485.100 ;
        RECT 181.950 484.050 184.950 486.150 ;
        RECT 170.100 483.300 171.900 484.050 ;
        RECT 168.000 482.400 168.900 483.150 ;
        RECT 173.100 482.400 174.900 483.000 ;
        RECT 168.000 481.200 174.900 482.400 ;
        RECT 173.850 480.000 174.900 481.200 ;
        RECT 184.050 480.000 184.950 484.050 ;
        RECT 193.950 483.750 196.050 484.050 ;
        RECT 192.150 481.950 196.050 483.750 ;
        RECT 197.250 481.950 198.450 491.400 ;
        RECT 227.100 486.150 228.900 487.950 ;
        RECT 232.950 486.150 234.150 491.400 ;
        RECT 235.950 489.150 237.750 490.950 ;
        RECT 235.950 487.050 238.050 489.150 ;
        RECT 269.100 486.150 270.900 487.950 ;
        RECT 226.950 484.050 229.050 486.150 ;
        RECT 229.950 482.850 232.050 484.950 ;
        RECT 232.950 484.050 235.050 486.150 ;
        RECT 268.950 484.050 271.050 486.150 ;
        RECT 173.850 479.100 184.950 480.000 ;
        RECT 193.950 479.850 198.450 481.950 ;
        RECT 230.100 481.050 231.900 482.850 ;
        RECT 233.850 480.750 235.050 484.050 ;
        RECT 173.850 478.200 174.900 479.100 ;
        RECT 184.050 478.800 184.950 479.100 ;
        RECT 160.350 471.750 162.150 477.600 ;
        RECT 165.150 471.750 166.950 477.600 ;
        RECT 169.950 475.500 172.050 477.600 ;
        RECT 173.550 476.400 175.350 478.200 ;
        RECT 176.850 477.450 178.650 478.200 ;
        RECT 176.850 476.400 181.800 477.450 ;
        RECT 184.050 477.000 185.850 478.800 ;
        RECT 197.250 477.600 198.450 479.850 ;
        RECT 234.000 479.700 237.750 480.750 ;
        RECT 272.700 480.300 273.900 497.400 ;
        RECT 276.150 491.400 277.950 503.250 ;
        RECT 279.150 491.400 280.950 503.250 ;
        RECT 285.150 491.400 286.950 503.250 ;
        RECT 288.150 497.400 289.950 503.250 ;
        RECT 293.250 497.400 295.050 503.250 ;
        RECT 298.050 497.400 299.850 503.250 ;
        RECT 293.550 496.500 294.750 497.400 ;
        RECT 301.050 496.500 302.850 503.250 ;
        RECT 304.950 497.400 306.750 503.250 ;
        RECT 309.150 497.400 310.950 503.250 ;
        RECT 313.650 500.400 315.450 503.250 ;
        RECT 289.950 494.400 294.750 496.500 ;
        RECT 297.150 494.700 304.050 496.500 ;
        RECT 309.150 495.300 313.050 497.400 ;
        RECT 293.550 493.500 294.750 494.400 ;
        RECT 306.450 493.800 308.250 494.400 ;
        RECT 293.550 492.300 301.050 493.500 ;
        RECT 299.250 491.700 301.050 492.300 ;
        RECT 301.950 492.900 308.250 493.800 ;
        RECT 274.950 485.850 277.050 487.950 ;
        RECT 279.150 486.150 280.350 491.400 ;
        RECT 275.100 484.050 276.900 485.850 ;
        RECT 277.950 484.050 280.350 486.150 ;
        RECT 190.950 476.700 193.050 477.600 ;
        RECT 171.000 474.600 172.050 475.500 ;
        RECT 180.750 474.600 181.800 476.400 ;
        RECT 189.300 475.500 193.050 476.700 ;
        RECT 189.300 474.600 190.350 475.500 ;
        RECT 168.150 471.750 169.950 474.600 ;
        RECT 171.000 473.700 174.750 474.600 ;
        RECT 172.950 471.750 174.750 473.700 ;
        RECT 177.450 471.750 179.250 474.600 ;
        RECT 180.750 471.750 182.550 474.600 ;
        RECT 184.650 471.750 186.450 474.600 ;
        RECT 188.850 471.750 190.650 474.600 ;
        RECT 193.350 471.750 195.150 474.600 ;
        RECT 196.650 471.750 198.450 477.600 ;
        RECT 227.550 476.700 235.350 478.050 ;
        RECT 227.550 471.750 229.350 476.700 ;
        RECT 230.550 471.750 232.350 475.800 ;
        RECT 233.550 471.750 235.350 476.700 ;
        RECT 236.550 477.600 237.750 479.700 ;
        RECT 269.550 479.100 277.050 480.300 ;
        RECT 236.550 471.750 238.350 477.600 ;
        RECT 269.550 471.750 271.350 479.100 ;
        RECT 275.250 478.500 277.050 479.100 ;
        RECT 279.150 477.600 280.350 484.050 ;
        RECT 274.050 471.750 275.850 477.600 ;
        RECT 277.050 476.100 280.350 477.600 ;
        RECT 285.150 490.800 296.250 491.400 ;
        RECT 301.950 490.800 302.850 492.900 ;
        RECT 306.450 492.600 308.250 492.900 ;
        RECT 309.150 492.600 311.850 494.400 ;
        RECT 309.150 491.700 310.050 492.600 ;
        RECT 285.150 490.200 302.850 490.800 ;
        RECT 285.150 477.600 286.050 490.200 ;
        RECT 294.450 489.900 302.850 490.200 ;
        RECT 304.050 490.800 310.050 491.700 ;
        RECT 310.950 490.800 313.050 491.700 ;
        RECT 316.650 491.400 318.450 503.250 ;
        RECT 353.400 497.400 355.200 503.250 ;
        RECT 356.700 491.400 358.500 503.250 ;
        RECT 360.900 491.400 362.700 503.250 ;
        RECT 392.550 491.400 394.350 503.250 ;
        RECT 294.450 489.600 296.250 489.900 ;
        RECT 304.050 486.150 304.950 490.800 ;
        RECT 310.950 489.600 315.150 490.800 ;
        RECT 314.250 487.800 316.050 489.600 ;
        RECT 295.950 485.100 298.050 486.150 ;
        RECT 287.100 483.150 288.900 484.950 ;
        RECT 290.100 484.050 298.050 485.100 ;
        RECT 301.950 484.050 304.950 486.150 ;
        RECT 290.100 483.300 291.900 484.050 ;
        RECT 288.000 482.400 288.900 483.150 ;
        RECT 293.100 482.400 294.900 483.000 ;
        RECT 288.000 481.200 294.900 482.400 ;
        RECT 293.850 480.000 294.900 481.200 ;
        RECT 304.050 480.000 304.950 484.050 ;
        RECT 313.950 483.750 316.050 484.050 ;
        RECT 312.150 481.950 316.050 483.750 ;
        RECT 317.250 481.950 318.450 491.400 ;
        RECT 353.250 489.150 355.050 490.950 ;
        RECT 352.950 487.050 355.050 489.150 ;
        RECT 356.850 486.150 358.050 491.400 ;
        RECT 395.550 490.500 397.350 503.250 ;
        RECT 398.550 491.400 400.350 503.250 ;
        RECT 401.550 490.500 403.350 503.250 ;
        RECT 404.550 491.400 406.350 503.250 ;
        RECT 407.550 490.500 409.350 503.250 ;
        RECT 410.550 491.400 412.350 503.250 ;
        RECT 413.550 490.500 415.350 503.250 ;
        RECT 416.550 491.400 418.350 503.250 ;
        RECT 454.350 491.400 456.150 503.250 ;
        RECT 457.350 491.400 459.150 503.250 ;
        RECT 460.650 497.400 462.450 503.250 ;
        RECT 496.650 497.400 498.450 503.250 ;
        RECT 499.650 497.400 501.450 503.250 ;
        RECT 502.650 497.400 504.450 503.250 ;
        RECT 538.650 497.400 540.450 503.250 ;
        RECT 541.650 497.400 543.450 503.250 ;
        RECT 544.650 497.400 546.450 503.250 ;
        RECT 395.550 489.300 399.450 490.500 ;
        RECT 401.550 489.300 405.300 490.500 ;
        RECT 407.550 489.300 411.300 490.500 ;
        RECT 413.550 489.300 416.250 490.500 ;
        RECT 362.100 486.150 363.900 487.950 ;
        RECT 293.850 479.100 304.950 480.000 ;
        RECT 313.950 479.850 318.450 481.950 ;
        RECT 355.950 484.050 358.050 486.150 ;
        RECT 355.950 480.750 357.150 484.050 ;
        RECT 358.950 482.850 361.050 484.950 ;
        RECT 361.950 484.050 364.050 486.150 ;
        RECT 394.950 482.850 397.050 484.950 ;
        RECT 359.100 481.050 360.900 482.850 ;
        RECT 395.100 481.050 396.900 482.850 ;
        RECT 398.250 482.400 399.450 489.300 ;
        RECT 404.100 482.400 405.300 489.300 ;
        RECT 410.100 482.400 411.300 489.300 ;
        RECT 415.200 484.950 416.250 489.300 ;
        RECT 454.650 486.150 455.850 491.400 ;
        RECT 461.250 490.500 462.450 497.400 ;
        RECT 456.750 489.600 462.450 490.500 ;
        RECT 456.750 488.700 459.000 489.600 ;
        RECT 500.250 489.150 501.450 497.400 ;
        RECT 542.250 489.150 543.450 497.400 ;
        RECT 549.150 491.400 550.950 503.250 ;
        RECT 552.150 497.400 553.950 503.250 ;
        RECT 557.250 497.400 559.050 503.250 ;
        RECT 562.050 497.400 563.850 503.250 ;
        RECT 557.550 496.500 558.750 497.400 ;
        RECT 565.050 496.500 566.850 503.250 ;
        RECT 568.950 497.400 570.750 503.250 ;
        RECT 573.150 497.400 574.950 503.250 ;
        RECT 577.650 500.400 579.450 503.250 ;
        RECT 553.950 494.400 558.750 496.500 ;
        RECT 561.150 494.700 568.050 496.500 ;
        RECT 573.150 495.300 577.050 497.400 ;
        RECT 557.550 493.500 558.750 494.400 ;
        RECT 570.450 493.800 572.250 494.400 ;
        RECT 557.550 492.300 565.050 493.500 ;
        RECT 563.250 491.700 565.050 492.300 ;
        RECT 565.950 492.900 572.250 493.800 ;
        RECT 549.150 490.800 560.250 491.400 ;
        RECT 565.950 490.800 566.850 492.900 ;
        RECT 570.450 492.600 572.250 492.900 ;
        RECT 573.150 492.600 575.850 494.400 ;
        RECT 573.150 491.700 574.050 492.600 ;
        RECT 549.150 490.200 566.850 490.800 ;
        RECT 415.200 482.850 418.050 484.950 ;
        RECT 454.650 484.050 457.050 486.150 ;
        RECT 293.850 478.200 294.900 479.100 ;
        RECT 304.050 478.800 304.950 479.100 ;
        RECT 277.050 471.750 278.850 476.100 ;
        RECT 285.150 471.750 286.950 477.600 ;
        RECT 289.950 475.500 292.050 477.600 ;
        RECT 293.550 476.400 295.350 478.200 ;
        RECT 296.850 477.450 298.650 478.200 ;
        RECT 296.850 476.400 301.800 477.450 ;
        RECT 304.050 477.000 305.850 478.800 ;
        RECT 317.250 477.600 318.450 479.850 ;
        RECT 353.250 479.700 357.000 480.750 ;
        RECT 398.250 480.600 402.300 482.400 ;
        RECT 404.100 480.600 408.300 482.400 ;
        RECT 410.100 480.600 414.300 482.400 ;
        RECT 398.250 479.700 399.450 480.600 ;
        RECT 404.100 479.700 405.300 480.600 ;
        RECT 410.100 479.700 411.300 480.600 ;
        RECT 415.200 479.700 416.250 482.850 ;
        RECT 353.250 477.600 354.450 479.700 ;
        RECT 395.400 478.500 399.450 479.700 ;
        RECT 401.550 478.500 405.300 479.700 ;
        RECT 407.400 478.500 411.300 479.700 ;
        RECT 413.400 478.650 416.250 479.700 ;
        RECT 413.400 478.500 416.100 478.650 ;
        RECT 310.950 476.700 313.050 477.600 ;
        RECT 291.000 474.600 292.050 475.500 ;
        RECT 300.750 474.600 301.800 476.400 ;
        RECT 309.300 475.500 313.050 476.700 ;
        RECT 309.300 474.600 310.350 475.500 ;
        RECT 288.150 471.750 289.950 474.600 ;
        RECT 291.000 473.700 294.750 474.600 ;
        RECT 292.950 471.750 294.750 473.700 ;
        RECT 297.450 471.750 299.250 474.600 ;
        RECT 300.750 471.750 302.550 474.600 ;
        RECT 304.650 471.750 306.450 474.600 ;
        RECT 308.850 471.750 310.650 474.600 ;
        RECT 313.350 471.750 315.150 474.600 ;
        RECT 316.650 471.750 318.450 477.600 ;
        RECT 352.650 471.750 354.450 477.600 ;
        RECT 355.650 476.700 363.450 478.050 ;
        RECT 395.400 477.600 397.200 478.500 ;
        RECT 355.650 471.750 357.450 476.700 ;
        RECT 358.650 471.750 360.450 475.800 ;
        RECT 361.650 471.750 363.450 476.700 ;
        RECT 392.550 471.750 394.350 477.600 ;
        RECT 395.550 471.750 397.350 477.600 ;
        RECT 398.550 471.750 400.350 477.600 ;
        RECT 401.550 471.750 403.350 478.500 ;
        RECT 407.400 477.600 409.200 478.500 ;
        RECT 413.400 477.600 415.200 478.500 ;
        RECT 454.650 477.600 455.850 484.050 ;
        RECT 457.950 480.300 459.000 488.700 ;
        RECT 461.100 486.150 462.900 487.950 ;
        RECT 460.950 484.050 463.050 486.150 ;
        RECT 496.950 485.850 499.050 487.950 ;
        RECT 499.950 487.050 502.050 489.150 ;
        RECT 497.100 484.050 498.900 485.850 ;
        RECT 456.750 479.400 459.000 480.300 ;
        RECT 500.250 479.700 501.450 487.050 ;
        RECT 502.950 485.850 505.050 487.950 ;
        RECT 538.950 485.850 541.050 487.950 ;
        RECT 541.950 487.050 544.050 489.150 ;
        RECT 503.100 484.050 504.900 485.850 ;
        RECT 539.100 484.050 540.900 485.850 ;
        RECT 542.250 479.700 543.450 487.050 ;
        RECT 544.950 485.850 547.050 487.950 ;
        RECT 545.100 484.050 546.900 485.850 ;
        RECT 456.750 478.500 461.850 479.400 ;
        RECT 404.550 471.750 406.350 477.600 ;
        RECT 407.550 471.750 409.350 477.600 ;
        RECT 410.550 471.750 412.350 477.600 ;
        RECT 413.550 471.750 415.350 477.600 ;
        RECT 416.550 471.750 418.350 477.600 ;
        RECT 454.350 471.750 456.150 477.600 ;
        RECT 457.350 471.750 459.150 477.600 ;
        RECT 460.650 474.600 461.850 478.500 ;
        RECT 497.850 478.800 501.450 479.700 ;
        RECT 539.850 478.800 543.450 479.700 ;
        RECT 460.650 471.750 462.450 474.600 ;
        RECT 497.850 471.750 499.650 478.800 ;
        RECT 502.350 471.750 504.150 477.600 ;
        RECT 539.850 471.750 541.650 478.800 ;
        RECT 549.150 477.600 550.050 490.200 ;
        RECT 558.450 489.900 566.850 490.200 ;
        RECT 568.050 490.800 574.050 491.700 ;
        RECT 574.950 490.800 577.050 491.700 ;
        RECT 580.650 491.400 582.450 503.250 ;
        RECT 612.300 491.400 614.100 503.250 ;
        RECT 616.500 491.400 618.300 503.250 ;
        RECT 619.800 497.400 621.600 503.250 ;
        RECT 658.650 497.400 660.450 503.250 ;
        RECT 661.650 497.400 663.450 503.250 ;
        RECT 664.650 497.400 666.450 503.250 ;
        RECT 698.550 497.400 700.350 503.250 ;
        RECT 558.450 489.600 560.250 489.900 ;
        RECT 568.050 486.150 568.950 490.800 ;
        RECT 574.950 489.600 579.150 490.800 ;
        RECT 578.250 487.800 580.050 489.600 ;
        RECT 559.950 485.100 562.050 486.150 ;
        RECT 551.100 483.150 552.900 484.950 ;
        RECT 554.100 484.050 562.050 485.100 ;
        RECT 565.950 484.050 568.950 486.150 ;
        RECT 554.100 483.300 555.900 484.050 ;
        RECT 552.000 482.400 552.900 483.150 ;
        RECT 557.100 482.400 558.900 483.000 ;
        RECT 552.000 481.200 558.900 482.400 ;
        RECT 557.850 480.000 558.900 481.200 ;
        RECT 568.050 480.000 568.950 484.050 ;
        RECT 577.950 483.750 580.050 484.050 ;
        RECT 576.150 481.950 580.050 483.750 ;
        RECT 581.250 481.950 582.450 491.400 ;
        RECT 611.100 486.150 612.900 487.950 ;
        RECT 616.950 486.150 618.150 491.400 ;
        RECT 619.950 489.150 621.750 490.950 ;
        RECT 662.250 489.150 663.450 497.400 ;
        RECT 698.550 490.500 699.750 497.400 ;
        RECT 701.850 491.400 703.650 503.250 ;
        RECT 704.850 491.400 706.650 503.250 ;
        RECT 740.550 497.400 742.350 503.250 ;
        RECT 698.550 489.600 704.250 490.500 ;
        RECT 619.950 487.050 622.050 489.150 ;
        RECT 610.950 484.050 613.050 486.150 ;
        RECT 613.950 482.850 616.050 484.950 ;
        RECT 616.950 484.050 619.050 486.150 ;
        RECT 658.950 485.850 661.050 487.950 ;
        RECT 661.950 487.050 664.050 489.150 ;
        RECT 702.000 488.700 704.250 489.600 ;
        RECT 659.100 484.050 660.900 485.850 ;
        RECT 557.850 479.100 568.950 480.000 ;
        RECT 577.950 479.850 582.450 481.950 ;
        RECT 614.100 481.050 615.900 482.850 ;
        RECT 617.850 480.750 619.050 484.050 ;
        RECT 557.850 478.200 558.900 479.100 ;
        RECT 568.050 478.800 568.950 479.100 ;
        RECT 544.350 471.750 546.150 477.600 ;
        RECT 549.150 471.750 550.950 477.600 ;
        RECT 553.950 475.500 556.050 477.600 ;
        RECT 557.550 476.400 559.350 478.200 ;
        RECT 560.850 477.450 562.650 478.200 ;
        RECT 560.850 476.400 565.800 477.450 ;
        RECT 568.050 477.000 569.850 478.800 ;
        RECT 581.250 477.600 582.450 479.850 ;
        RECT 618.000 479.700 621.750 480.750 ;
        RECT 662.250 479.700 663.450 487.050 ;
        RECT 664.950 485.850 667.050 487.950 ;
        RECT 698.100 486.150 699.900 487.950 ;
        RECT 665.100 484.050 666.900 485.850 ;
        RECT 697.950 484.050 700.050 486.150 ;
        RECT 574.950 476.700 577.050 477.600 ;
        RECT 555.000 474.600 556.050 475.500 ;
        RECT 564.750 474.600 565.800 476.400 ;
        RECT 573.300 475.500 577.050 476.700 ;
        RECT 573.300 474.600 574.350 475.500 ;
        RECT 552.150 471.750 553.950 474.600 ;
        RECT 555.000 473.700 558.750 474.600 ;
        RECT 556.950 471.750 558.750 473.700 ;
        RECT 561.450 471.750 563.250 474.600 ;
        RECT 564.750 471.750 566.550 474.600 ;
        RECT 568.650 471.750 570.450 474.600 ;
        RECT 572.850 471.750 574.650 474.600 ;
        RECT 577.350 471.750 579.150 474.600 ;
        RECT 580.650 471.750 582.450 477.600 ;
        RECT 611.550 476.700 619.350 478.050 ;
        RECT 611.550 471.750 613.350 476.700 ;
        RECT 614.550 471.750 616.350 475.800 ;
        RECT 617.550 471.750 619.350 476.700 ;
        RECT 620.550 477.600 621.750 479.700 ;
        RECT 659.850 478.800 663.450 479.700 ;
        RECT 702.000 480.300 703.050 488.700 ;
        RECT 705.150 486.150 706.350 491.400 ;
        RECT 740.550 490.500 741.750 497.400 ;
        RECT 743.850 491.400 745.650 503.250 ;
        RECT 746.850 491.400 748.650 503.250 ;
        RECT 740.550 489.600 746.250 490.500 ;
        RECT 744.000 488.700 746.250 489.600 ;
        RECT 740.100 486.150 741.900 487.950 ;
        RECT 703.950 484.050 706.350 486.150 ;
        RECT 739.950 484.050 742.050 486.150 ;
        RECT 702.000 479.400 704.250 480.300 ;
        RECT 620.550 471.750 622.350 477.600 ;
        RECT 659.850 471.750 661.650 478.800 ;
        RECT 699.150 478.500 704.250 479.400 ;
        RECT 664.350 471.750 666.150 477.600 ;
        RECT 699.150 474.600 700.350 478.500 ;
        RECT 705.150 477.600 706.350 484.050 ;
        RECT 744.000 480.300 745.050 488.700 ;
        RECT 747.150 486.150 748.350 491.400 ;
        RECT 745.950 484.050 748.350 486.150 ;
        RECT 744.000 479.400 746.250 480.300 ;
        RECT 741.150 478.500 746.250 479.400 ;
        RECT 698.550 471.750 700.350 474.600 ;
        RECT 701.850 471.750 703.650 477.600 ;
        RECT 704.850 471.750 706.650 477.600 ;
        RECT 741.150 474.600 742.350 478.500 ;
        RECT 747.150 477.600 748.350 484.050 ;
        RECT 740.550 471.750 742.350 474.600 ;
        RECT 743.850 471.750 745.650 477.600 ;
        RECT 746.850 471.750 748.650 477.600 ;
        RECT 32.550 461.400 34.350 467.250 ;
        RECT 35.550 461.400 37.350 467.250 ;
        RECT 38.550 461.400 40.350 467.250 ;
        RECT 35.400 460.500 37.200 461.400 ;
        RECT 41.550 460.500 43.350 467.250 ;
        RECT 44.550 461.400 46.350 467.250 ;
        RECT 47.550 461.400 49.350 467.250 ;
        RECT 50.550 461.400 52.350 467.250 ;
        RECT 53.550 461.400 55.350 467.250 ;
        RECT 56.550 461.400 58.350 467.250 ;
        RECT 94.650 464.400 96.450 467.250 ;
        RECT 97.650 464.400 99.450 467.250 ;
        RECT 47.400 460.500 49.200 461.400 ;
        RECT 53.400 460.500 55.200 461.400 ;
        RECT 35.400 459.300 39.450 460.500 ;
        RECT 41.550 459.300 45.300 460.500 ;
        RECT 47.400 459.300 51.300 460.500 ;
        RECT 53.400 460.350 56.100 460.500 ;
        RECT 53.400 459.300 56.250 460.350 ;
        RECT 38.250 458.400 39.450 459.300 ;
        RECT 44.100 458.400 45.300 459.300 ;
        RECT 50.100 458.400 51.300 459.300 ;
        RECT 35.100 456.150 36.900 457.950 ;
        RECT 38.250 456.600 42.300 458.400 ;
        RECT 44.100 456.600 48.300 458.400 ;
        RECT 50.100 456.600 54.300 458.400 ;
        RECT 34.950 454.050 37.050 456.150 ;
        RECT 38.250 449.700 39.450 456.600 ;
        RECT 44.100 449.700 45.300 456.600 ;
        RECT 50.100 449.700 51.300 456.600 ;
        RECT 55.200 456.150 56.250 459.300 ;
        RECT 95.400 456.150 96.600 464.400 ;
        RECT 131.850 460.200 133.650 467.250 ;
        RECT 136.350 461.400 138.150 467.250 ;
        RECT 170.850 461.400 172.650 467.250 ;
        RECT 175.350 460.200 177.150 467.250 ;
        RECT 214.650 464.400 216.450 467.250 ;
        RECT 217.650 464.400 219.450 467.250 ;
        RECT 131.850 459.300 135.450 460.200 ;
        RECT 55.200 454.050 58.050 456.150 ;
        RECT 94.950 454.050 97.050 456.150 ;
        RECT 97.950 455.850 100.050 457.950 ;
        RECT 98.100 454.050 99.900 455.850 ;
        RECT 55.200 449.700 56.250 454.050 ;
        RECT 35.550 448.500 39.450 449.700 ;
        RECT 41.550 448.500 45.300 449.700 ;
        RECT 47.550 448.500 51.300 449.700 ;
        RECT 53.550 448.500 56.250 449.700 ;
        RECT 32.550 435.750 34.350 447.600 ;
        RECT 35.550 435.750 37.350 448.500 ;
        RECT 38.550 435.750 40.350 447.600 ;
        RECT 41.550 435.750 43.350 448.500 ;
        RECT 44.550 435.750 46.350 447.600 ;
        RECT 47.550 435.750 49.350 448.500 ;
        RECT 50.550 435.750 52.350 447.600 ;
        RECT 53.550 435.750 55.350 448.500 ;
        RECT 56.550 435.750 58.350 447.600 ;
        RECT 95.400 441.600 96.600 454.050 ;
        RECT 131.100 453.150 132.900 454.950 ;
        RECT 130.950 451.050 133.050 453.150 ;
        RECT 134.250 451.950 135.450 459.300 ;
        RECT 173.550 459.300 177.150 460.200 ;
        RECT 137.100 453.150 138.900 454.950 ;
        RECT 170.100 453.150 171.900 454.950 ;
        RECT 133.950 449.850 136.050 451.950 ;
        RECT 136.950 451.050 139.050 453.150 ;
        RECT 169.950 451.050 172.050 453.150 ;
        RECT 173.550 451.950 174.750 459.300 ;
        RECT 215.400 456.150 216.600 464.400 ;
        RECT 251.850 461.400 253.650 467.250 ;
        RECT 256.350 460.200 258.150 467.250 ;
        RECT 295.650 461.400 297.450 467.250 ;
        RECT 254.550 459.300 258.150 460.200 ;
        RECT 296.250 459.300 297.450 461.400 ;
        RECT 298.650 462.300 300.450 467.250 ;
        RECT 301.650 463.200 303.450 467.250 ;
        RECT 304.650 462.300 306.450 467.250 ;
        RECT 340.650 464.400 342.450 467.250 ;
        RECT 343.650 464.400 345.450 467.250 ;
        RECT 346.650 464.400 348.450 467.250 ;
        RECT 298.650 460.950 306.450 462.300 ;
        RECT 176.100 453.150 177.900 454.950 ;
        RECT 214.950 454.050 217.050 456.150 ;
        RECT 217.950 455.850 220.050 457.950 ;
        RECT 218.100 454.050 219.900 455.850 ;
        RECT 172.950 449.850 175.050 451.950 ;
        RECT 175.950 451.050 178.050 453.150 ;
        RECT 134.250 441.600 135.450 449.850 ;
        RECT 173.550 441.600 174.750 449.850 ;
        RECT 215.400 441.600 216.600 454.050 ;
        RECT 251.100 453.150 252.900 454.950 ;
        RECT 250.950 451.050 253.050 453.150 ;
        RECT 254.550 451.950 255.750 459.300 ;
        RECT 296.250 458.250 300.000 459.300 ;
        RECT 298.950 454.950 300.150 458.250 ;
        RECT 343.950 457.950 345.000 464.400 ;
        RECT 351.150 461.400 352.950 467.250 ;
        RECT 354.150 464.400 355.950 467.250 ;
        RECT 358.950 465.300 360.750 467.250 ;
        RECT 357.000 464.400 360.750 465.300 ;
        RECT 363.450 464.400 365.250 467.250 ;
        RECT 366.750 464.400 368.550 467.250 ;
        RECT 370.650 464.400 372.450 467.250 ;
        RECT 374.850 464.400 376.650 467.250 ;
        RECT 379.350 464.400 381.150 467.250 ;
        RECT 357.000 463.500 358.050 464.400 ;
        RECT 355.950 461.400 358.050 463.500 ;
        RECT 366.750 462.600 367.800 464.400 ;
        RECT 302.100 456.150 303.900 457.950 ;
        RECT 257.100 453.150 258.900 454.950 ;
        RECT 253.950 449.850 256.050 451.950 ;
        RECT 256.950 451.050 259.050 453.150 ;
        RECT 298.950 452.850 301.050 454.950 ;
        RECT 301.950 454.050 304.050 456.150 ;
        RECT 343.950 455.850 346.050 457.950 ;
        RECT 304.950 452.850 307.050 454.950 ;
        RECT 340.950 452.850 343.050 454.950 ;
        RECT 295.950 449.850 298.050 451.950 ;
        RECT 254.550 441.600 255.750 449.850 ;
        RECT 296.250 448.050 298.050 449.850 ;
        RECT 299.850 447.600 301.050 452.850 ;
        RECT 305.100 451.050 306.900 452.850 ;
        RECT 341.100 451.050 342.900 452.850 ;
        RECT 343.950 448.650 345.000 455.850 ;
        RECT 346.950 452.850 349.050 454.950 ;
        RECT 347.100 451.050 348.900 452.850 ;
        RECT 342.450 447.600 345.000 448.650 ;
        RECT 351.150 448.800 352.050 461.400 ;
        RECT 359.550 460.800 361.350 462.600 ;
        RECT 362.850 461.550 367.800 462.600 ;
        RECT 375.300 463.500 376.350 464.400 ;
        RECT 375.300 462.300 379.050 463.500 ;
        RECT 362.850 460.800 364.650 461.550 ;
        RECT 359.850 459.900 360.900 460.800 ;
        RECT 370.050 460.200 371.850 462.000 ;
        RECT 376.950 461.400 379.050 462.300 ;
        RECT 382.650 461.400 384.450 467.250 ;
        RECT 413.850 461.400 415.650 467.250 ;
        RECT 370.050 459.900 370.950 460.200 ;
        RECT 359.850 459.000 370.950 459.900 ;
        RECT 383.250 459.150 384.450 461.400 ;
        RECT 418.350 460.200 420.150 467.250 ;
        RECT 455.550 464.400 457.350 467.250 ;
        RECT 359.850 457.800 360.900 459.000 ;
        RECT 354.000 456.600 360.900 457.800 ;
        RECT 354.000 455.850 354.900 456.600 ;
        RECT 359.100 456.000 360.900 456.600 ;
        RECT 353.100 454.050 354.900 455.850 ;
        RECT 356.100 454.950 357.900 455.700 ;
        RECT 370.050 454.950 370.950 459.000 ;
        RECT 379.950 457.050 384.450 459.150 ;
        RECT 378.150 455.250 382.050 457.050 ;
        RECT 379.950 454.950 382.050 455.250 ;
        RECT 356.100 453.900 364.050 454.950 ;
        RECT 361.950 452.850 364.050 453.900 ;
        RECT 367.950 452.850 370.950 454.950 ;
        RECT 360.450 449.100 362.250 449.400 ;
        RECT 360.450 448.800 368.850 449.100 ;
        RECT 351.150 448.200 368.850 448.800 ;
        RECT 351.150 447.600 362.250 448.200 ;
        RECT 94.650 435.750 96.450 441.600 ;
        RECT 97.650 435.750 99.450 441.600 ;
        RECT 130.650 435.750 132.450 441.600 ;
        RECT 133.650 435.750 135.450 441.600 ;
        RECT 136.650 435.750 138.450 441.600 ;
        RECT 170.550 435.750 172.350 441.600 ;
        RECT 173.550 435.750 175.350 441.600 ;
        RECT 176.550 435.750 178.350 441.600 ;
        RECT 214.650 435.750 216.450 441.600 ;
        RECT 217.650 435.750 219.450 441.600 ;
        RECT 251.550 435.750 253.350 441.600 ;
        RECT 254.550 435.750 256.350 441.600 ;
        RECT 257.550 435.750 259.350 441.600 ;
        RECT 296.400 435.750 298.200 441.600 ;
        RECT 299.700 435.750 301.500 447.600 ;
        RECT 303.900 435.750 305.700 447.600 ;
        RECT 342.450 435.750 344.250 447.600 ;
        RECT 346.650 435.750 348.450 447.600 ;
        RECT 351.150 435.750 352.950 447.600 ;
        RECT 365.250 446.700 367.050 447.300 ;
        RECT 359.550 445.500 367.050 446.700 ;
        RECT 367.950 446.100 368.850 448.200 ;
        RECT 370.050 448.200 370.950 452.850 ;
        RECT 380.250 449.400 382.050 451.200 ;
        RECT 376.950 448.200 381.150 449.400 ;
        RECT 370.050 447.300 376.050 448.200 ;
        RECT 376.950 447.300 379.050 448.200 ;
        RECT 383.250 447.600 384.450 457.050 ;
        RECT 416.550 459.300 420.150 460.200 ;
        RECT 456.150 460.500 457.350 464.400 ;
        RECT 458.850 461.400 460.650 467.250 ;
        RECT 461.850 461.400 463.650 467.250 ;
        RECT 496.350 461.400 498.150 467.250 ;
        RECT 499.350 461.400 501.150 467.250 ;
        RECT 502.650 464.400 504.450 467.250 ;
        RECT 456.150 459.600 461.250 460.500 ;
        RECT 413.100 453.150 414.900 454.950 ;
        RECT 412.950 451.050 415.050 453.150 ;
        RECT 416.550 451.950 417.750 459.300 ;
        RECT 459.000 458.700 461.250 459.600 ;
        RECT 419.100 453.150 420.900 454.950 ;
        RECT 415.950 449.850 418.050 451.950 ;
        RECT 418.950 451.050 421.050 453.150 ;
        RECT 454.950 452.850 457.050 454.950 ;
        RECT 455.100 451.050 456.900 452.850 ;
        RECT 459.000 450.300 460.050 458.700 ;
        RECT 462.150 454.950 463.350 461.400 ;
        RECT 460.950 452.850 463.350 454.950 ;
        RECT 375.150 446.400 376.050 447.300 ;
        RECT 372.450 446.100 374.250 446.400 ;
        RECT 359.550 444.600 360.750 445.500 ;
        RECT 367.950 445.200 374.250 446.100 ;
        RECT 372.450 444.600 374.250 445.200 ;
        RECT 375.150 444.600 377.850 446.400 ;
        RECT 355.950 442.500 360.750 444.600 ;
        RECT 363.150 442.500 370.050 444.300 ;
        RECT 359.550 441.600 360.750 442.500 ;
        RECT 354.150 435.750 355.950 441.600 ;
        RECT 359.250 435.750 361.050 441.600 ;
        RECT 364.050 435.750 365.850 441.600 ;
        RECT 367.050 435.750 368.850 442.500 ;
        RECT 375.150 441.600 379.050 443.700 ;
        RECT 370.950 435.750 372.750 441.600 ;
        RECT 375.150 435.750 376.950 441.600 ;
        RECT 379.650 435.750 381.450 438.600 ;
        RECT 382.650 435.750 384.450 447.600 ;
        RECT 416.550 441.600 417.750 449.850 ;
        RECT 459.000 449.400 461.250 450.300 ;
        RECT 455.550 448.500 461.250 449.400 ;
        RECT 455.550 441.600 456.750 448.500 ;
        RECT 462.150 447.600 463.350 452.850 ;
        RECT 496.650 454.950 497.850 461.400 ;
        RECT 502.650 460.500 503.850 464.400 ;
        RECT 536.850 461.400 538.650 467.250 ;
        RECT 498.750 459.600 503.850 460.500 ;
        RECT 541.350 460.200 543.150 467.250 ;
        RECT 580.650 461.400 582.450 467.250 ;
        RECT 498.750 458.700 501.000 459.600 ;
        RECT 496.650 452.850 499.050 454.950 ;
        RECT 496.650 447.600 497.850 452.850 ;
        RECT 499.950 450.300 501.000 458.700 ;
        RECT 539.550 459.300 543.150 460.200 ;
        RECT 581.250 459.300 582.450 461.400 ;
        RECT 583.650 462.300 585.450 467.250 ;
        RECT 586.650 463.200 588.450 467.250 ;
        RECT 589.650 462.300 591.450 467.250 ;
        RECT 583.650 460.950 591.450 462.300 ;
        RECT 622.650 461.400 624.450 467.250 ;
        RECT 625.650 461.400 627.450 467.250 ;
        RECT 628.650 461.400 630.450 467.250 ;
        RECT 631.650 461.400 633.450 467.250 ;
        RECT 634.650 461.400 636.450 467.250 ;
        RECT 667.650 464.400 669.450 467.250 ;
        RECT 670.650 464.400 672.450 467.250 ;
        RECT 626.250 460.500 627.450 461.400 ;
        RECT 632.250 460.500 633.450 461.400 ;
        RECT 626.250 459.300 633.450 460.500 ;
        RECT 502.950 452.850 505.050 454.950 ;
        RECT 536.100 453.150 537.900 454.950 ;
        RECT 503.100 451.050 504.900 452.850 ;
        RECT 535.950 451.050 538.050 453.150 ;
        RECT 539.550 451.950 540.750 459.300 ;
        RECT 581.250 458.250 585.000 459.300 ;
        RECT 583.950 454.950 585.150 458.250 ;
        RECT 587.100 456.150 588.900 457.950 ;
        RECT 542.100 453.150 543.900 454.950 ;
        RECT 498.750 449.400 501.000 450.300 ;
        RECT 538.950 449.850 541.050 451.950 ;
        RECT 541.950 451.050 544.050 453.150 ;
        RECT 583.950 452.850 586.050 454.950 ;
        RECT 586.950 454.050 589.050 456.150 ;
        RECT 626.250 454.950 627.450 459.300 ;
        RECT 668.400 456.150 669.600 464.400 ;
        RECT 707.850 460.200 709.650 467.250 ;
        RECT 712.350 461.400 714.150 467.250 ;
        RECT 748.650 461.400 750.450 467.250 ;
        RECT 707.850 459.300 711.450 460.200 ;
        RECT 589.950 452.850 592.050 454.950 ;
        RECT 625.950 452.850 628.050 454.950 ;
        RECT 631.950 452.850 634.050 454.950 ;
        RECT 667.950 454.050 670.050 456.150 ;
        RECT 670.950 455.850 673.050 457.950 ;
        RECT 671.100 454.050 672.900 455.850 ;
        RECT 580.950 449.850 583.050 451.950 ;
        RECT 498.750 448.500 504.450 449.400 ;
        RECT 413.550 435.750 415.350 441.600 ;
        RECT 416.550 435.750 418.350 441.600 ;
        RECT 419.550 435.750 421.350 441.600 ;
        RECT 455.550 435.750 457.350 441.600 ;
        RECT 458.850 435.750 460.650 447.600 ;
        RECT 461.850 435.750 463.650 447.600 ;
        RECT 496.350 435.750 498.150 447.600 ;
        RECT 499.350 435.750 501.150 447.600 ;
        RECT 503.250 441.600 504.450 448.500 ;
        RECT 539.550 441.600 540.750 449.850 ;
        RECT 581.250 448.050 583.050 449.850 ;
        RECT 584.850 447.600 586.050 452.850 ;
        RECT 590.100 451.050 591.900 452.850 ;
        RECT 626.250 449.400 627.450 452.850 ;
        RECT 632.100 451.050 633.900 452.850 ;
        RECT 626.250 448.500 633.450 449.400 ;
        RECT 626.250 447.600 627.450 448.500 ;
        RECT 502.650 435.750 504.450 441.600 ;
        RECT 536.550 435.750 538.350 441.600 ;
        RECT 539.550 435.750 541.350 441.600 ;
        RECT 542.550 435.750 544.350 441.600 ;
        RECT 581.400 435.750 583.200 441.600 ;
        RECT 584.700 435.750 586.500 447.600 ;
        RECT 588.900 435.750 590.700 447.600 ;
        RECT 622.650 435.750 624.450 447.600 ;
        RECT 625.650 435.750 627.450 447.600 ;
        RECT 628.650 435.750 630.450 447.600 ;
        RECT 631.650 435.750 633.450 448.500 ;
        RECT 634.650 435.750 636.450 447.600 ;
        RECT 668.400 441.600 669.600 454.050 ;
        RECT 707.100 453.150 708.900 454.950 ;
        RECT 706.950 451.050 709.050 453.150 ;
        RECT 710.250 451.950 711.450 459.300 ;
        RECT 749.250 459.300 750.450 461.400 ;
        RECT 751.650 462.300 753.450 467.250 ;
        RECT 754.650 463.200 756.450 467.250 ;
        RECT 757.650 462.300 759.450 467.250 ;
        RECT 751.650 460.950 759.450 462.300 ;
        RECT 749.250 458.250 753.000 459.300 ;
        RECT 751.950 454.950 753.150 458.250 ;
        RECT 755.100 456.150 756.900 457.950 ;
        RECT 713.100 453.150 714.900 454.950 ;
        RECT 709.950 449.850 712.050 451.950 ;
        RECT 712.950 451.050 715.050 453.150 ;
        RECT 751.950 452.850 754.050 454.950 ;
        RECT 754.950 454.050 757.050 456.150 ;
        RECT 757.950 452.850 760.050 454.950 ;
        RECT 748.950 449.850 751.050 451.950 ;
        RECT 710.250 441.600 711.450 449.850 ;
        RECT 749.250 448.050 751.050 449.850 ;
        RECT 752.850 447.600 754.050 452.850 ;
        RECT 758.100 451.050 759.900 452.850 ;
        RECT 667.650 435.750 669.450 441.600 ;
        RECT 670.650 435.750 672.450 441.600 ;
        RECT 706.650 435.750 708.450 441.600 ;
        RECT 709.650 435.750 711.450 441.600 ;
        RECT 712.650 435.750 714.450 441.600 ;
        RECT 749.400 435.750 751.200 441.600 ;
        RECT 752.700 435.750 754.500 447.600 ;
        RECT 756.900 435.750 758.700 447.600 ;
        RECT 3.150 419.400 4.950 431.250 ;
        RECT 6.150 425.400 7.950 431.250 ;
        RECT 11.250 425.400 13.050 431.250 ;
        RECT 16.050 425.400 17.850 431.250 ;
        RECT 11.550 424.500 12.750 425.400 ;
        RECT 19.050 424.500 20.850 431.250 ;
        RECT 22.950 425.400 24.750 431.250 ;
        RECT 27.150 425.400 28.950 431.250 ;
        RECT 31.650 428.400 33.450 431.250 ;
        RECT 7.950 422.400 12.750 424.500 ;
        RECT 15.150 422.700 22.050 424.500 ;
        RECT 27.150 423.300 31.050 425.400 ;
        RECT 11.550 421.500 12.750 422.400 ;
        RECT 24.450 421.800 26.250 422.400 ;
        RECT 11.550 420.300 19.050 421.500 ;
        RECT 17.250 419.700 19.050 420.300 ;
        RECT 19.950 420.900 26.250 421.800 ;
        RECT 3.150 418.800 14.250 419.400 ;
        RECT 19.950 418.800 20.850 420.900 ;
        RECT 24.450 420.600 26.250 420.900 ;
        RECT 27.150 420.600 29.850 422.400 ;
        RECT 27.150 419.700 28.050 420.600 ;
        RECT 3.150 418.200 20.850 418.800 ;
        RECT 3.150 405.600 4.050 418.200 ;
        RECT 12.450 417.900 20.850 418.200 ;
        RECT 22.050 418.800 28.050 419.700 ;
        RECT 28.950 418.800 31.050 419.700 ;
        RECT 34.650 419.400 36.450 431.250 ;
        RECT 12.450 417.600 14.250 417.900 ;
        RECT 22.050 414.150 22.950 418.800 ;
        RECT 28.950 417.600 33.150 418.800 ;
        RECT 32.250 415.800 34.050 417.600 ;
        RECT 13.950 413.100 16.050 414.150 ;
        RECT 5.100 411.150 6.900 412.950 ;
        RECT 8.100 412.050 16.050 413.100 ;
        RECT 19.950 412.050 22.950 414.150 ;
        RECT 8.100 411.300 9.900 412.050 ;
        RECT 6.000 410.400 6.900 411.150 ;
        RECT 11.100 410.400 12.900 411.000 ;
        RECT 6.000 409.200 12.900 410.400 ;
        RECT 11.850 408.000 12.900 409.200 ;
        RECT 22.050 408.000 22.950 412.050 ;
        RECT 31.950 411.750 34.050 412.050 ;
        RECT 30.150 409.950 34.050 411.750 ;
        RECT 35.250 409.950 36.450 419.400 ;
        RECT 11.850 407.100 22.950 408.000 ;
        RECT 31.950 407.850 36.450 409.950 ;
        RECT 11.850 406.200 12.900 407.100 ;
        RECT 22.050 406.800 22.950 407.100 ;
        RECT 3.150 399.750 4.950 405.600 ;
        RECT 7.950 403.500 10.050 405.600 ;
        RECT 11.550 404.400 13.350 406.200 ;
        RECT 14.850 405.450 16.650 406.200 ;
        RECT 14.850 404.400 19.800 405.450 ;
        RECT 22.050 405.000 23.850 406.800 ;
        RECT 35.250 405.600 36.450 407.850 ;
        RECT 28.950 404.700 31.050 405.600 ;
        RECT 9.000 402.600 10.050 403.500 ;
        RECT 18.750 402.600 19.800 404.400 ;
        RECT 27.300 403.500 31.050 404.700 ;
        RECT 27.300 402.600 28.350 403.500 ;
        RECT 6.150 399.750 7.950 402.600 ;
        RECT 9.000 401.700 12.750 402.600 ;
        RECT 10.950 399.750 12.750 401.700 ;
        RECT 15.450 399.750 17.250 402.600 ;
        RECT 18.750 399.750 20.550 402.600 ;
        RECT 22.650 399.750 24.450 402.600 ;
        RECT 26.850 399.750 28.650 402.600 ;
        RECT 31.350 399.750 33.150 402.600 ;
        RECT 34.650 399.750 36.450 405.600 ;
        RECT 39.150 419.400 40.950 431.250 ;
        RECT 42.150 425.400 43.950 431.250 ;
        RECT 47.250 425.400 49.050 431.250 ;
        RECT 52.050 425.400 53.850 431.250 ;
        RECT 47.550 424.500 48.750 425.400 ;
        RECT 55.050 424.500 56.850 431.250 ;
        RECT 58.950 425.400 60.750 431.250 ;
        RECT 63.150 425.400 64.950 431.250 ;
        RECT 67.650 428.400 69.450 431.250 ;
        RECT 43.950 422.400 48.750 424.500 ;
        RECT 51.150 422.700 58.050 424.500 ;
        RECT 63.150 423.300 67.050 425.400 ;
        RECT 47.550 421.500 48.750 422.400 ;
        RECT 60.450 421.800 62.250 422.400 ;
        RECT 47.550 420.300 55.050 421.500 ;
        RECT 53.250 419.700 55.050 420.300 ;
        RECT 55.950 420.900 62.250 421.800 ;
        RECT 39.150 418.800 50.250 419.400 ;
        RECT 55.950 418.800 56.850 420.900 ;
        RECT 60.450 420.600 62.250 420.900 ;
        RECT 63.150 420.600 65.850 422.400 ;
        RECT 63.150 419.700 64.050 420.600 ;
        RECT 39.150 418.200 56.850 418.800 ;
        RECT 39.150 405.600 40.050 418.200 ;
        RECT 48.450 417.900 56.850 418.200 ;
        RECT 58.050 418.800 64.050 419.700 ;
        RECT 64.950 418.800 67.050 419.700 ;
        RECT 70.650 419.400 72.450 431.250 ;
        RECT 48.450 417.600 50.250 417.900 ;
        RECT 58.050 414.150 58.950 418.800 ;
        RECT 64.950 417.600 69.150 418.800 ;
        RECT 68.250 415.800 70.050 417.600 ;
        RECT 49.950 413.100 52.050 414.150 ;
        RECT 41.100 411.150 42.900 412.950 ;
        RECT 44.100 412.050 52.050 413.100 ;
        RECT 55.950 412.050 58.950 414.150 ;
        RECT 44.100 411.300 45.900 412.050 ;
        RECT 42.000 410.400 42.900 411.150 ;
        RECT 47.100 410.400 48.900 411.000 ;
        RECT 42.000 409.200 48.900 410.400 ;
        RECT 47.850 408.000 48.900 409.200 ;
        RECT 58.050 408.000 58.950 412.050 ;
        RECT 67.950 411.750 70.050 412.050 ;
        RECT 66.150 409.950 70.050 411.750 ;
        RECT 71.250 409.950 72.450 419.400 ;
        RECT 47.850 407.100 58.950 408.000 ;
        RECT 67.950 407.850 72.450 409.950 ;
        RECT 47.850 406.200 48.900 407.100 ;
        RECT 58.050 406.800 58.950 407.100 ;
        RECT 39.150 399.750 40.950 405.600 ;
        RECT 43.950 403.500 46.050 405.600 ;
        RECT 47.550 404.400 49.350 406.200 ;
        RECT 50.850 405.450 52.650 406.200 ;
        RECT 50.850 404.400 55.800 405.450 ;
        RECT 58.050 405.000 59.850 406.800 ;
        RECT 71.250 405.600 72.450 407.850 ;
        RECT 64.950 404.700 67.050 405.600 ;
        RECT 45.000 402.600 46.050 403.500 ;
        RECT 54.750 402.600 55.800 404.400 ;
        RECT 63.300 403.500 67.050 404.700 ;
        RECT 63.300 402.600 64.350 403.500 ;
        RECT 42.150 399.750 43.950 402.600 ;
        RECT 45.000 401.700 48.750 402.600 ;
        RECT 46.950 399.750 48.750 401.700 ;
        RECT 51.450 399.750 53.250 402.600 ;
        RECT 54.750 399.750 56.550 402.600 ;
        RECT 58.650 399.750 60.450 402.600 ;
        RECT 62.850 399.750 64.650 402.600 ;
        RECT 67.350 399.750 69.150 402.600 ;
        RECT 70.650 399.750 72.450 405.600 ;
        RECT 75.150 419.400 76.950 431.250 ;
        RECT 78.150 425.400 79.950 431.250 ;
        RECT 83.250 425.400 85.050 431.250 ;
        RECT 88.050 425.400 89.850 431.250 ;
        RECT 83.550 424.500 84.750 425.400 ;
        RECT 91.050 424.500 92.850 431.250 ;
        RECT 94.950 425.400 96.750 431.250 ;
        RECT 99.150 425.400 100.950 431.250 ;
        RECT 103.650 428.400 105.450 431.250 ;
        RECT 79.950 422.400 84.750 424.500 ;
        RECT 87.150 422.700 94.050 424.500 ;
        RECT 99.150 423.300 103.050 425.400 ;
        RECT 83.550 421.500 84.750 422.400 ;
        RECT 96.450 421.800 98.250 422.400 ;
        RECT 83.550 420.300 91.050 421.500 ;
        RECT 89.250 419.700 91.050 420.300 ;
        RECT 91.950 420.900 98.250 421.800 ;
        RECT 75.150 418.800 86.250 419.400 ;
        RECT 91.950 418.800 92.850 420.900 ;
        RECT 96.450 420.600 98.250 420.900 ;
        RECT 99.150 420.600 101.850 422.400 ;
        RECT 99.150 419.700 100.050 420.600 ;
        RECT 75.150 418.200 92.850 418.800 ;
        RECT 75.150 405.600 76.050 418.200 ;
        RECT 84.450 417.900 92.850 418.200 ;
        RECT 94.050 418.800 100.050 419.700 ;
        RECT 100.950 418.800 103.050 419.700 ;
        RECT 106.650 419.400 108.450 431.250 ;
        RECT 143.400 425.400 145.200 431.250 ;
        RECT 146.700 419.400 148.500 431.250 ;
        RECT 150.900 419.400 152.700 431.250 ;
        RECT 187.650 430.500 195.450 431.250 ;
        RECT 187.650 419.400 189.450 430.500 ;
        RECT 190.650 419.400 192.450 429.600 ;
        RECT 193.650 420.600 195.450 430.500 ;
        RECT 196.650 421.500 198.450 431.250 ;
        RECT 199.650 420.600 201.450 431.250 ;
        RECT 193.650 419.700 201.450 420.600 ;
        RECT 230.550 419.400 232.350 431.250 ;
        RECT 234.750 419.400 236.550 431.250 ;
        RECT 276.150 420.900 277.950 431.250 ;
        RECT 84.450 417.600 86.250 417.900 ;
        RECT 94.050 414.150 94.950 418.800 ;
        RECT 100.950 417.600 105.150 418.800 ;
        RECT 104.250 415.800 106.050 417.600 ;
        RECT 85.950 413.100 88.050 414.150 ;
        RECT 77.100 411.150 78.900 412.950 ;
        RECT 80.100 412.050 88.050 413.100 ;
        RECT 91.950 412.050 94.950 414.150 ;
        RECT 80.100 411.300 81.900 412.050 ;
        RECT 78.000 410.400 78.900 411.150 ;
        RECT 83.100 410.400 84.900 411.000 ;
        RECT 78.000 409.200 84.900 410.400 ;
        RECT 83.850 408.000 84.900 409.200 ;
        RECT 94.050 408.000 94.950 412.050 ;
        RECT 103.950 411.750 106.050 412.050 ;
        RECT 102.150 409.950 106.050 411.750 ;
        RECT 107.250 409.950 108.450 419.400 ;
        RECT 143.250 417.150 145.050 418.950 ;
        RECT 142.950 415.050 145.050 417.150 ;
        RECT 146.850 414.150 148.050 419.400 ;
        RECT 190.800 418.500 192.600 419.400 ;
        RECT 190.800 417.600 194.850 418.500 ;
        RECT 152.100 414.150 153.900 415.950 ;
        RECT 188.100 414.150 189.900 415.950 ;
        RECT 193.950 414.150 194.850 417.600 ;
        RECT 234.000 418.350 236.550 419.400 ;
        RECT 275.550 419.550 277.950 420.900 ;
        RECT 279.150 419.550 280.950 431.250 ;
        RECT 199.950 414.150 201.750 415.950 ;
        RECT 230.100 414.150 231.900 415.950 ;
        RECT 83.850 407.100 94.950 408.000 ;
        RECT 103.950 407.850 108.450 409.950 ;
        RECT 145.950 412.050 148.050 414.150 ;
        RECT 145.950 408.750 147.150 412.050 ;
        RECT 148.950 410.850 151.050 412.950 ;
        RECT 151.950 412.050 154.050 414.150 ;
        RECT 187.950 412.050 190.050 414.150 ;
        RECT 190.950 410.850 193.050 412.950 ;
        RECT 193.950 412.050 196.050 414.150 ;
        RECT 149.100 409.050 150.900 410.850 ;
        RECT 191.250 409.050 193.050 410.850 ;
        RECT 83.850 406.200 84.900 407.100 ;
        RECT 94.050 406.800 94.950 407.100 ;
        RECT 75.150 399.750 76.950 405.600 ;
        RECT 79.950 403.500 82.050 405.600 ;
        RECT 83.550 404.400 85.350 406.200 ;
        RECT 86.850 405.450 88.650 406.200 ;
        RECT 86.850 404.400 91.800 405.450 ;
        RECT 94.050 405.000 95.850 406.800 ;
        RECT 107.250 405.600 108.450 407.850 ;
        RECT 143.250 407.700 147.000 408.750 ;
        RECT 160.950 408.450 163.050 409.050 ;
        RECT 187.950 408.450 190.050 409.050 ;
        RECT 143.250 405.600 144.450 407.700 ;
        RECT 160.950 407.550 190.050 408.450 ;
        RECT 160.950 406.950 163.050 407.550 ;
        RECT 187.950 406.950 190.050 407.550 ;
        RECT 100.950 404.700 103.050 405.600 ;
        RECT 81.000 402.600 82.050 403.500 ;
        RECT 90.750 402.600 91.800 404.400 ;
        RECT 99.300 403.500 103.050 404.700 ;
        RECT 99.300 402.600 100.350 403.500 ;
        RECT 78.150 399.750 79.950 402.600 ;
        RECT 81.000 401.700 84.750 402.600 ;
        RECT 82.950 399.750 84.750 401.700 ;
        RECT 87.450 399.750 89.250 402.600 ;
        RECT 90.750 399.750 92.550 402.600 ;
        RECT 94.650 399.750 96.450 402.600 ;
        RECT 98.850 399.750 100.650 402.600 ;
        RECT 103.350 399.750 105.150 402.600 ;
        RECT 106.650 399.750 108.450 405.600 ;
        RECT 142.650 399.750 144.450 405.600 ;
        RECT 145.650 404.700 153.450 406.050 ;
        RECT 195.000 405.600 196.050 412.050 ;
        RECT 196.950 410.850 199.050 412.950 ;
        RECT 199.950 412.050 202.050 414.150 ;
        RECT 229.950 412.050 232.050 414.150 ;
        RECT 234.000 411.150 235.050 418.350 ;
        RECT 236.100 414.150 237.900 415.950 ;
        RECT 235.950 412.050 238.050 414.150 ;
        RECT 275.550 412.950 276.900 419.550 ;
        RECT 283.650 419.400 285.450 431.250 ;
        RECT 314.550 425.400 316.350 431.250 ;
        RECT 317.550 425.400 319.350 431.250 ;
        RECT 320.550 426.000 322.350 431.250 ;
        RECT 317.700 425.100 319.350 425.400 ;
        RECT 323.550 425.400 325.350 431.250 ;
        RECT 356.550 425.400 358.350 431.250 ;
        RECT 359.550 425.400 361.350 431.250 ;
        RECT 362.550 425.400 364.350 431.250 ;
        RECT 398.550 425.400 400.350 431.250 ;
        RECT 401.550 425.400 403.350 431.250 ;
        RECT 404.550 426.000 406.350 431.250 ;
        RECT 323.550 425.100 324.750 425.400 ;
        RECT 317.700 424.200 324.750 425.100 ;
        RECT 317.100 420.150 318.900 421.950 ;
        RECT 278.250 418.200 280.050 418.650 ;
        RECT 284.250 418.200 285.450 419.400 ;
        RECT 278.250 417.000 285.450 418.200 ;
        RECT 314.100 417.150 315.900 418.950 ;
        RECT 316.950 418.050 319.050 420.150 ;
        RECT 320.250 417.150 322.050 418.950 ;
        RECT 278.250 416.850 280.050 417.000 ;
        RECT 196.950 409.050 198.750 410.850 ;
        RECT 232.950 409.050 235.050 411.150 ;
        RECT 145.650 399.750 147.450 404.700 ;
        RECT 148.650 399.750 150.450 403.800 ;
        RECT 151.650 399.750 153.450 404.700 ;
        RECT 190.800 399.750 192.600 405.600 ;
        RECT 195.000 399.750 196.800 405.600 ;
        RECT 199.200 399.750 201.000 405.600 ;
        RECT 234.000 402.600 235.050 409.050 ;
        RECT 274.950 410.850 277.050 412.950 ;
        RECT 274.950 405.600 276.000 410.850 ;
        RECT 278.400 408.600 279.300 416.850 ;
        RECT 281.100 414.150 282.900 415.950 ;
        RECT 313.950 415.050 316.050 417.150 ;
        RECT 319.950 415.050 322.050 417.150 ;
        RECT 323.700 415.950 324.750 424.200 ;
        RECT 359.550 417.150 360.750 425.400 ;
        RECT 401.700 425.100 403.350 425.400 ;
        RECT 407.550 425.400 409.350 431.250 ;
        RECT 443.550 425.400 445.350 431.250 ;
        RECT 407.550 425.100 408.750 425.400 ;
        RECT 401.700 424.200 408.750 425.100 ;
        RECT 401.100 420.150 402.900 421.950 ;
        RECT 398.100 417.150 399.900 418.950 ;
        RECT 400.950 418.050 403.050 420.150 ;
        RECT 404.250 417.150 406.050 418.950 ;
        RECT 280.950 412.050 283.050 414.150 ;
        RECT 322.950 413.850 325.050 415.950 ;
        RECT 355.950 413.850 358.050 415.950 ;
        RECT 358.950 415.050 361.050 417.150 ;
        RECT 284.100 411.150 285.900 412.950 ;
        RECT 283.950 409.050 286.050 411.150 ;
        RECT 323.400 409.650 324.600 413.850 ;
        RECT 356.100 412.050 357.900 413.850 ;
        RECT 278.250 407.700 280.050 408.600 ;
        RECT 278.250 406.800 281.550 407.700 ;
        RECT 230.550 399.750 232.350 402.600 ;
        RECT 233.550 399.750 235.350 402.600 ;
        RECT 236.550 399.750 238.350 402.600 ;
        RECT 274.650 399.750 276.450 405.600 ;
        RECT 280.650 402.600 281.550 406.800 ;
        RECT 277.650 399.750 279.450 402.600 ;
        RECT 280.650 399.750 282.450 402.600 ;
        RECT 283.650 399.750 285.450 402.600 ;
        RECT 314.700 399.750 316.500 408.600 ;
        RECT 320.100 408.000 324.600 409.650 ;
        RECT 320.100 399.750 321.900 408.000 ;
        RECT 359.550 407.700 360.750 415.050 ;
        RECT 361.950 413.850 364.050 415.950 ;
        RECT 397.950 415.050 400.050 417.150 ;
        RECT 403.950 415.050 406.050 417.150 ;
        RECT 407.700 415.950 408.750 424.200 ;
        RECT 443.550 418.500 444.750 425.400 ;
        RECT 446.850 419.400 448.650 431.250 ;
        RECT 449.850 419.400 451.650 431.250 ;
        RECT 488.400 425.400 490.200 431.250 ;
        RECT 491.700 419.400 493.500 431.250 ;
        RECT 495.900 419.400 497.700 431.250 ;
        RECT 501.150 419.400 502.950 431.250 ;
        RECT 504.150 425.400 505.950 431.250 ;
        RECT 509.250 425.400 511.050 431.250 ;
        RECT 514.050 425.400 515.850 431.250 ;
        RECT 509.550 424.500 510.750 425.400 ;
        RECT 517.050 424.500 518.850 431.250 ;
        RECT 520.950 425.400 522.750 431.250 ;
        RECT 525.150 425.400 526.950 431.250 ;
        RECT 529.650 428.400 531.450 431.250 ;
        RECT 505.950 422.400 510.750 424.500 ;
        RECT 513.150 422.700 520.050 424.500 ;
        RECT 525.150 423.300 529.050 425.400 ;
        RECT 509.550 421.500 510.750 422.400 ;
        RECT 522.450 421.800 524.250 422.400 ;
        RECT 509.550 420.300 517.050 421.500 ;
        RECT 515.250 419.700 517.050 420.300 ;
        RECT 517.950 420.900 524.250 421.800 ;
        RECT 443.550 417.600 449.250 418.500 ;
        RECT 447.000 416.700 449.250 417.600 ;
        RECT 406.950 413.850 409.050 415.950 ;
        RECT 443.100 414.150 444.900 415.950 ;
        RECT 362.100 412.050 363.900 413.850 ;
        RECT 407.400 409.650 408.600 413.850 ;
        RECT 442.950 412.050 445.050 414.150 ;
        RECT 359.550 406.800 363.150 407.700 ;
        RECT 356.850 399.750 358.650 405.600 ;
        RECT 361.350 399.750 363.150 406.800 ;
        RECT 398.700 399.750 400.500 408.600 ;
        RECT 404.100 408.000 408.600 409.650 ;
        RECT 447.000 408.300 448.050 416.700 ;
        RECT 450.150 414.150 451.350 419.400 ;
        RECT 488.250 417.150 490.050 418.950 ;
        RECT 487.950 415.050 490.050 417.150 ;
        RECT 491.850 414.150 493.050 419.400 ;
        RECT 501.150 418.800 512.250 419.400 ;
        RECT 517.950 418.800 518.850 420.900 ;
        RECT 522.450 420.600 524.250 420.900 ;
        RECT 525.150 420.600 527.850 422.400 ;
        RECT 525.150 419.700 526.050 420.600 ;
        RECT 501.150 418.200 518.850 418.800 ;
        RECT 497.100 414.150 498.900 415.950 ;
        RECT 448.950 412.050 451.350 414.150 ;
        RECT 404.100 399.750 405.900 408.000 ;
        RECT 447.000 407.400 449.250 408.300 ;
        RECT 444.150 406.500 449.250 407.400 ;
        RECT 444.150 402.600 445.350 406.500 ;
        RECT 450.150 405.600 451.350 412.050 ;
        RECT 490.950 412.050 493.050 414.150 ;
        RECT 490.950 408.750 492.150 412.050 ;
        RECT 493.950 410.850 496.050 412.950 ;
        RECT 496.950 412.050 499.050 414.150 ;
        RECT 494.100 409.050 495.900 410.850 ;
        RECT 488.250 407.700 492.000 408.750 ;
        RECT 488.250 405.600 489.450 407.700 ;
        RECT 443.550 399.750 445.350 402.600 ;
        RECT 446.850 399.750 448.650 405.600 ;
        RECT 449.850 399.750 451.650 405.600 ;
        RECT 487.650 399.750 489.450 405.600 ;
        RECT 490.650 404.700 498.450 406.050 ;
        RECT 490.650 399.750 492.450 404.700 ;
        RECT 493.650 399.750 495.450 403.800 ;
        RECT 496.650 399.750 498.450 404.700 ;
        RECT 501.150 405.600 502.050 418.200 ;
        RECT 510.450 417.900 518.850 418.200 ;
        RECT 520.050 418.800 526.050 419.700 ;
        RECT 526.950 418.800 529.050 419.700 ;
        RECT 532.650 419.400 534.450 431.250 ;
        RECT 569.400 425.400 571.200 431.250 ;
        RECT 572.700 419.400 574.500 431.250 ;
        RECT 576.900 419.400 578.700 431.250 ;
        RECT 611.550 425.400 613.350 431.250 ;
        RECT 614.550 425.400 616.350 431.250 ;
        RECT 653.400 425.400 655.200 431.250 ;
        RECT 510.450 417.600 512.250 417.900 ;
        RECT 520.050 414.150 520.950 418.800 ;
        RECT 526.950 417.600 531.150 418.800 ;
        RECT 530.250 415.800 532.050 417.600 ;
        RECT 511.950 413.100 514.050 414.150 ;
        RECT 503.100 411.150 504.900 412.950 ;
        RECT 506.100 412.050 514.050 413.100 ;
        RECT 517.950 412.050 520.950 414.150 ;
        RECT 506.100 411.300 507.900 412.050 ;
        RECT 504.000 410.400 504.900 411.150 ;
        RECT 509.100 410.400 510.900 411.000 ;
        RECT 504.000 409.200 510.900 410.400 ;
        RECT 509.850 408.000 510.900 409.200 ;
        RECT 520.050 408.000 520.950 412.050 ;
        RECT 529.950 411.750 532.050 412.050 ;
        RECT 528.150 409.950 532.050 411.750 ;
        RECT 533.250 409.950 534.450 419.400 ;
        RECT 569.250 417.150 571.050 418.950 ;
        RECT 568.950 415.050 571.050 417.150 ;
        RECT 572.850 414.150 574.050 419.400 ;
        RECT 578.100 414.150 579.900 415.950 ;
        RECT 509.850 407.100 520.950 408.000 ;
        RECT 529.950 407.850 534.450 409.950 ;
        RECT 571.950 412.050 574.050 414.150 ;
        RECT 571.950 408.750 573.150 412.050 ;
        RECT 574.950 410.850 577.050 412.950 ;
        RECT 577.950 412.050 580.050 414.150 ;
        RECT 614.400 412.950 615.600 425.400 ;
        RECT 656.700 419.400 658.500 431.250 ;
        RECT 660.900 419.400 662.700 431.250 ;
        RECT 692.550 425.400 694.350 431.250 ;
        RECT 653.250 417.150 655.050 418.950 ;
        RECT 652.950 415.050 655.050 417.150 ;
        RECT 656.850 414.150 658.050 419.400 ;
        RECT 692.550 418.500 693.750 425.400 ;
        RECT 695.850 419.400 697.650 431.250 ;
        RECT 698.850 419.400 700.650 431.250 ;
        RECT 733.350 419.400 735.150 431.250 ;
        RECT 736.350 419.400 738.150 431.250 ;
        RECT 739.650 425.400 741.450 431.250 ;
        RECT 692.550 417.600 698.250 418.500 ;
        RECT 696.000 416.700 698.250 417.600 ;
        RECT 662.100 414.150 663.900 415.950 ;
        RECT 692.100 414.150 693.900 415.950 ;
        RECT 611.100 411.150 612.900 412.950 ;
        RECT 575.100 409.050 576.900 410.850 ;
        RECT 610.950 409.050 613.050 411.150 ;
        RECT 613.950 410.850 616.050 412.950 ;
        RECT 655.950 412.050 658.050 414.150 ;
        RECT 509.850 406.200 510.900 407.100 ;
        RECT 520.050 406.800 520.950 407.100 ;
        RECT 501.150 399.750 502.950 405.600 ;
        RECT 505.950 403.500 508.050 405.600 ;
        RECT 509.550 404.400 511.350 406.200 ;
        RECT 512.850 405.450 514.650 406.200 ;
        RECT 512.850 404.400 517.800 405.450 ;
        RECT 520.050 405.000 521.850 406.800 ;
        RECT 533.250 405.600 534.450 407.850 ;
        RECT 569.250 407.700 573.000 408.750 ;
        RECT 569.250 405.600 570.450 407.700 ;
        RECT 526.950 404.700 529.050 405.600 ;
        RECT 507.000 402.600 508.050 403.500 ;
        RECT 516.750 402.600 517.800 404.400 ;
        RECT 525.300 403.500 529.050 404.700 ;
        RECT 525.300 402.600 526.350 403.500 ;
        RECT 504.150 399.750 505.950 402.600 ;
        RECT 507.000 401.700 510.750 402.600 ;
        RECT 508.950 399.750 510.750 401.700 ;
        RECT 513.450 399.750 515.250 402.600 ;
        RECT 516.750 399.750 518.550 402.600 ;
        RECT 520.650 399.750 522.450 402.600 ;
        RECT 524.850 399.750 526.650 402.600 ;
        RECT 529.350 399.750 531.150 402.600 ;
        RECT 532.650 399.750 534.450 405.600 ;
        RECT 568.650 399.750 570.450 405.600 ;
        RECT 571.650 404.700 579.450 406.050 ;
        RECT 571.650 399.750 573.450 404.700 ;
        RECT 574.650 399.750 576.450 403.800 ;
        RECT 577.650 399.750 579.450 404.700 ;
        RECT 614.400 402.600 615.600 410.850 ;
        RECT 655.950 408.750 657.150 412.050 ;
        RECT 658.950 410.850 661.050 412.950 ;
        RECT 661.950 412.050 664.050 414.150 ;
        RECT 691.950 412.050 694.050 414.150 ;
        RECT 659.100 409.050 660.900 410.850 ;
        RECT 653.250 407.700 657.000 408.750 ;
        RECT 696.000 408.300 697.050 416.700 ;
        RECT 699.150 414.150 700.350 419.400 ;
        RECT 697.950 412.050 700.350 414.150 ;
        RECT 653.250 405.600 654.450 407.700 ;
        RECT 696.000 407.400 698.250 408.300 ;
        RECT 693.150 406.500 698.250 407.400 ;
        RECT 611.550 399.750 613.350 402.600 ;
        RECT 614.550 399.750 616.350 402.600 ;
        RECT 652.650 399.750 654.450 405.600 ;
        RECT 655.650 404.700 663.450 406.050 ;
        RECT 655.650 399.750 657.450 404.700 ;
        RECT 658.650 399.750 660.450 403.800 ;
        RECT 661.650 399.750 663.450 404.700 ;
        RECT 693.150 402.600 694.350 406.500 ;
        RECT 699.150 405.600 700.350 412.050 ;
        RECT 733.650 414.150 734.850 419.400 ;
        RECT 740.250 418.500 741.450 425.400 ;
        RECT 735.750 417.600 741.450 418.500 ;
        RECT 735.750 416.700 738.000 417.600 ;
        RECT 733.650 412.050 736.050 414.150 ;
        RECT 733.650 405.600 734.850 412.050 ;
        RECT 736.950 408.300 738.000 416.700 ;
        RECT 740.100 414.150 741.900 415.950 ;
        RECT 739.950 412.050 742.050 414.150 ;
        RECT 735.750 407.400 738.000 408.300 ;
        RECT 735.750 406.500 740.850 407.400 ;
        RECT 692.550 399.750 694.350 402.600 ;
        RECT 695.850 399.750 697.650 405.600 ;
        RECT 698.850 399.750 700.650 405.600 ;
        RECT 733.350 399.750 735.150 405.600 ;
        RECT 736.350 399.750 738.150 405.600 ;
        RECT 739.650 402.600 740.850 406.500 ;
        RECT 739.650 399.750 741.450 402.600 ;
        RECT 34.650 389.400 36.450 395.250 ;
        RECT 35.250 387.300 36.450 389.400 ;
        RECT 37.650 390.300 39.450 395.250 ;
        RECT 40.650 391.200 42.450 395.250 ;
        RECT 43.650 390.300 45.450 395.250 ;
        RECT 37.650 388.950 45.450 390.300 ;
        RECT 74.550 390.300 76.350 395.250 ;
        RECT 77.550 391.200 79.350 395.250 ;
        RECT 80.550 390.300 82.350 395.250 ;
        RECT 74.550 388.950 82.350 390.300 ;
        RECT 83.550 389.400 85.350 395.250 ;
        RECT 121.650 392.400 123.450 395.250 ;
        RECT 124.650 392.400 126.450 395.250 ;
        RECT 83.550 387.300 84.750 389.400 ;
        RECT 35.250 386.250 39.000 387.300 ;
        RECT 81.000 386.250 84.750 387.300 ;
        RECT 37.950 382.950 39.150 386.250 ;
        RECT 41.100 384.150 42.900 385.950 ;
        RECT 77.100 384.150 78.900 385.950 ;
        RECT 37.950 380.850 40.050 382.950 ;
        RECT 40.950 382.050 43.050 384.150 ;
        RECT 43.950 380.850 46.050 382.950 ;
        RECT 73.950 380.850 76.050 382.950 ;
        RECT 76.950 382.050 79.050 384.150 ;
        RECT 80.850 382.950 82.050 386.250 ;
        RECT 122.400 384.150 123.600 392.400 ;
        RECT 157.650 389.400 159.450 395.250 ;
        RECT 160.650 392.400 162.450 395.250 ;
        RECT 163.650 392.400 165.450 395.250 ;
        RECT 166.650 392.400 168.450 395.250 ;
        RECT 79.950 380.850 82.050 382.950 ;
        RECT 121.950 382.050 124.050 384.150 ;
        RECT 124.950 383.850 127.050 385.950 ;
        RECT 157.950 384.150 159.000 389.400 ;
        RECT 163.650 388.200 164.550 392.400 ;
        RECT 201.000 389.400 202.800 395.250 ;
        RECT 205.200 391.050 207.000 395.250 ;
        RECT 208.500 392.400 210.300 395.250 ;
        RECT 245.550 392.400 247.350 395.250 ;
        RECT 248.550 392.400 250.350 395.250 ;
        RECT 205.200 389.400 210.900 391.050 ;
        RECT 161.250 387.300 164.550 388.200 ;
        RECT 161.250 386.400 163.050 387.300 ;
        RECT 125.100 382.050 126.900 383.850 ;
        RECT 157.950 382.050 160.050 384.150 ;
        RECT 34.950 377.850 37.050 379.950 ;
        RECT 35.250 376.050 37.050 377.850 ;
        RECT 38.850 375.600 40.050 380.850 ;
        RECT 44.100 379.050 45.900 380.850 ;
        RECT 74.100 379.050 75.900 380.850 ;
        RECT 79.950 375.600 81.150 380.850 ;
        RECT 82.950 377.850 85.050 379.950 ;
        RECT 82.950 376.050 84.750 377.850 ;
        RECT 35.400 363.750 37.200 369.600 ;
        RECT 38.700 363.750 40.500 375.600 ;
        RECT 42.900 363.750 44.700 375.600 ;
        RECT 75.300 363.750 77.100 375.600 ;
        RECT 79.500 363.750 81.300 375.600 ;
        RECT 122.400 369.600 123.600 382.050 ;
        RECT 158.550 375.450 159.900 382.050 ;
        RECT 161.400 378.150 162.300 386.400 ;
        RECT 166.950 383.850 169.050 385.950 ;
        RECT 200.100 384.150 201.900 385.950 ;
        RECT 163.950 380.850 166.050 382.950 ;
        RECT 167.100 382.050 168.900 383.850 ;
        RECT 199.950 382.050 202.050 384.150 ;
        RECT 202.950 383.850 205.050 385.950 ;
        RECT 206.100 384.150 207.900 385.950 ;
        RECT 203.100 382.050 204.900 383.850 ;
        RECT 205.950 382.050 208.050 384.150 ;
        RECT 209.700 382.950 210.900 389.400 ;
        RECT 244.950 383.850 247.050 385.950 ;
        RECT 248.400 384.150 249.600 392.400 ;
        RECT 286.650 389.400 288.450 395.250 ;
        RECT 287.250 387.300 288.450 389.400 ;
        RECT 289.650 390.300 291.450 395.250 ;
        RECT 292.650 391.200 294.450 395.250 ;
        RECT 295.650 390.300 297.450 395.250 ;
        RECT 289.650 388.950 297.450 390.300 ;
        RECT 328.650 389.400 330.450 395.250 ;
        RECT 329.250 387.300 330.450 389.400 ;
        RECT 331.650 390.300 333.450 395.250 ;
        RECT 334.650 391.200 336.450 395.250 ;
        RECT 337.650 390.300 339.450 395.250 ;
        RECT 371.550 392.400 373.350 395.250 ;
        RECT 374.550 392.400 376.350 395.250 ;
        RECT 377.550 392.400 379.350 395.250 ;
        RECT 331.650 388.950 339.450 390.300 ;
        RECT 375.450 388.200 376.350 392.400 ;
        RECT 380.550 389.400 382.350 395.250 ;
        RECT 387.150 389.400 388.950 395.250 ;
        RECT 390.150 392.400 391.950 395.250 ;
        RECT 394.950 393.300 396.750 395.250 ;
        RECT 393.000 392.400 396.750 393.300 ;
        RECT 399.450 392.400 401.250 395.250 ;
        RECT 402.750 392.400 404.550 395.250 ;
        RECT 406.650 392.400 408.450 395.250 ;
        RECT 410.850 392.400 412.650 395.250 ;
        RECT 415.350 392.400 417.150 395.250 ;
        RECT 393.000 391.500 394.050 392.400 ;
        RECT 391.950 389.400 394.050 391.500 ;
        RECT 402.750 390.600 403.800 392.400 ;
        RECT 375.450 387.300 378.750 388.200 ;
        RECT 287.250 386.250 291.000 387.300 ;
        RECT 329.250 386.250 333.000 387.300 ;
        RECT 376.950 386.400 378.750 387.300 ;
        RECT 208.950 380.850 211.050 382.950 ;
        RECT 245.100 382.050 246.900 383.850 ;
        RECT 247.950 382.050 250.050 384.150 ;
        RECT 289.950 382.950 291.150 386.250 ;
        RECT 293.100 384.150 294.900 385.950 ;
        RECT 164.100 379.050 165.900 380.850 ;
        RECT 161.250 378.000 163.050 378.150 ;
        RECT 161.250 376.800 168.450 378.000 ;
        RECT 161.250 376.350 163.050 376.800 ;
        RECT 167.250 375.600 168.450 376.800 ;
        RECT 209.700 375.600 210.900 380.850 ;
        RECT 158.550 374.100 160.950 375.450 ;
        RECT 82.800 363.750 84.600 369.600 ;
        RECT 121.650 363.750 123.450 369.600 ;
        RECT 124.650 363.750 126.450 369.600 ;
        RECT 159.150 363.750 160.950 374.100 ;
        RECT 162.150 363.750 163.950 375.450 ;
        RECT 166.650 363.750 168.450 375.600 ;
        RECT 200.550 374.700 208.350 375.600 ;
        RECT 200.550 363.750 202.350 374.700 ;
        RECT 203.550 363.750 205.350 373.800 ;
        RECT 206.550 363.750 208.350 374.700 ;
        RECT 209.550 363.750 211.350 375.600 ;
        RECT 248.400 369.600 249.600 382.050 ;
        RECT 289.950 380.850 292.050 382.950 ;
        RECT 292.950 382.050 295.050 384.150 ;
        RECT 331.950 382.950 333.150 386.250 ;
        RECT 335.100 384.150 336.900 385.950 ;
        RECT 295.950 380.850 298.050 382.950 ;
        RECT 331.950 380.850 334.050 382.950 ;
        RECT 334.950 382.050 337.050 384.150 ;
        RECT 370.950 383.850 373.050 385.950 ;
        RECT 337.950 380.850 340.050 382.950 ;
        RECT 371.100 382.050 372.900 383.850 ;
        RECT 373.950 380.850 376.050 382.950 ;
        RECT 286.950 377.850 289.050 379.950 ;
        RECT 287.250 376.050 289.050 377.850 ;
        RECT 290.850 375.600 292.050 380.850 ;
        RECT 296.100 379.050 297.900 380.850 ;
        RECT 328.950 377.850 331.050 379.950 ;
        RECT 329.250 376.050 331.050 377.850 ;
        RECT 332.850 375.600 334.050 380.850 ;
        RECT 338.100 379.050 339.900 380.850 ;
        RECT 374.100 379.050 375.900 380.850 ;
        RECT 377.700 378.150 378.600 386.400 ;
        RECT 381.000 384.150 382.050 389.400 ;
        RECT 379.950 382.050 382.050 384.150 ;
        RECT 376.950 378.000 378.750 378.150 ;
        RECT 371.550 376.800 378.750 378.000 ;
        RECT 371.550 375.600 372.750 376.800 ;
        RECT 376.950 376.350 378.750 376.800 ;
        RECT 245.550 363.750 247.350 369.600 ;
        RECT 248.550 363.750 250.350 369.600 ;
        RECT 287.400 363.750 289.200 369.600 ;
        RECT 290.700 363.750 292.500 375.600 ;
        RECT 294.900 363.750 296.700 375.600 ;
        RECT 329.400 363.750 331.200 369.600 ;
        RECT 332.700 363.750 334.500 375.600 ;
        RECT 336.900 363.750 338.700 375.600 ;
        RECT 371.550 363.750 373.350 375.600 ;
        RECT 380.100 375.450 381.450 382.050 ;
        RECT 376.050 363.750 377.850 375.450 ;
        RECT 379.050 374.100 381.450 375.450 ;
        RECT 387.150 376.800 388.050 389.400 ;
        RECT 395.550 388.800 397.350 390.600 ;
        RECT 398.850 389.550 403.800 390.600 ;
        RECT 411.300 391.500 412.350 392.400 ;
        RECT 411.300 390.300 415.050 391.500 ;
        RECT 398.850 388.800 400.650 389.550 ;
        RECT 395.850 387.900 396.900 388.800 ;
        RECT 406.050 388.200 407.850 390.000 ;
        RECT 412.950 389.400 415.050 390.300 ;
        RECT 418.650 389.400 420.450 395.250 ;
        RECT 454.650 389.400 456.450 395.250 ;
        RECT 406.050 387.900 406.950 388.200 ;
        RECT 395.850 387.000 406.950 387.900 ;
        RECT 419.250 387.150 420.450 389.400 ;
        RECT 395.850 385.800 396.900 387.000 ;
        RECT 390.000 384.600 396.900 385.800 ;
        RECT 390.000 383.850 390.900 384.600 ;
        RECT 395.100 384.000 396.900 384.600 ;
        RECT 389.100 382.050 390.900 383.850 ;
        RECT 392.100 382.950 393.900 383.700 ;
        RECT 406.050 382.950 406.950 387.000 ;
        RECT 415.950 385.050 420.450 387.150 ;
        RECT 455.250 387.300 456.450 389.400 ;
        RECT 457.650 390.300 459.450 395.250 ;
        RECT 460.650 391.200 462.450 395.250 ;
        RECT 463.650 390.300 465.450 395.250 ;
        RECT 499.650 392.400 501.450 395.250 ;
        RECT 502.650 392.400 504.450 395.250 ;
        RECT 457.650 388.950 465.450 390.300 ;
        RECT 455.250 386.250 459.000 387.300 ;
        RECT 414.150 383.250 418.050 385.050 ;
        RECT 415.950 382.950 418.050 383.250 ;
        RECT 392.100 381.900 400.050 382.950 ;
        RECT 397.950 380.850 400.050 381.900 ;
        RECT 403.950 380.850 406.950 382.950 ;
        RECT 396.450 377.100 398.250 377.400 ;
        RECT 396.450 376.800 404.850 377.100 ;
        RECT 387.150 376.200 404.850 376.800 ;
        RECT 387.150 375.600 398.250 376.200 ;
        RECT 379.050 363.750 380.850 374.100 ;
        RECT 387.150 363.750 388.950 375.600 ;
        RECT 401.250 374.700 403.050 375.300 ;
        RECT 395.550 373.500 403.050 374.700 ;
        RECT 403.950 374.100 404.850 376.200 ;
        RECT 406.050 376.200 406.950 380.850 ;
        RECT 416.250 377.400 418.050 379.200 ;
        RECT 412.950 376.200 417.150 377.400 ;
        RECT 406.050 375.300 412.050 376.200 ;
        RECT 412.950 375.300 415.050 376.200 ;
        RECT 419.250 375.600 420.450 385.050 ;
        RECT 457.950 382.950 459.150 386.250 ;
        RECT 461.100 384.150 462.900 385.950 ;
        RECT 500.400 384.150 501.600 392.400 ;
        RECT 538.350 389.400 540.150 395.250 ;
        RECT 541.350 389.400 543.150 395.250 ;
        RECT 544.650 392.400 546.450 395.250 ;
        RECT 457.950 380.850 460.050 382.950 ;
        RECT 460.950 382.050 463.050 384.150 ;
        RECT 463.950 380.850 466.050 382.950 ;
        RECT 499.950 382.050 502.050 384.150 ;
        RECT 502.950 383.850 505.050 385.950 ;
        RECT 503.100 382.050 504.900 383.850 ;
        RECT 538.650 382.950 539.850 389.400 ;
        RECT 544.650 388.500 545.850 392.400 ;
        RECT 540.750 387.600 545.850 388.500 ;
        RECT 549.150 389.400 550.950 395.250 ;
        RECT 552.150 392.400 553.950 395.250 ;
        RECT 556.950 393.300 558.750 395.250 ;
        RECT 555.000 392.400 558.750 393.300 ;
        RECT 561.450 392.400 563.250 395.250 ;
        RECT 564.750 392.400 566.550 395.250 ;
        RECT 568.650 392.400 570.450 395.250 ;
        RECT 572.850 392.400 574.650 395.250 ;
        RECT 577.350 392.400 579.150 395.250 ;
        RECT 555.000 391.500 556.050 392.400 ;
        RECT 553.950 389.400 556.050 391.500 ;
        RECT 564.750 390.600 565.800 392.400 ;
        RECT 540.750 386.700 543.000 387.600 ;
        RECT 454.950 377.850 457.050 379.950 ;
        RECT 455.250 376.050 457.050 377.850 ;
        RECT 458.850 375.600 460.050 380.850 ;
        RECT 464.100 379.050 465.900 380.850 ;
        RECT 411.150 374.400 412.050 375.300 ;
        RECT 408.450 374.100 410.250 374.400 ;
        RECT 395.550 372.600 396.750 373.500 ;
        RECT 403.950 373.200 410.250 374.100 ;
        RECT 408.450 372.600 410.250 373.200 ;
        RECT 411.150 372.600 413.850 374.400 ;
        RECT 391.950 370.500 396.750 372.600 ;
        RECT 399.150 370.500 406.050 372.300 ;
        RECT 395.550 369.600 396.750 370.500 ;
        RECT 390.150 363.750 391.950 369.600 ;
        RECT 395.250 363.750 397.050 369.600 ;
        RECT 400.050 363.750 401.850 369.600 ;
        RECT 403.050 363.750 404.850 370.500 ;
        RECT 411.150 369.600 415.050 371.700 ;
        RECT 406.950 363.750 408.750 369.600 ;
        RECT 411.150 363.750 412.950 369.600 ;
        RECT 415.650 363.750 417.450 366.600 ;
        RECT 418.650 363.750 420.450 375.600 ;
        RECT 455.400 363.750 457.200 369.600 ;
        RECT 458.700 363.750 460.500 375.600 ;
        RECT 462.900 363.750 464.700 375.600 ;
        RECT 500.400 369.600 501.600 382.050 ;
        RECT 538.650 380.850 541.050 382.950 ;
        RECT 538.650 375.600 539.850 380.850 ;
        RECT 541.950 378.300 543.000 386.700 ;
        RECT 544.950 380.850 547.050 382.950 ;
        RECT 545.100 379.050 546.900 380.850 ;
        RECT 540.750 377.400 543.000 378.300 ;
        RECT 540.750 376.500 546.450 377.400 ;
        RECT 499.650 363.750 501.450 369.600 ;
        RECT 502.650 363.750 504.450 369.600 ;
        RECT 538.350 363.750 540.150 375.600 ;
        RECT 541.350 363.750 543.150 375.600 ;
        RECT 545.250 369.600 546.450 376.500 ;
        RECT 544.650 363.750 546.450 369.600 ;
        RECT 549.150 376.800 550.050 389.400 ;
        RECT 557.550 388.800 559.350 390.600 ;
        RECT 560.850 389.550 565.800 390.600 ;
        RECT 573.300 391.500 574.350 392.400 ;
        RECT 573.300 390.300 577.050 391.500 ;
        RECT 560.850 388.800 562.650 389.550 ;
        RECT 557.850 387.900 558.900 388.800 ;
        RECT 568.050 388.200 569.850 390.000 ;
        RECT 574.950 389.400 577.050 390.300 ;
        RECT 580.650 389.400 582.450 395.250 ;
        RECT 614.550 392.400 616.350 395.250 ;
        RECT 568.050 387.900 568.950 388.200 ;
        RECT 557.850 387.000 568.950 387.900 ;
        RECT 581.250 387.150 582.450 389.400 ;
        RECT 615.150 388.500 616.350 392.400 ;
        RECT 617.850 389.400 619.650 395.250 ;
        RECT 620.850 389.400 622.650 395.250 ;
        RECT 627.150 389.400 628.950 395.250 ;
        RECT 630.150 392.400 631.950 395.250 ;
        RECT 634.950 393.300 636.750 395.250 ;
        RECT 633.000 392.400 636.750 393.300 ;
        RECT 639.450 392.400 641.250 395.250 ;
        RECT 642.750 392.400 644.550 395.250 ;
        RECT 646.650 392.400 648.450 395.250 ;
        RECT 650.850 392.400 652.650 395.250 ;
        RECT 655.350 392.400 657.150 395.250 ;
        RECT 633.000 391.500 634.050 392.400 ;
        RECT 631.950 389.400 634.050 391.500 ;
        RECT 642.750 390.600 643.800 392.400 ;
        RECT 615.150 387.600 620.250 388.500 ;
        RECT 557.850 385.800 558.900 387.000 ;
        RECT 552.000 384.600 558.900 385.800 ;
        RECT 552.000 383.850 552.900 384.600 ;
        RECT 557.100 384.000 558.900 384.600 ;
        RECT 551.100 382.050 552.900 383.850 ;
        RECT 554.100 382.950 555.900 383.700 ;
        RECT 568.050 382.950 568.950 387.000 ;
        RECT 577.950 385.050 582.450 387.150 ;
        RECT 576.150 383.250 580.050 385.050 ;
        RECT 577.950 382.950 580.050 383.250 ;
        RECT 554.100 381.900 562.050 382.950 ;
        RECT 559.950 380.850 562.050 381.900 ;
        RECT 565.950 380.850 568.950 382.950 ;
        RECT 558.450 377.100 560.250 377.400 ;
        RECT 558.450 376.800 566.850 377.100 ;
        RECT 549.150 376.200 566.850 376.800 ;
        RECT 549.150 375.600 560.250 376.200 ;
        RECT 549.150 363.750 550.950 375.600 ;
        RECT 563.250 374.700 565.050 375.300 ;
        RECT 557.550 373.500 565.050 374.700 ;
        RECT 565.950 374.100 566.850 376.200 ;
        RECT 568.050 376.200 568.950 380.850 ;
        RECT 578.250 377.400 580.050 379.200 ;
        RECT 574.950 376.200 579.150 377.400 ;
        RECT 568.050 375.300 574.050 376.200 ;
        RECT 574.950 375.300 577.050 376.200 ;
        RECT 581.250 375.600 582.450 385.050 ;
        RECT 618.000 386.700 620.250 387.600 ;
        RECT 613.950 380.850 616.050 382.950 ;
        RECT 614.100 379.050 615.900 380.850 ;
        RECT 618.000 378.300 619.050 386.700 ;
        RECT 621.150 382.950 622.350 389.400 ;
        RECT 619.950 380.850 622.350 382.950 ;
        RECT 618.000 377.400 620.250 378.300 ;
        RECT 573.150 374.400 574.050 375.300 ;
        RECT 570.450 374.100 572.250 374.400 ;
        RECT 557.550 372.600 558.750 373.500 ;
        RECT 565.950 373.200 572.250 374.100 ;
        RECT 570.450 372.600 572.250 373.200 ;
        RECT 573.150 372.600 575.850 374.400 ;
        RECT 553.950 370.500 558.750 372.600 ;
        RECT 561.150 370.500 568.050 372.300 ;
        RECT 557.550 369.600 558.750 370.500 ;
        RECT 552.150 363.750 553.950 369.600 ;
        RECT 557.250 363.750 559.050 369.600 ;
        RECT 562.050 363.750 563.850 369.600 ;
        RECT 565.050 363.750 566.850 370.500 ;
        RECT 573.150 369.600 577.050 371.700 ;
        RECT 568.950 363.750 570.750 369.600 ;
        RECT 573.150 363.750 574.950 369.600 ;
        RECT 577.650 363.750 579.450 366.600 ;
        RECT 580.650 363.750 582.450 375.600 ;
        RECT 614.550 376.500 620.250 377.400 ;
        RECT 614.550 369.600 615.750 376.500 ;
        RECT 621.150 375.600 622.350 380.850 ;
        RECT 627.150 376.800 628.050 389.400 ;
        RECT 635.550 388.800 637.350 390.600 ;
        RECT 638.850 389.550 643.800 390.600 ;
        RECT 651.300 391.500 652.350 392.400 ;
        RECT 651.300 390.300 655.050 391.500 ;
        RECT 638.850 388.800 640.650 389.550 ;
        RECT 635.850 387.900 636.900 388.800 ;
        RECT 646.050 388.200 647.850 390.000 ;
        RECT 652.950 389.400 655.050 390.300 ;
        RECT 658.650 389.400 660.450 395.250 ;
        RECT 692.550 392.400 694.350 395.250 ;
        RECT 695.550 392.400 697.350 395.250 ;
        RECT 646.050 387.900 646.950 388.200 ;
        RECT 635.850 387.000 646.950 387.900 ;
        RECT 659.250 387.150 660.450 389.400 ;
        RECT 635.850 385.800 636.900 387.000 ;
        RECT 630.000 384.600 636.900 385.800 ;
        RECT 630.000 383.850 630.900 384.600 ;
        RECT 635.100 384.000 636.900 384.600 ;
        RECT 629.100 382.050 630.900 383.850 ;
        RECT 632.100 382.950 633.900 383.700 ;
        RECT 646.050 382.950 646.950 387.000 ;
        RECT 655.950 385.050 660.450 387.150 ;
        RECT 654.150 383.250 658.050 385.050 ;
        RECT 655.950 382.950 658.050 383.250 ;
        RECT 632.100 381.900 640.050 382.950 ;
        RECT 637.950 380.850 640.050 381.900 ;
        RECT 643.950 380.850 646.950 382.950 ;
        RECT 636.450 377.100 638.250 377.400 ;
        RECT 636.450 376.800 644.850 377.100 ;
        RECT 627.150 376.200 644.850 376.800 ;
        RECT 627.150 375.600 638.250 376.200 ;
        RECT 614.550 363.750 616.350 369.600 ;
        RECT 617.850 363.750 619.650 375.600 ;
        RECT 620.850 363.750 622.650 375.600 ;
        RECT 627.150 363.750 628.950 375.600 ;
        RECT 641.250 374.700 643.050 375.300 ;
        RECT 635.550 373.500 643.050 374.700 ;
        RECT 643.950 374.100 644.850 376.200 ;
        RECT 646.050 376.200 646.950 380.850 ;
        RECT 656.250 377.400 658.050 379.200 ;
        RECT 652.950 376.200 657.150 377.400 ;
        RECT 646.050 375.300 652.050 376.200 ;
        RECT 652.950 375.300 655.050 376.200 ;
        RECT 659.250 375.600 660.450 385.050 ;
        RECT 691.950 383.850 694.050 385.950 ;
        RECT 695.400 384.150 696.600 392.400 ;
        RECT 733.650 389.400 735.450 395.250 ;
        RECT 734.250 387.300 735.450 389.400 ;
        RECT 736.650 390.300 738.450 395.250 ;
        RECT 739.650 391.200 741.450 395.250 ;
        RECT 742.650 390.300 744.450 395.250 ;
        RECT 736.650 388.950 744.450 390.300 ;
        RECT 734.250 386.250 738.000 387.300 ;
        RECT 692.100 382.050 693.900 383.850 ;
        RECT 694.950 382.050 697.050 384.150 ;
        RECT 736.950 382.950 738.150 386.250 ;
        RECT 740.100 384.150 741.900 385.950 ;
        RECT 651.150 374.400 652.050 375.300 ;
        RECT 648.450 374.100 650.250 374.400 ;
        RECT 635.550 372.600 636.750 373.500 ;
        RECT 643.950 373.200 650.250 374.100 ;
        RECT 648.450 372.600 650.250 373.200 ;
        RECT 651.150 372.600 653.850 374.400 ;
        RECT 631.950 370.500 636.750 372.600 ;
        RECT 639.150 370.500 646.050 372.300 ;
        RECT 635.550 369.600 636.750 370.500 ;
        RECT 630.150 363.750 631.950 369.600 ;
        RECT 635.250 363.750 637.050 369.600 ;
        RECT 640.050 363.750 641.850 369.600 ;
        RECT 643.050 363.750 644.850 370.500 ;
        RECT 651.150 369.600 655.050 371.700 ;
        RECT 646.950 363.750 648.750 369.600 ;
        RECT 651.150 363.750 652.950 369.600 ;
        RECT 655.650 363.750 657.450 366.600 ;
        RECT 658.650 363.750 660.450 375.600 ;
        RECT 695.400 369.600 696.600 382.050 ;
        RECT 736.950 380.850 739.050 382.950 ;
        RECT 739.950 382.050 742.050 384.150 ;
        RECT 742.950 380.850 745.050 382.950 ;
        RECT 733.950 377.850 736.050 379.950 ;
        RECT 734.250 376.050 736.050 377.850 ;
        RECT 737.850 375.600 739.050 380.850 ;
        RECT 743.100 379.050 744.900 380.850 ;
        RECT 692.550 363.750 694.350 369.600 ;
        RECT 695.550 363.750 697.350 369.600 ;
        RECT 734.400 363.750 736.200 369.600 ;
        RECT 737.700 363.750 739.500 375.600 ;
        RECT 741.900 363.750 743.700 375.600 ;
        RECT 3.150 347.400 4.950 359.250 ;
        RECT 6.150 353.400 7.950 359.250 ;
        RECT 11.250 353.400 13.050 359.250 ;
        RECT 16.050 353.400 17.850 359.250 ;
        RECT 11.550 352.500 12.750 353.400 ;
        RECT 19.050 352.500 20.850 359.250 ;
        RECT 22.950 353.400 24.750 359.250 ;
        RECT 27.150 353.400 28.950 359.250 ;
        RECT 31.650 356.400 33.450 359.250 ;
        RECT 7.950 350.400 12.750 352.500 ;
        RECT 15.150 350.700 22.050 352.500 ;
        RECT 27.150 351.300 31.050 353.400 ;
        RECT 11.550 349.500 12.750 350.400 ;
        RECT 24.450 349.800 26.250 350.400 ;
        RECT 11.550 348.300 19.050 349.500 ;
        RECT 17.250 347.700 19.050 348.300 ;
        RECT 19.950 348.900 26.250 349.800 ;
        RECT 3.150 346.800 14.250 347.400 ;
        RECT 19.950 346.800 20.850 348.900 ;
        RECT 24.450 348.600 26.250 348.900 ;
        RECT 27.150 348.600 29.850 350.400 ;
        RECT 27.150 347.700 28.050 348.600 ;
        RECT 3.150 346.200 20.850 346.800 ;
        RECT 3.150 333.600 4.050 346.200 ;
        RECT 12.450 345.900 20.850 346.200 ;
        RECT 22.050 346.800 28.050 347.700 ;
        RECT 28.950 346.800 31.050 347.700 ;
        RECT 34.650 347.400 36.450 359.250 ;
        RECT 71.400 353.400 73.200 359.250 ;
        RECT 74.700 347.400 76.500 359.250 ;
        RECT 78.900 347.400 80.700 359.250 ;
        RECT 114.300 347.400 116.100 359.250 ;
        RECT 118.500 347.400 120.300 359.250 ;
        RECT 121.800 353.400 123.600 359.250 ;
        RECT 157.650 353.400 159.450 359.250 ;
        RECT 160.650 353.400 162.450 359.250 ;
        RECT 163.650 353.400 165.450 359.250 ;
        RECT 197.550 353.400 199.350 359.250 ;
        RECT 200.550 353.400 202.350 359.250 ;
        RECT 239.400 353.400 241.200 359.250 ;
        RECT 12.450 345.600 14.250 345.900 ;
        RECT 22.050 342.150 22.950 346.800 ;
        RECT 28.950 345.600 33.150 346.800 ;
        RECT 32.250 343.800 34.050 345.600 ;
        RECT 13.950 341.100 16.050 342.150 ;
        RECT 5.100 339.150 6.900 340.950 ;
        RECT 8.100 340.050 16.050 341.100 ;
        RECT 19.950 340.050 22.950 342.150 ;
        RECT 8.100 339.300 9.900 340.050 ;
        RECT 6.000 338.400 6.900 339.150 ;
        RECT 11.100 338.400 12.900 339.000 ;
        RECT 6.000 337.200 12.900 338.400 ;
        RECT 11.850 336.000 12.900 337.200 ;
        RECT 22.050 336.000 22.950 340.050 ;
        RECT 31.950 339.750 34.050 340.050 ;
        RECT 30.150 337.950 34.050 339.750 ;
        RECT 35.250 337.950 36.450 347.400 ;
        RECT 71.250 345.150 73.050 346.950 ;
        RECT 70.950 343.050 73.050 345.150 ;
        RECT 74.850 342.150 76.050 347.400 ;
        RECT 80.100 342.150 81.900 343.950 ;
        RECT 113.100 342.150 114.900 343.950 ;
        RECT 118.950 342.150 120.150 347.400 ;
        RECT 121.950 345.150 123.750 346.950 ;
        RECT 161.250 345.150 162.450 353.400 ;
        RECT 121.950 343.050 124.050 345.150 ;
        RECT 11.850 335.100 22.950 336.000 ;
        RECT 31.950 335.850 36.450 337.950 ;
        RECT 73.950 340.050 76.050 342.150 ;
        RECT 73.950 336.750 75.150 340.050 ;
        RECT 76.950 338.850 79.050 340.950 ;
        RECT 79.950 340.050 82.050 342.150 ;
        RECT 112.950 340.050 115.050 342.150 ;
        RECT 115.950 338.850 118.050 340.950 ;
        RECT 118.950 340.050 121.050 342.150 ;
        RECT 157.950 341.850 160.050 343.950 ;
        RECT 160.950 343.050 163.050 345.150 ;
        RECT 158.100 340.050 159.900 341.850 ;
        RECT 77.100 337.050 78.900 338.850 ;
        RECT 116.100 337.050 117.900 338.850 ;
        RECT 119.850 336.750 121.050 340.050 ;
        RECT 11.850 334.200 12.900 335.100 ;
        RECT 22.050 334.800 22.950 335.100 ;
        RECT 3.150 327.750 4.950 333.600 ;
        RECT 7.950 331.500 10.050 333.600 ;
        RECT 11.550 332.400 13.350 334.200 ;
        RECT 14.850 333.450 16.650 334.200 ;
        RECT 14.850 332.400 19.800 333.450 ;
        RECT 22.050 333.000 23.850 334.800 ;
        RECT 35.250 333.600 36.450 335.850 ;
        RECT 71.250 335.700 75.000 336.750 ;
        RECT 120.000 335.700 123.750 336.750 ;
        RECT 161.250 335.700 162.450 343.050 ;
        RECT 163.950 341.850 166.050 343.950 ;
        RECT 164.100 340.050 165.900 341.850 ;
        RECT 200.400 340.950 201.600 353.400 ;
        RECT 242.700 347.400 244.500 359.250 ;
        RECT 246.900 347.400 248.700 359.250 ;
        RECT 281.550 353.400 283.350 359.250 ;
        RECT 284.550 353.400 286.350 359.250 ;
        RECT 287.550 353.400 289.350 359.250 ;
        RECT 239.250 345.150 241.050 346.950 ;
        RECT 238.950 343.050 241.050 345.150 ;
        RECT 242.850 342.150 244.050 347.400 ;
        RECT 284.550 345.150 285.750 353.400 ;
        RECT 294.150 347.400 295.950 359.250 ;
        RECT 297.150 353.400 298.950 359.250 ;
        RECT 302.250 353.400 304.050 359.250 ;
        RECT 307.050 353.400 308.850 359.250 ;
        RECT 302.550 352.500 303.750 353.400 ;
        RECT 310.050 352.500 311.850 359.250 ;
        RECT 313.950 353.400 315.750 359.250 ;
        RECT 318.150 353.400 319.950 359.250 ;
        RECT 322.650 356.400 324.450 359.250 ;
        RECT 298.950 350.400 303.750 352.500 ;
        RECT 306.150 350.700 313.050 352.500 ;
        RECT 318.150 351.300 322.050 353.400 ;
        RECT 302.550 349.500 303.750 350.400 ;
        RECT 315.450 349.800 317.250 350.400 ;
        RECT 302.550 348.300 310.050 349.500 ;
        RECT 308.250 347.700 310.050 348.300 ;
        RECT 310.950 348.900 317.250 349.800 ;
        RECT 294.150 346.800 305.250 347.400 ;
        RECT 310.950 346.800 311.850 348.900 ;
        RECT 315.450 348.600 317.250 348.900 ;
        RECT 318.150 348.600 320.850 350.400 ;
        RECT 318.150 347.700 319.050 348.600 ;
        RECT 294.150 346.200 311.850 346.800 ;
        RECT 248.100 342.150 249.900 343.950 ;
        RECT 197.100 339.150 198.900 340.950 ;
        RECT 196.950 337.050 199.050 339.150 ;
        RECT 199.950 338.850 202.050 340.950 ;
        RECT 241.950 340.050 244.050 342.150 ;
        RECT 71.250 333.600 72.450 335.700 ;
        RECT 28.950 332.700 31.050 333.600 ;
        RECT 9.000 330.600 10.050 331.500 ;
        RECT 18.750 330.600 19.800 332.400 ;
        RECT 27.300 331.500 31.050 332.700 ;
        RECT 27.300 330.600 28.350 331.500 ;
        RECT 6.150 327.750 7.950 330.600 ;
        RECT 9.000 329.700 12.750 330.600 ;
        RECT 10.950 327.750 12.750 329.700 ;
        RECT 15.450 327.750 17.250 330.600 ;
        RECT 18.750 327.750 20.550 330.600 ;
        RECT 22.650 327.750 24.450 330.600 ;
        RECT 26.850 327.750 28.650 330.600 ;
        RECT 31.350 327.750 33.150 330.600 ;
        RECT 34.650 327.750 36.450 333.600 ;
        RECT 70.650 327.750 72.450 333.600 ;
        RECT 73.650 332.700 81.450 334.050 ;
        RECT 73.650 327.750 75.450 332.700 ;
        RECT 76.650 327.750 78.450 331.800 ;
        RECT 79.650 327.750 81.450 332.700 ;
        RECT 113.550 332.700 121.350 334.050 ;
        RECT 113.550 327.750 115.350 332.700 ;
        RECT 116.550 327.750 118.350 331.800 ;
        RECT 119.550 327.750 121.350 332.700 ;
        RECT 122.550 333.600 123.750 335.700 ;
        RECT 158.850 334.800 162.450 335.700 ;
        RECT 122.550 327.750 124.350 333.600 ;
        RECT 158.850 327.750 160.650 334.800 ;
        RECT 163.350 327.750 165.150 333.600 ;
        RECT 200.400 330.600 201.600 338.850 ;
        RECT 241.950 336.750 243.150 340.050 ;
        RECT 244.950 338.850 247.050 340.950 ;
        RECT 247.950 340.050 250.050 342.150 ;
        RECT 280.950 341.850 283.050 343.950 ;
        RECT 283.950 343.050 286.050 345.150 ;
        RECT 281.100 340.050 282.900 341.850 ;
        RECT 245.100 337.050 246.900 338.850 ;
        RECT 239.250 335.700 243.000 336.750 ;
        RECT 284.550 335.700 285.750 343.050 ;
        RECT 286.950 341.850 289.050 343.950 ;
        RECT 287.100 340.050 288.900 341.850 ;
        RECT 239.250 333.600 240.450 335.700 ;
        RECT 284.550 334.800 288.150 335.700 ;
        RECT 197.550 327.750 199.350 330.600 ;
        RECT 200.550 327.750 202.350 330.600 ;
        RECT 238.650 327.750 240.450 333.600 ;
        RECT 241.650 332.700 249.450 334.050 ;
        RECT 241.650 327.750 243.450 332.700 ;
        RECT 244.650 327.750 246.450 331.800 ;
        RECT 247.650 327.750 249.450 332.700 ;
        RECT 281.850 327.750 283.650 333.600 ;
        RECT 286.350 327.750 288.150 334.800 ;
        RECT 294.150 333.600 295.050 346.200 ;
        RECT 303.450 345.900 311.850 346.200 ;
        RECT 313.050 346.800 319.050 347.700 ;
        RECT 319.950 346.800 322.050 347.700 ;
        RECT 325.650 347.400 327.450 359.250 ;
        RECT 361.650 353.400 363.450 359.250 ;
        RECT 364.650 354.000 366.450 359.250 ;
        RECT 303.450 345.600 305.250 345.900 ;
        RECT 313.050 342.150 313.950 346.800 ;
        RECT 319.950 345.600 324.150 346.800 ;
        RECT 323.250 343.800 325.050 345.600 ;
        RECT 304.950 341.100 307.050 342.150 ;
        RECT 296.100 339.150 297.900 340.950 ;
        RECT 299.100 340.050 307.050 341.100 ;
        RECT 310.950 340.050 313.950 342.150 ;
        RECT 299.100 339.300 300.900 340.050 ;
        RECT 297.000 338.400 297.900 339.150 ;
        RECT 302.100 338.400 303.900 339.000 ;
        RECT 297.000 337.200 303.900 338.400 ;
        RECT 302.850 336.000 303.900 337.200 ;
        RECT 313.050 336.000 313.950 340.050 ;
        RECT 322.950 339.750 325.050 340.050 ;
        RECT 321.150 337.950 325.050 339.750 ;
        RECT 326.250 337.950 327.450 347.400 ;
        RECT 362.250 353.100 363.450 353.400 ;
        RECT 367.650 353.400 369.450 359.250 ;
        RECT 370.650 353.400 372.450 359.250 ;
        RECT 404.550 353.400 406.350 359.250 ;
        RECT 407.550 353.400 409.350 359.250 ;
        RECT 410.550 354.000 412.350 359.250 ;
        RECT 367.650 353.100 369.300 353.400 ;
        RECT 362.250 352.200 369.300 353.100 ;
        RECT 407.700 353.100 409.350 353.400 ;
        RECT 413.550 353.400 415.350 359.250 ;
        RECT 413.550 353.100 414.750 353.400 ;
        RECT 407.700 352.200 414.750 353.100 ;
        RECT 362.250 343.950 363.300 352.200 ;
        RECT 368.100 348.150 369.900 349.950 ;
        RECT 407.100 348.150 408.900 349.950 ;
        RECT 364.950 345.150 366.750 346.950 ;
        RECT 367.950 346.050 370.050 348.150 ;
        RECT 371.100 345.150 372.900 346.950 ;
        RECT 404.100 345.150 405.900 346.950 ;
        RECT 406.950 346.050 409.050 348.150 ;
        RECT 410.250 345.150 412.050 346.950 ;
        RECT 361.950 341.850 364.050 343.950 ;
        RECT 364.950 343.050 367.050 345.150 ;
        RECT 370.950 343.050 373.050 345.150 ;
        RECT 403.950 343.050 406.050 345.150 ;
        RECT 409.950 343.050 412.050 345.150 ;
        RECT 413.700 343.950 414.750 352.200 ;
        RECT 419.550 347.400 421.350 359.250 ;
        RECT 422.550 356.400 424.350 359.250 ;
        RECT 427.050 353.400 428.850 359.250 ;
        RECT 431.250 353.400 433.050 359.250 ;
        RECT 424.950 351.300 428.850 353.400 ;
        RECT 435.150 352.500 436.950 359.250 ;
        RECT 438.150 353.400 439.950 359.250 ;
        RECT 442.950 353.400 444.750 359.250 ;
        RECT 448.050 353.400 449.850 359.250 ;
        RECT 443.250 352.500 444.450 353.400 ;
        RECT 433.950 350.700 440.850 352.500 ;
        RECT 443.250 350.400 448.050 352.500 ;
        RECT 426.150 348.600 428.850 350.400 ;
        RECT 429.750 349.800 431.550 350.400 ;
        RECT 429.750 348.900 436.050 349.800 ;
        RECT 443.250 349.500 444.450 350.400 ;
        RECT 429.750 348.600 431.550 348.900 ;
        RECT 427.950 347.700 428.850 348.600 ;
        RECT 412.950 341.850 415.050 343.950 ;
        RECT 302.850 335.100 313.950 336.000 ;
        RECT 322.950 335.850 327.450 337.950 ;
        RECT 362.400 337.650 363.600 341.850 ;
        RECT 413.400 337.650 414.600 341.850 ;
        RECT 362.400 336.000 366.900 337.650 ;
        RECT 302.850 334.200 303.900 335.100 ;
        RECT 313.050 334.800 313.950 335.100 ;
        RECT 294.150 327.750 295.950 333.600 ;
        RECT 298.950 331.500 301.050 333.600 ;
        RECT 302.550 332.400 304.350 334.200 ;
        RECT 305.850 333.450 307.650 334.200 ;
        RECT 305.850 332.400 310.800 333.450 ;
        RECT 313.050 333.000 314.850 334.800 ;
        RECT 326.250 333.600 327.450 335.850 ;
        RECT 319.950 332.700 322.050 333.600 ;
        RECT 300.000 330.600 301.050 331.500 ;
        RECT 309.750 330.600 310.800 332.400 ;
        RECT 318.300 331.500 322.050 332.700 ;
        RECT 318.300 330.600 319.350 331.500 ;
        RECT 297.150 327.750 298.950 330.600 ;
        RECT 300.000 329.700 303.750 330.600 ;
        RECT 301.950 327.750 303.750 329.700 ;
        RECT 306.450 327.750 308.250 330.600 ;
        RECT 309.750 327.750 311.550 330.600 ;
        RECT 313.650 327.750 315.450 330.600 ;
        RECT 317.850 327.750 319.650 330.600 ;
        RECT 322.350 327.750 324.150 330.600 ;
        RECT 325.650 327.750 327.450 333.600 ;
        RECT 365.100 327.750 366.900 336.000 ;
        RECT 370.500 327.750 372.300 336.600 ;
        RECT 404.700 327.750 406.500 336.600 ;
        RECT 410.100 336.000 414.600 337.650 ;
        RECT 419.550 337.950 420.750 347.400 ;
        RECT 424.950 346.800 427.050 347.700 ;
        RECT 427.950 346.800 433.950 347.700 ;
        RECT 422.850 345.600 427.050 346.800 ;
        RECT 421.950 343.800 423.750 345.600 ;
        RECT 433.050 342.150 433.950 346.800 ;
        RECT 435.150 346.800 436.050 348.900 ;
        RECT 436.950 348.300 444.450 349.500 ;
        RECT 436.950 347.700 438.750 348.300 ;
        RECT 451.050 347.400 452.850 359.250 ;
        RECT 488.400 353.400 490.200 359.250 ;
        RECT 491.700 347.400 493.500 359.250 ;
        RECT 495.900 347.400 497.700 359.250 ;
        RECT 501.150 347.400 502.950 359.250 ;
        RECT 504.150 353.400 505.950 359.250 ;
        RECT 509.250 353.400 511.050 359.250 ;
        RECT 514.050 353.400 515.850 359.250 ;
        RECT 509.550 352.500 510.750 353.400 ;
        RECT 517.050 352.500 518.850 359.250 ;
        RECT 520.950 353.400 522.750 359.250 ;
        RECT 525.150 353.400 526.950 359.250 ;
        RECT 529.650 356.400 531.450 359.250 ;
        RECT 505.950 350.400 510.750 352.500 ;
        RECT 513.150 350.700 520.050 352.500 ;
        RECT 525.150 351.300 529.050 353.400 ;
        RECT 509.550 349.500 510.750 350.400 ;
        RECT 522.450 349.800 524.250 350.400 ;
        RECT 509.550 348.300 517.050 349.500 ;
        RECT 515.250 347.700 517.050 348.300 ;
        RECT 517.950 348.900 524.250 349.800 ;
        RECT 441.750 346.800 452.850 347.400 ;
        RECT 435.150 346.200 452.850 346.800 ;
        RECT 435.150 345.900 443.550 346.200 ;
        RECT 441.750 345.600 443.550 345.900 ;
        RECT 433.050 340.050 436.050 342.150 ;
        RECT 439.950 341.100 442.050 342.150 ;
        RECT 439.950 340.050 447.900 341.100 ;
        RECT 421.950 339.750 424.050 340.050 ;
        RECT 421.950 337.950 425.850 339.750 ;
        RECT 410.100 327.750 411.900 336.000 ;
        RECT 419.550 335.850 424.050 337.950 ;
        RECT 433.050 336.000 433.950 340.050 ;
        RECT 446.100 339.300 447.900 340.050 ;
        RECT 449.100 339.150 450.900 340.950 ;
        RECT 443.100 338.400 444.900 339.000 ;
        RECT 449.100 338.400 450.000 339.150 ;
        RECT 443.100 337.200 450.000 338.400 ;
        RECT 443.100 336.000 444.150 337.200 ;
        RECT 419.550 333.600 420.750 335.850 ;
        RECT 433.050 335.100 444.150 336.000 ;
        RECT 433.050 334.800 433.950 335.100 ;
        RECT 419.550 327.750 421.350 333.600 ;
        RECT 424.950 332.700 427.050 333.600 ;
        RECT 432.150 333.000 433.950 334.800 ;
        RECT 443.100 334.200 444.150 335.100 ;
        RECT 439.350 333.450 441.150 334.200 ;
        RECT 424.950 331.500 428.700 332.700 ;
        RECT 427.650 330.600 428.700 331.500 ;
        RECT 436.200 332.400 441.150 333.450 ;
        RECT 442.650 332.400 444.450 334.200 ;
        RECT 451.950 333.600 452.850 346.200 ;
        RECT 488.250 345.150 490.050 346.950 ;
        RECT 487.950 343.050 490.050 345.150 ;
        RECT 491.850 342.150 493.050 347.400 ;
        RECT 501.150 346.800 512.250 347.400 ;
        RECT 517.950 346.800 518.850 348.900 ;
        RECT 522.450 348.600 524.250 348.900 ;
        RECT 525.150 348.600 527.850 350.400 ;
        RECT 525.150 347.700 526.050 348.600 ;
        RECT 501.150 346.200 518.850 346.800 ;
        RECT 497.100 342.150 498.900 343.950 ;
        RECT 490.950 340.050 493.050 342.150 ;
        RECT 490.950 336.750 492.150 340.050 ;
        RECT 493.950 338.850 496.050 340.950 ;
        RECT 496.950 340.050 499.050 342.150 ;
        RECT 494.100 337.050 495.900 338.850 ;
        RECT 488.250 335.700 492.000 336.750 ;
        RECT 488.250 333.600 489.450 335.700 ;
        RECT 436.200 330.600 437.250 332.400 ;
        RECT 445.950 331.500 448.050 333.600 ;
        RECT 445.950 330.600 447.000 331.500 ;
        RECT 422.850 327.750 424.650 330.600 ;
        RECT 427.350 327.750 429.150 330.600 ;
        RECT 431.550 327.750 433.350 330.600 ;
        RECT 435.450 327.750 437.250 330.600 ;
        RECT 438.750 327.750 440.550 330.600 ;
        RECT 443.250 329.700 447.000 330.600 ;
        RECT 443.250 327.750 445.050 329.700 ;
        RECT 448.050 327.750 449.850 330.600 ;
        RECT 451.050 327.750 452.850 333.600 ;
        RECT 487.650 327.750 489.450 333.600 ;
        RECT 490.650 332.700 498.450 334.050 ;
        RECT 490.650 327.750 492.450 332.700 ;
        RECT 493.650 327.750 495.450 331.800 ;
        RECT 496.650 327.750 498.450 332.700 ;
        RECT 501.150 333.600 502.050 346.200 ;
        RECT 510.450 345.900 518.850 346.200 ;
        RECT 520.050 346.800 526.050 347.700 ;
        RECT 526.950 346.800 529.050 347.700 ;
        RECT 532.650 347.400 534.450 359.250 ;
        RECT 566.550 347.400 568.350 359.250 ;
        RECT 510.450 345.600 512.250 345.900 ;
        RECT 520.050 342.150 520.950 346.800 ;
        RECT 526.950 345.600 531.150 346.800 ;
        RECT 530.250 343.800 532.050 345.600 ;
        RECT 511.950 341.100 514.050 342.150 ;
        RECT 503.100 339.150 504.900 340.950 ;
        RECT 506.100 340.050 514.050 341.100 ;
        RECT 517.950 340.050 520.950 342.150 ;
        RECT 506.100 339.300 507.900 340.050 ;
        RECT 504.000 338.400 504.900 339.150 ;
        RECT 509.100 338.400 510.900 339.000 ;
        RECT 504.000 337.200 510.900 338.400 ;
        RECT 509.850 336.000 510.900 337.200 ;
        RECT 520.050 336.000 520.950 340.050 ;
        RECT 529.950 339.750 532.050 340.050 ;
        RECT 528.150 337.950 532.050 339.750 ;
        RECT 533.250 337.950 534.450 347.400 ;
        RECT 569.550 346.500 571.350 359.250 ;
        RECT 572.550 347.400 574.350 359.250 ;
        RECT 575.550 346.500 577.350 359.250 ;
        RECT 578.550 347.400 580.350 359.250 ;
        RECT 581.550 346.500 583.350 359.250 ;
        RECT 584.550 347.400 586.350 359.250 ;
        RECT 587.550 346.500 589.350 359.250 ;
        RECT 590.550 347.400 592.350 359.250 ;
        RECT 628.650 353.400 630.450 359.250 ;
        RECT 631.650 353.400 633.450 359.250 ;
        RECT 634.650 353.400 636.450 359.250 ;
        RECT 610.950 348.450 613.050 349.050 ;
        RECT 628.950 348.450 631.050 349.050 ;
        RECT 610.950 347.550 631.050 348.450 ;
        RECT 610.950 346.950 613.050 347.550 ;
        RECT 628.950 346.950 631.050 347.550 ;
        RECT 569.550 345.300 573.450 346.500 ;
        RECT 575.550 345.300 579.300 346.500 ;
        RECT 581.550 345.300 585.300 346.500 ;
        RECT 587.550 345.300 590.250 346.500 ;
        RECT 568.950 338.850 571.050 340.950 ;
        RECT 509.850 335.100 520.950 336.000 ;
        RECT 529.950 335.850 534.450 337.950 ;
        RECT 569.100 337.050 570.900 338.850 ;
        RECT 572.250 338.400 573.450 345.300 ;
        RECT 578.100 338.400 579.300 345.300 ;
        RECT 584.100 338.400 585.300 345.300 ;
        RECT 589.200 340.950 590.250 345.300 ;
        RECT 632.250 345.150 633.450 353.400 ;
        RECT 638.550 347.400 640.350 359.250 ;
        RECT 641.550 356.400 643.350 359.250 ;
        RECT 646.050 353.400 647.850 359.250 ;
        RECT 650.250 353.400 652.050 359.250 ;
        RECT 643.950 351.300 647.850 353.400 ;
        RECT 654.150 352.500 655.950 359.250 ;
        RECT 657.150 353.400 658.950 359.250 ;
        RECT 661.950 353.400 663.750 359.250 ;
        RECT 667.050 353.400 668.850 359.250 ;
        RECT 662.250 352.500 663.450 353.400 ;
        RECT 652.950 350.700 659.850 352.500 ;
        RECT 662.250 350.400 667.050 352.500 ;
        RECT 645.150 348.600 647.850 350.400 ;
        RECT 648.750 349.800 650.550 350.400 ;
        RECT 648.750 348.900 655.050 349.800 ;
        RECT 662.250 349.500 663.450 350.400 ;
        RECT 648.750 348.600 650.550 348.900 ;
        RECT 646.950 347.700 647.850 348.600 ;
        RECT 628.950 341.850 631.050 343.950 ;
        RECT 631.950 343.050 634.050 345.150 ;
        RECT 589.200 338.850 592.050 340.950 ;
        RECT 629.100 340.050 630.900 341.850 ;
        RECT 509.850 334.200 510.900 335.100 ;
        RECT 520.050 334.800 520.950 335.100 ;
        RECT 501.150 327.750 502.950 333.600 ;
        RECT 505.950 331.500 508.050 333.600 ;
        RECT 509.550 332.400 511.350 334.200 ;
        RECT 512.850 333.450 514.650 334.200 ;
        RECT 512.850 332.400 517.800 333.450 ;
        RECT 520.050 333.000 521.850 334.800 ;
        RECT 533.250 333.600 534.450 335.850 ;
        RECT 572.250 336.600 576.300 338.400 ;
        RECT 578.100 336.600 582.300 338.400 ;
        RECT 584.100 336.600 588.300 338.400 ;
        RECT 572.250 335.700 573.450 336.600 ;
        RECT 578.100 335.700 579.300 336.600 ;
        RECT 584.100 335.700 585.300 336.600 ;
        RECT 589.200 335.700 590.250 338.850 ;
        RECT 632.250 335.700 633.450 343.050 ;
        RECT 634.950 341.850 637.050 343.950 ;
        RECT 635.100 340.050 636.900 341.850 ;
        RECT 569.400 334.500 573.450 335.700 ;
        RECT 575.550 334.500 579.300 335.700 ;
        RECT 581.400 334.500 585.300 335.700 ;
        RECT 587.400 334.650 590.250 335.700 ;
        RECT 629.850 334.800 633.450 335.700 ;
        RECT 638.550 337.950 639.750 347.400 ;
        RECT 643.950 346.800 646.050 347.700 ;
        RECT 646.950 346.800 652.950 347.700 ;
        RECT 641.850 345.600 646.050 346.800 ;
        RECT 640.950 343.800 642.750 345.600 ;
        RECT 652.050 342.150 652.950 346.800 ;
        RECT 654.150 346.800 655.050 348.900 ;
        RECT 655.950 348.300 663.450 349.500 ;
        RECT 655.950 347.700 657.750 348.300 ;
        RECT 670.050 347.400 671.850 359.250 ;
        RECT 706.650 353.400 708.450 359.250 ;
        RECT 709.650 353.400 711.450 359.250 ;
        RECT 712.650 353.400 714.450 359.250 ;
        RECT 660.750 346.800 671.850 347.400 ;
        RECT 654.150 346.200 671.850 346.800 ;
        RECT 654.150 345.900 662.550 346.200 ;
        RECT 660.750 345.600 662.550 345.900 ;
        RECT 652.050 340.050 655.050 342.150 ;
        RECT 658.950 341.100 661.050 342.150 ;
        RECT 658.950 340.050 666.900 341.100 ;
        RECT 640.950 339.750 643.050 340.050 ;
        RECT 640.950 337.950 644.850 339.750 ;
        RECT 638.550 335.850 643.050 337.950 ;
        RECT 652.050 336.000 652.950 340.050 ;
        RECT 665.100 339.300 666.900 340.050 ;
        RECT 668.100 339.150 669.900 340.950 ;
        RECT 662.100 338.400 663.900 339.000 ;
        RECT 668.100 338.400 669.000 339.150 ;
        RECT 662.100 337.200 669.000 338.400 ;
        RECT 662.100 336.000 663.150 337.200 ;
        RECT 587.400 334.500 590.100 334.650 ;
        RECT 569.400 333.600 571.200 334.500 ;
        RECT 526.950 332.700 529.050 333.600 ;
        RECT 507.000 330.600 508.050 331.500 ;
        RECT 516.750 330.600 517.800 332.400 ;
        RECT 525.300 331.500 529.050 332.700 ;
        RECT 525.300 330.600 526.350 331.500 ;
        RECT 504.150 327.750 505.950 330.600 ;
        RECT 507.000 329.700 510.750 330.600 ;
        RECT 508.950 327.750 510.750 329.700 ;
        RECT 513.450 327.750 515.250 330.600 ;
        RECT 516.750 327.750 518.550 330.600 ;
        RECT 520.650 327.750 522.450 330.600 ;
        RECT 524.850 327.750 526.650 330.600 ;
        RECT 529.350 327.750 531.150 330.600 ;
        RECT 532.650 327.750 534.450 333.600 ;
        RECT 566.550 327.750 568.350 333.600 ;
        RECT 569.550 327.750 571.350 333.600 ;
        RECT 572.550 327.750 574.350 333.600 ;
        RECT 575.550 327.750 577.350 334.500 ;
        RECT 581.400 333.600 583.200 334.500 ;
        RECT 587.400 333.600 589.200 334.500 ;
        RECT 578.550 327.750 580.350 333.600 ;
        RECT 581.550 327.750 583.350 333.600 ;
        RECT 584.550 327.750 586.350 333.600 ;
        RECT 587.550 327.750 589.350 333.600 ;
        RECT 590.550 327.750 592.350 333.600 ;
        RECT 629.850 327.750 631.650 334.800 ;
        RECT 638.550 333.600 639.750 335.850 ;
        RECT 652.050 335.100 663.150 336.000 ;
        RECT 652.050 334.800 652.950 335.100 ;
        RECT 634.350 327.750 636.150 333.600 ;
        RECT 638.550 327.750 640.350 333.600 ;
        RECT 643.950 332.700 646.050 333.600 ;
        RECT 651.150 333.000 652.950 334.800 ;
        RECT 662.100 334.200 663.150 335.100 ;
        RECT 658.350 333.450 660.150 334.200 ;
        RECT 643.950 331.500 647.700 332.700 ;
        RECT 646.650 330.600 647.700 331.500 ;
        RECT 655.200 332.400 660.150 333.450 ;
        RECT 661.650 332.400 663.450 334.200 ;
        RECT 670.950 333.600 671.850 346.200 ;
        RECT 710.250 345.150 711.450 353.400 ;
        RECT 747.300 347.400 749.100 359.250 ;
        RECT 751.500 347.400 753.300 359.250 ;
        RECT 754.800 353.400 756.600 359.250 ;
        RECT 706.950 341.850 709.050 343.950 ;
        RECT 709.950 343.050 712.050 345.150 ;
        RECT 707.100 340.050 708.900 341.850 ;
        RECT 710.250 335.700 711.450 343.050 ;
        RECT 712.950 341.850 715.050 343.950 ;
        RECT 746.100 342.150 747.900 343.950 ;
        RECT 751.950 342.150 753.150 347.400 ;
        RECT 754.950 345.150 756.750 346.950 ;
        RECT 754.950 343.050 757.050 345.150 ;
        RECT 713.100 340.050 714.900 341.850 ;
        RECT 745.950 340.050 748.050 342.150 ;
        RECT 748.950 338.850 751.050 340.950 ;
        RECT 751.950 340.050 754.050 342.150 ;
        RECT 749.100 337.050 750.900 338.850 ;
        RECT 752.850 336.750 754.050 340.050 ;
        RECT 753.000 335.700 756.750 336.750 ;
        RECT 655.200 330.600 656.250 332.400 ;
        RECT 664.950 331.500 667.050 333.600 ;
        RECT 664.950 330.600 666.000 331.500 ;
        RECT 641.850 327.750 643.650 330.600 ;
        RECT 646.350 327.750 648.150 330.600 ;
        RECT 650.550 327.750 652.350 330.600 ;
        RECT 654.450 327.750 656.250 330.600 ;
        RECT 657.750 327.750 659.550 330.600 ;
        RECT 662.250 329.700 666.000 330.600 ;
        RECT 662.250 327.750 664.050 329.700 ;
        RECT 667.050 327.750 668.850 330.600 ;
        RECT 670.050 327.750 671.850 333.600 ;
        RECT 707.850 334.800 711.450 335.700 ;
        RECT 707.850 327.750 709.650 334.800 ;
        RECT 712.350 327.750 714.150 333.600 ;
        RECT 746.550 332.700 754.350 334.050 ;
        RECT 746.550 327.750 748.350 332.700 ;
        RECT 749.550 327.750 751.350 331.800 ;
        RECT 752.550 327.750 754.350 332.700 ;
        RECT 755.550 333.600 756.750 335.700 ;
        RECT 755.550 327.750 757.350 333.600 ;
        RECT 3.150 317.400 4.950 323.250 ;
        RECT 6.150 320.400 7.950 323.250 ;
        RECT 10.950 321.300 12.750 323.250 ;
        RECT 9.000 320.400 12.750 321.300 ;
        RECT 15.450 320.400 17.250 323.250 ;
        RECT 18.750 320.400 20.550 323.250 ;
        RECT 22.650 320.400 24.450 323.250 ;
        RECT 26.850 320.400 28.650 323.250 ;
        RECT 31.350 320.400 33.150 323.250 ;
        RECT 9.000 319.500 10.050 320.400 ;
        RECT 7.950 317.400 10.050 319.500 ;
        RECT 18.750 318.600 19.800 320.400 ;
        RECT 3.150 304.800 4.050 317.400 ;
        RECT 11.550 316.800 13.350 318.600 ;
        RECT 14.850 317.550 19.800 318.600 ;
        RECT 27.300 319.500 28.350 320.400 ;
        RECT 27.300 318.300 31.050 319.500 ;
        RECT 14.850 316.800 16.650 317.550 ;
        RECT 11.850 315.900 12.900 316.800 ;
        RECT 22.050 316.200 23.850 318.000 ;
        RECT 28.950 317.400 31.050 318.300 ;
        RECT 34.650 317.400 36.450 323.250 ;
        RECT 65.550 320.400 67.350 323.250 ;
        RECT 68.550 320.400 70.350 323.250 ;
        RECT 71.550 320.400 73.350 323.250 ;
        RECT 22.050 315.900 22.950 316.200 ;
        RECT 11.850 315.000 22.950 315.900 ;
        RECT 35.250 315.150 36.450 317.400 ;
        RECT 69.450 316.200 70.350 320.400 ;
        RECT 74.550 317.400 76.350 323.250 ;
        RECT 112.350 317.400 114.150 323.250 ;
        RECT 115.350 317.400 117.150 323.250 ;
        RECT 118.650 320.400 120.450 323.250 ;
        RECT 69.450 315.300 72.750 316.200 ;
        RECT 11.850 313.800 12.900 315.000 ;
        RECT 6.000 312.600 12.900 313.800 ;
        RECT 6.000 311.850 6.900 312.600 ;
        RECT 11.100 312.000 12.900 312.600 ;
        RECT 5.100 310.050 6.900 311.850 ;
        RECT 8.100 310.950 9.900 311.700 ;
        RECT 22.050 310.950 22.950 315.000 ;
        RECT 31.950 313.050 36.450 315.150 ;
        RECT 70.950 314.400 72.750 315.300 ;
        RECT 30.150 311.250 34.050 313.050 ;
        RECT 31.950 310.950 34.050 311.250 ;
        RECT 8.100 309.900 16.050 310.950 ;
        RECT 13.950 308.850 16.050 309.900 ;
        RECT 19.950 308.850 22.950 310.950 ;
        RECT 12.450 305.100 14.250 305.400 ;
        RECT 12.450 304.800 20.850 305.100 ;
        RECT 3.150 304.200 20.850 304.800 ;
        RECT 3.150 303.600 14.250 304.200 ;
        RECT 3.150 291.750 4.950 303.600 ;
        RECT 17.250 302.700 19.050 303.300 ;
        RECT 11.550 301.500 19.050 302.700 ;
        RECT 19.950 302.100 20.850 304.200 ;
        RECT 22.050 304.200 22.950 308.850 ;
        RECT 32.250 305.400 34.050 307.200 ;
        RECT 28.950 304.200 33.150 305.400 ;
        RECT 22.050 303.300 28.050 304.200 ;
        RECT 28.950 303.300 31.050 304.200 ;
        RECT 35.250 303.600 36.450 313.050 ;
        RECT 64.950 311.850 67.050 313.950 ;
        RECT 65.100 310.050 66.900 311.850 ;
        RECT 67.950 308.850 70.050 310.950 ;
        RECT 68.100 307.050 69.900 308.850 ;
        RECT 71.700 306.150 72.600 314.400 ;
        RECT 75.000 312.150 76.050 317.400 ;
        RECT 73.950 310.050 76.050 312.150 ;
        RECT 112.650 310.950 113.850 317.400 ;
        RECT 118.650 316.500 119.850 320.400 ;
        RECT 114.750 315.600 119.850 316.500 ;
        RECT 155.850 316.200 157.650 323.250 ;
        RECT 160.350 317.400 162.150 323.250 ;
        RECT 194.550 320.400 196.350 323.250 ;
        RECT 197.550 320.400 199.350 323.250 ;
        RECT 114.750 314.700 117.000 315.600 ;
        RECT 155.850 315.300 159.450 316.200 ;
        RECT 70.950 306.000 72.750 306.150 ;
        RECT 27.150 302.400 28.050 303.300 ;
        RECT 24.450 302.100 26.250 302.400 ;
        RECT 11.550 300.600 12.750 301.500 ;
        RECT 19.950 301.200 26.250 302.100 ;
        RECT 24.450 300.600 26.250 301.200 ;
        RECT 27.150 300.600 29.850 302.400 ;
        RECT 7.950 298.500 12.750 300.600 ;
        RECT 15.150 298.500 22.050 300.300 ;
        RECT 11.550 297.600 12.750 298.500 ;
        RECT 6.150 291.750 7.950 297.600 ;
        RECT 11.250 291.750 13.050 297.600 ;
        RECT 16.050 291.750 17.850 297.600 ;
        RECT 19.050 291.750 20.850 298.500 ;
        RECT 27.150 297.600 31.050 299.700 ;
        RECT 22.950 291.750 24.750 297.600 ;
        RECT 27.150 291.750 28.950 297.600 ;
        RECT 31.650 291.750 33.450 294.600 ;
        RECT 34.650 291.750 36.450 303.600 ;
        RECT 65.550 304.800 72.750 306.000 ;
        RECT 65.550 303.600 66.750 304.800 ;
        RECT 70.950 304.350 72.750 304.800 ;
        RECT 65.550 291.750 67.350 303.600 ;
        RECT 74.100 303.450 75.450 310.050 ;
        RECT 112.650 308.850 115.050 310.950 ;
        RECT 112.650 303.600 113.850 308.850 ;
        RECT 115.950 306.300 117.000 314.700 ;
        RECT 118.950 308.850 121.050 310.950 ;
        RECT 155.100 309.150 156.900 310.950 ;
        RECT 119.100 307.050 120.900 308.850 ;
        RECT 154.950 307.050 157.050 309.150 ;
        RECT 158.250 307.950 159.450 315.300 ;
        RECT 193.950 311.850 196.050 313.950 ;
        RECT 197.400 312.150 198.600 320.400 ;
        RECT 233.850 317.400 235.650 323.250 ;
        RECT 238.350 316.200 240.150 323.250 ;
        RECT 272.550 320.400 274.350 323.250 ;
        RECT 275.550 320.400 277.350 323.250 ;
        RECT 278.550 320.400 280.350 323.250 ;
        RECT 236.550 315.300 240.150 316.200 ;
        RECT 276.450 316.200 277.350 320.400 ;
        RECT 281.550 317.400 283.350 323.250 ;
        RECT 319.650 317.400 321.450 323.250 ;
        RECT 276.450 315.300 279.750 316.200 ;
        RECT 161.100 309.150 162.900 310.950 ;
        RECT 194.100 310.050 195.900 311.850 ;
        RECT 196.950 310.050 199.050 312.150 ;
        RECT 114.750 305.400 117.000 306.300 ;
        RECT 157.950 305.850 160.050 307.950 ;
        RECT 160.950 307.050 163.050 309.150 ;
        RECT 114.750 304.500 120.450 305.400 ;
        RECT 70.050 291.750 71.850 303.450 ;
        RECT 73.050 302.100 75.450 303.450 ;
        RECT 73.050 291.750 74.850 302.100 ;
        RECT 112.350 291.750 114.150 303.600 ;
        RECT 115.350 291.750 117.150 303.600 ;
        RECT 119.250 297.600 120.450 304.500 ;
        RECT 158.250 297.600 159.450 305.850 ;
        RECT 197.400 297.600 198.600 310.050 ;
        RECT 233.100 309.150 234.900 310.950 ;
        RECT 232.950 307.050 235.050 309.150 ;
        RECT 236.550 307.950 237.750 315.300 ;
        RECT 277.950 314.400 279.750 315.300 ;
        RECT 271.950 311.850 274.050 313.950 ;
        RECT 239.100 309.150 240.900 310.950 ;
        RECT 272.100 310.050 273.900 311.850 ;
        RECT 235.950 305.850 238.050 307.950 ;
        RECT 238.950 307.050 241.050 309.150 ;
        RECT 274.950 308.850 277.050 310.950 ;
        RECT 275.100 307.050 276.900 308.850 ;
        RECT 278.700 306.150 279.600 314.400 ;
        RECT 282.000 312.150 283.050 317.400 ;
        RECT 320.250 315.300 321.450 317.400 ;
        RECT 322.650 318.300 324.450 323.250 ;
        RECT 325.650 319.200 327.450 323.250 ;
        RECT 328.650 318.300 330.450 323.250 ;
        RECT 359.550 320.400 361.350 323.250 ;
        RECT 362.550 320.400 364.350 323.250 ;
        RECT 322.650 316.950 330.450 318.300 ;
        RECT 320.250 314.250 324.000 315.300 ;
        RECT 280.950 310.050 283.050 312.150 ;
        RECT 322.950 310.950 324.150 314.250 ;
        RECT 326.100 312.150 327.900 313.950 ;
        RECT 277.950 306.000 279.750 306.150 ;
        RECT 236.550 297.600 237.750 305.850 ;
        RECT 272.550 304.800 279.750 306.000 ;
        RECT 272.550 303.600 273.750 304.800 ;
        RECT 277.950 304.350 279.750 304.800 ;
        RECT 118.650 291.750 120.450 297.600 ;
        RECT 154.650 291.750 156.450 297.600 ;
        RECT 157.650 291.750 159.450 297.600 ;
        RECT 160.650 291.750 162.450 297.600 ;
        RECT 194.550 291.750 196.350 297.600 ;
        RECT 197.550 291.750 199.350 297.600 ;
        RECT 233.550 291.750 235.350 297.600 ;
        RECT 236.550 291.750 238.350 297.600 ;
        RECT 239.550 291.750 241.350 297.600 ;
        RECT 272.550 291.750 274.350 303.600 ;
        RECT 281.100 303.450 282.450 310.050 ;
        RECT 322.950 308.850 325.050 310.950 ;
        RECT 325.950 310.050 328.050 312.150 ;
        RECT 358.950 311.850 361.050 313.950 ;
        RECT 362.400 312.150 363.600 320.400 ;
        RECT 397.650 317.400 399.450 323.250 ;
        RECT 398.250 315.300 399.450 317.400 ;
        RECT 400.650 318.300 402.450 323.250 ;
        RECT 403.650 319.200 405.450 323.250 ;
        RECT 406.650 318.300 408.450 323.250 ;
        RECT 440.550 320.400 442.350 323.250 ;
        RECT 443.550 320.400 445.350 323.250 ;
        RECT 400.650 316.950 408.450 318.300 ;
        RECT 398.250 314.250 402.000 315.300 ;
        RECT 328.950 308.850 331.050 310.950 ;
        RECT 359.100 310.050 360.900 311.850 ;
        RECT 361.950 310.050 364.050 312.150 ;
        RECT 400.950 310.950 402.150 314.250 ;
        RECT 404.100 312.150 405.900 313.950 ;
        RECT 319.950 305.850 322.050 307.950 ;
        RECT 320.250 304.050 322.050 305.850 ;
        RECT 323.850 303.600 325.050 308.850 ;
        RECT 329.100 307.050 330.900 308.850 ;
        RECT 277.050 291.750 278.850 303.450 ;
        RECT 280.050 302.100 282.450 303.450 ;
        RECT 280.050 291.750 281.850 302.100 ;
        RECT 320.400 291.750 322.200 297.600 ;
        RECT 323.700 291.750 325.500 303.600 ;
        RECT 327.900 291.750 329.700 303.600 ;
        RECT 362.400 297.600 363.600 310.050 ;
        RECT 400.950 308.850 403.050 310.950 ;
        RECT 403.950 310.050 406.050 312.150 ;
        RECT 439.950 311.850 442.050 313.950 ;
        RECT 443.400 312.150 444.600 320.400 ;
        RECT 479.550 318.300 481.350 323.250 ;
        RECT 482.550 319.200 484.350 323.250 ;
        RECT 485.550 318.300 487.350 323.250 ;
        RECT 479.550 316.950 487.350 318.300 ;
        RECT 488.550 317.400 490.350 323.250 ;
        RECT 524.850 317.400 526.650 323.250 ;
        RECT 488.550 315.300 489.750 317.400 ;
        RECT 529.350 316.200 531.150 323.250 ;
        RECT 568.650 320.400 570.450 323.250 ;
        RECT 571.650 320.400 573.450 323.250 ;
        RECT 607.650 320.400 609.450 323.250 ;
        RECT 610.650 320.400 612.450 323.250 ;
        RECT 486.000 314.250 489.750 315.300 ;
        RECT 527.550 315.300 531.150 316.200 ;
        RECT 482.100 312.150 483.900 313.950 ;
        RECT 406.950 308.850 409.050 310.950 ;
        RECT 440.100 310.050 441.900 311.850 ;
        RECT 442.950 310.050 445.050 312.150 ;
        RECT 397.950 305.850 400.050 307.950 ;
        RECT 398.250 304.050 400.050 305.850 ;
        RECT 401.850 303.600 403.050 308.850 ;
        RECT 407.100 307.050 408.900 308.850 ;
        RECT 427.950 306.450 430.050 307.050 ;
        RECT 439.950 306.450 442.050 307.050 ;
        RECT 427.950 305.550 442.050 306.450 ;
        RECT 427.950 304.950 430.050 305.550 ;
        RECT 439.950 304.950 442.050 305.550 ;
        RECT 359.550 291.750 361.350 297.600 ;
        RECT 362.550 291.750 364.350 297.600 ;
        RECT 398.400 291.750 400.200 297.600 ;
        RECT 401.700 291.750 403.500 303.600 ;
        RECT 405.900 291.750 407.700 303.600 ;
        RECT 443.400 297.600 444.600 310.050 ;
        RECT 478.950 308.850 481.050 310.950 ;
        RECT 481.950 310.050 484.050 312.150 ;
        RECT 485.850 310.950 487.050 314.250 ;
        RECT 484.950 308.850 487.050 310.950 ;
        RECT 524.100 309.150 525.900 310.950 ;
        RECT 479.100 307.050 480.900 308.850 ;
        RECT 484.950 303.600 486.150 308.850 ;
        RECT 487.950 305.850 490.050 307.950 ;
        RECT 523.950 307.050 526.050 309.150 ;
        RECT 527.550 307.950 528.750 315.300 ;
        RECT 569.400 312.150 570.600 320.400 ;
        RECT 530.100 309.150 531.900 310.950 ;
        RECT 568.950 310.050 571.050 312.150 ;
        RECT 571.950 311.850 574.050 313.950 ;
        RECT 608.400 312.150 609.600 320.400 ;
        RECT 643.650 317.400 645.450 323.250 ;
        RECT 644.250 315.300 645.450 317.400 ;
        RECT 646.650 318.300 648.450 323.250 ;
        RECT 649.650 319.200 651.450 323.250 ;
        RECT 652.650 318.300 654.450 323.250 ;
        RECT 646.650 316.950 654.450 318.300 ;
        RECT 657.150 317.400 658.950 323.250 ;
        RECT 660.150 320.400 661.950 323.250 ;
        RECT 664.950 321.300 666.750 323.250 ;
        RECT 663.000 320.400 666.750 321.300 ;
        RECT 669.450 320.400 671.250 323.250 ;
        RECT 672.750 320.400 674.550 323.250 ;
        RECT 676.650 320.400 678.450 323.250 ;
        RECT 680.850 320.400 682.650 323.250 ;
        RECT 685.350 320.400 687.150 323.250 ;
        RECT 663.000 319.500 664.050 320.400 ;
        RECT 661.950 317.400 664.050 319.500 ;
        RECT 672.750 318.600 673.800 320.400 ;
        RECT 644.250 314.250 648.000 315.300 ;
        RECT 572.100 310.050 573.900 311.850 ;
        RECT 607.950 310.050 610.050 312.150 ;
        RECT 610.950 311.850 613.050 313.950 ;
        RECT 611.100 310.050 612.900 311.850 ;
        RECT 646.950 310.950 648.150 314.250 ;
        RECT 650.100 312.150 651.900 313.950 ;
        RECT 526.950 305.850 529.050 307.950 ;
        RECT 529.950 307.050 532.050 309.150 ;
        RECT 487.950 304.050 489.750 305.850 ;
        RECT 440.550 291.750 442.350 297.600 ;
        RECT 443.550 291.750 445.350 297.600 ;
        RECT 480.300 291.750 482.100 303.600 ;
        RECT 484.500 291.750 486.300 303.600 ;
        RECT 527.550 297.600 528.750 305.850 ;
        RECT 569.400 297.600 570.600 310.050 ;
        RECT 608.400 297.600 609.600 310.050 ;
        RECT 646.950 308.850 649.050 310.950 ;
        RECT 649.950 310.050 652.050 312.150 ;
        RECT 652.950 308.850 655.050 310.950 ;
        RECT 643.950 305.850 646.050 307.950 ;
        RECT 644.250 304.050 646.050 305.850 ;
        RECT 647.850 303.600 649.050 308.850 ;
        RECT 653.100 307.050 654.900 308.850 ;
        RECT 657.150 304.800 658.050 317.400 ;
        RECT 665.550 316.800 667.350 318.600 ;
        RECT 668.850 317.550 673.800 318.600 ;
        RECT 681.300 319.500 682.350 320.400 ;
        RECT 681.300 318.300 685.050 319.500 ;
        RECT 668.850 316.800 670.650 317.550 ;
        RECT 665.850 315.900 666.900 316.800 ;
        RECT 676.050 316.200 677.850 318.000 ;
        RECT 682.950 317.400 685.050 318.300 ;
        RECT 688.650 317.400 690.450 323.250 ;
        RECT 676.050 315.900 676.950 316.200 ;
        RECT 665.850 315.000 676.950 315.900 ;
        RECT 689.250 315.150 690.450 317.400 ;
        RECT 722.850 316.200 724.650 323.250 ;
        RECT 727.350 317.400 729.150 323.250 ;
        RECT 722.850 315.300 726.450 316.200 ;
        RECT 665.850 313.800 666.900 315.000 ;
        RECT 660.000 312.600 666.900 313.800 ;
        RECT 660.000 311.850 660.900 312.600 ;
        RECT 665.100 312.000 666.900 312.600 ;
        RECT 659.100 310.050 660.900 311.850 ;
        RECT 662.100 310.950 663.900 311.700 ;
        RECT 676.050 310.950 676.950 315.000 ;
        RECT 685.950 313.050 690.450 315.150 ;
        RECT 684.150 311.250 688.050 313.050 ;
        RECT 685.950 310.950 688.050 311.250 ;
        RECT 662.100 309.900 670.050 310.950 ;
        RECT 667.950 308.850 670.050 309.900 ;
        RECT 673.950 308.850 676.950 310.950 ;
        RECT 666.450 305.100 668.250 305.400 ;
        RECT 666.450 304.800 674.850 305.100 ;
        RECT 657.150 304.200 674.850 304.800 ;
        RECT 657.150 303.600 668.250 304.200 ;
        RECT 487.800 291.750 489.600 297.600 ;
        RECT 524.550 291.750 526.350 297.600 ;
        RECT 527.550 291.750 529.350 297.600 ;
        RECT 530.550 291.750 532.350 297.600 ;
        RECT 568.650 291.750 570.450 297.600 ;
        RECT 571.650 291.750 573.450 297.600 ;
        RECT 607.650 291.750 609.450 297.600 ;
        RECT 610.650 291.750 612.450 297.600 ;
        RECT 644.400 291.750 646.200 297.600 ;
        RECT 647.700 291.750 649.500 303.600 ;
        RECT 651.900 291.750 653.700 303.600 ;
        RECT 657.150 291.750 658.950 303.600 ;
        RECT 671.250 302.700 673.050 303.300 ;
        RECT 665.550 301.500 673.050 302.700 ;
        RECT 673.950 302.100 674.850 304.200 ;
        RECT 676.050 304.200 676.950 308.850 ;
        RECT 686.250 305.400 688.050 307.200 ;
        RECT 682.950 304.200 687.150 305.400 ;
        RECT 676.050 303.300 682.050 304.200 ;
        RECT 682.950 303.300 685.050 304.200 ;
        RECT 689.250 303.600 690.450 313.050 ;
        RECT 722.100 309.150 723.900 310.950 ;
        RECT 721.950 307.050 724.050 309.150 ;
        RECT 725.250 307.950 726.450 315.300 ;
        RECT 728.100 309.150 729.900 310.950 ;
        RECT 724.950 305.850 727.050 307.950 ;
        RECT 727.950 307.050 730.050 309.150 ;
        RECT 681.150 302.400 682.050 303.300 ;
        RECT 678.450 302.100 680.250 302.400 ;
        RECT 665.550 300.600 666.750 301.500 ;
        RECT 673.950 301.200 680.250 302.100 ;
        RECT 678.450 300.600 680.250 301.200 ;
        RECT 681.150 300.600 683.850 302.400 ;
        RECT 661.950 298.500 666.750 300.600 ;
        RECT 669.150 298.500 676.050 300.300 ;
        RECT 665.550 297.600 666.750 298.500 ;
        RECT 660.150 291.750 661.950 297.600 ;
        RECT 665.250 291.750 667.050 297.600 ;
        RECT 670.050 291.750 671.850 297.600 ;
        RECT 673.050 291.750 674.850 298.500 ;
        RECT 681.150 297.600 685.050 299.700 ;
        RECT 676.950 291.750 678.750 297.600 ;
        RECT 681.150 291.750 682.950 297.600 ;
        RECT 685.650 291.750 687.450 294.600 ;
        RECT 688.650 291.750 690.450 303.600 ;
        RECT 725.250 297.600 726.450 305.850 ;
        RECT 721.650 291.750 723.450 297.600 ;
        RECT 724.650 291.750 726.450 297.600 ;
        RECT 727.650 291.750 729.450 297.600 ;
        RECT 32.400 281.400 34.200 287.250 ;
        RECT 35.700 275.400 37.500 287.250 ;
        RECT 39.900 275.400 41.700 287.250 ;
        RECT 75.300 275.400 77.100 287.250 ;
        RECT 79.500 275.400 81.300 287.250 ;
        RECT 82.800 281.400 84.600 287.250 ;
        RECT 90.150 275.400 91.950 287.250 ;
        RECT 93.150 281.400 94.950 287.250 ;
        RECT 98.250 281.400 100.050 287.250 ;
        RECT 103.050 281.400 104.850 287.250 ;
        RECT 98.550 280.500 99.750 281.400 ;
        RECT 106.050 280.500 107.850 287.250 ;
        RECT 109.950 281.400 111.750 287.250 ;
        RECT 114.150 281.400 115.950 287.250 ;
        RECT 118.650 284.400 120.450 287.250 ;
        RECT 94.950 278.400 99.750 280.500 ;
        RECT 102.150 278.700 109.050 280.500 ;
        RECT 114.150 279.300 118.050 281.400 ;
        RECT 98.550 277.500 99.750 278.400 ;
        RECT 111.450 277.800 113.250 278.400 ;
        RECT 98.550 276.300 106.050 277.500 ;
        RECT 104.250 275.700 106.050 276.300 ;
        RECT 106.950 276.900 113.250 277.800 ;
        RECT 32.250 273.150 34.050 274.950 ;
        RECT 31.950 271.050 34.050 273.150 ;
        RECT 35.850 270.150 37.050 275.400 ;
        RECT 41.100 270.150 42.900 271.950 ;
        RECT 74.100 270.150 75.900 271.950 ;
        RECT 79.950 270.150 81.150 275.400 ;
        RECT 82.950 273.150 84.750 274.950 ;
        RECT 90.150 274.800 101.250 275.400 ;
        RECT 106.950 274.800 107.850 276.900 ;
        RECT 111.450 276.600 113.250 276.900 ;
        RECT 114.150 276.600 116.850 278.400 ;
        RECT 114.150 275.700 115.050 276.600 ;
        RECT 90.150 274.200 107.850 274.800 ;
        RECT 82.950 271.050 85.050 273.150 ;
        RECT 34.950 268.050 37.050 270.150 ;
        RECT 34.950 264.750 36.150 268.050 ;
        RECT 37.950 266.850 40.050 268.950 ;
        RECT 40.950 268.050 43.050 270.150 ;
        RECT 73.950 268.050 76.050 270.150 ;
        RECT 76.950 266.850 79.050 268.950 ;
        RECT 79.950 268.050 82.050 270.150 ;
        RECT 38.100 265.050 39.900 266.850 ;
        RECT 77.100 265.050 78.900 266.850 ;
        RECT 80.850 264.750 82.050 268.050 ;
        RECT 32.250 263.700 36.000 264.750 ;
        RECT 81.000 263.700 84.750 264.750 ;
        RECT 32.250 261.600 33.450 263.700 ;
        RECT 31.650 255.750 33.450 261.600 ;
        RECT 34.650 260.700 42.450 262.050 ;
        RECT 34.650 255.750 36.450 260.700 ;
        RECT 37.650 255.750 39.450 259.800 ;
        RECT 40.650 255.750 42.450 260.700 ;
        RECT 74.550 260.700 82.350 262.050 ;
        RECT 74.550 255.750 76.350 260.700 ;
        RECT 77.550 255.750 79.350 259.800 ;
        RECT 80.550 255.750 82.350 260.700 ;
        RECT 83.550 261.600 84.750 263.700 ;
        RECT 90.150 261.600 91.050 274.200 ;
        RECT 99.450 273.900 107.850 274.200 ;
        RECT 109.050 274.800 115.050 275.700 ;
        RECT 115.950 274.800 118.050 275.700 ;
        RECT 121.650 275.400 123.450 287.250 ;
        RECT 155.550 281.400 157.350 287.250 ;
        RECT 158.550 281.400 160.350 287.250 ;
        RECT 191.550 281.400 193.350 287.250 ;
        RECT 194.550 281.400 196.350 287.250 ;
        RECT 197.550 282.000 199.350 287.250 ;
        RECT 99.450 273.600 101.250 273.900 ;
        RECT 109.050 270.150 109.950 274.800 ;
        RECT 115.950 273.600 120.150 274.800 ;
        RECT 119.250 271.800 121.050 273.600 ;
        RECT 100.950 269.100 103.050 270.150 ;
        RECT 92.100 267.150 93.900 268.950 ;
        RECT 95.100 268.050 103.050 269.100 ;
        RECT 106.950 268.050 109.950 270.150 ;
        RECT 95.100 267.300 96.900 268.050 ;
        RECT 93.000 266.400 93.900 267.150 ;
        RECT 98.100 266.400 99.900 267.000 ;
        RECT 93.000 265.200 99.900 266.400 ;
        RECT 98.850 264.000 99.900 265.200 ;
        RECT 109.050 264.000 109.950 268.050 ;
        RECT 118.950 267.750 121.050 268.050 ;
        RECT 117.150 265.950 121.050 267.750 ;
        RECT 122.250 265.950 123.450 275.400 ;
        RECT 158.400 268.950 159.600 281.400 ;
        RECT 194.700 281.100 196.350 281.400 ;
        RECT 200.550 281.400 202.350 287.250 ;
        RECT 236.550 281.400 238.350 287.250 ;
        RECT 239.550 281.400 241.350 287.250 ;
        RECT 242.550 281.400 244.350 287.250 ;
        RECT 278.550 281.400 280.350 287.250 ;
        RECT 281.550 281.400 283.350 287.250 ;
        RECT 284.550 282.000 286.350 287.250 ;
        RECT 200.550 281.100 201.750 281.400 ;
        RECT 194.700 280.200 201.750 281.100 ;
        RECT 194.100 276.150 195.900 277.950 ;
        RECT 191.100 273.150 192.900 274.950 ;
        RECT 193.950 274.050 196.050 276.150 ;
        RECT 197.250 273.150 199.050 274.950 ;
        RECT 190.950 271.050 193.050 273.150 ;
        RECT 196.950 271.050 199.050 273.150 ;
        RECT 200.700 271.950 201.750 280.200 ;
        RECT 211.950 276.450 214.050 277.050 ;
        RECT 235.950 276.450 238.050 277.050 ;
        RECT 211.950 275.550 238.050 276.450 ;
        RECT 211.950 274.950 214.050 275.550 ;
        RECT 235.950 274.950 238.050 275.550 ;
        RECT 239.550 273.150 240.750 281.400 ;
        RECT 281.700 281.100 283.350 281.400 ;
        RECT 287.550 281.400 289.350 287.250 ;
        RECT 323.550 281.400 325.350 287.250 ;
        RECT 326.550 281.400 328.350 287.250 ;
        RECT 329.550 281.400 331.350 287.250 ;
        RECT 287.550 281.100 288.750 281.400 ;
        RECT 281.700 280.200 288.750 281.100 ;
        RECT 281.100 276.150 282.900 277.950 ;
        RECT 278.100 273.150 279.900 274.950 ;
        RECT 280.950 274.050 283.050 276.150 ;
        RECT 284.250 273.150 286.050 274.950 ;
        RECT 199.950 269.850 202.050 271.950 ;
        RECT 235.950 269.850 238.050 271.950 ;
        RECT 238.950 271.050 241.050 273.150 ;
        RECT 155.100 267.150 156.900 268.950 ;
        RECT 98.850 263.100 109.950 264.000 ;
        RECT 118.950 263.850 123.450 265.950 ;
        RECT 154.950 265.050 157.050 267.150 ;
        RECT 157.950 266.850 160.050 268.950 ;
        RECT 98.850 262.200 99.900 263.100 ;
        RECT 109.050 262.800 109.950 263.100 ;
        RECT 83.550 255.750 85.350 261.600 ;
        RECT 90.150 255.750 91.950 261.600 ;
        RECT 94.950 259.500 97.050 261.600 ;
        RECT 98.550 260.400 100.350 262.200 ;
        RECT 101.850 261.450 103.650 262.200 ;
        RECT 101.850 260.400 106.800 261.450 ;
        RECT 109.050 261.000 110.850 262.800 ;
        RECT 122.250 261.600 123.450 263.850 ;
        RECT 115.950 260.700 118.050 261.600 ;
        RECT 96.000 258.600 97.050 259.500 ;
        RECT 105.750 258.600 106.800 260.400 ;
        RECT 114.300 259.500 118.050 260.700 ;
        RECT 114.300 258.600 115.350 259.500 ;
        RECT 93.150 255.750 94.950 258.600 ;
        RECT 96.000 257.700 99.750 258.600 ;
        RECT 97.950 255.750 99.750 257.700 ;
        RECT 102.450 255.750 104.250 258.600 ;
        RECT 105.750 255.750 107.550 258.600 ;
        RECT 109.650 255.750 111.450 258.600 ;
        RECT 113.850 255.750 115.650 258.600 ;
        RECT 118.350 255.750 120.150 258.600 ;
        RECT 121.650 255.750 123.450 261.600 ;
        RECT 158.400 258.600 159.600 266.850 ;
        RECT 200.400 265.650 201.600 269.850 ;
        RECT 236.100 268.050 237.900 269.850 ;
        RECT 155.550 255.750 157.350 258.600 ;
        RECT 158.550 255.750 160.350 258.600 ;
        RECT 191.700 255.750 193.500 264.600 ;
        RECT 197.100 264.000 201.600 265.650 ;
        RECT 197.100 255.750 198.900 264.000 ;
        RECT 239.550 263.700 240.750 271.050 ;
        RECT 241.950 269.850 244.050 271.950 ;
        RECT 277.950 271.050 280.050 273.150 ;
        RECT 283.950 271.050 286.050 273.150 ;
        RECT 287.700 271.950 288.750 280.200 ;
        RECT 326.550 273.150 327.750 281.400 ;
        RECT 362.550 275.400 364.350 287.250 ;
        RECT 366.750 275.400 368.550 287.250 ;
        RECT 404.550 281.400 406.350 287.250 ;
        RECT 407.550 281.400 409.350 287.250 ;
        RECT 445.650 281.400 447.450 287.250 ;
        RECT 448.650 281.400 450.450 287.250 ;
        RECT 451.650 281.400 453.450 287.250 ;
        RECT 366.000 274.350 368.550 275.400 ;
        RECT 286.950 269.850 289.050 271.950 ;
        RECT 322.950 269.850 325.050 271.950 ;
        RECT 325.950 271.050 328.050 273.150 ;
        RECT 242.100 268.050 243.900 269.850 ;
        RECT 287.400 265.650 288.600 269.850 ;
        RECT 323.100 268.050 324.900 269.850 ;
        RECT 239.550 262.800 243.150 263.700 ;
        RECT 236.850 255.750 238.650 261.600 ;
        RECT 241.350 255.750 243.150 262.800 ;
        RECT 278.700 255.750 280.500 264.600 ;
        RECT 284.100 264.000 288.600 265.650 ;
        RECT 284.100 255.750 285.900 264.000 ;
        RECT 326.550 263.700 327.750 271.050 ;
        RECT 328.950 269.850 331.050 271.950 ;
        RECT 362.100 270.150 363.900 271.950 ;
        RECT 329.100 268.050 330.900 269.850 ;
        RECT 361.950 268.050 364.050 270.150 ;
        RECT 366.000 267.150 367.050 274.350 ;
        RECT 368.100 270.150 369.900 271.950 ;
        RECT 367.950 268.050 370.050 270.150 ;
        RECT 407.400 268.950 408.600 281.400 ;
        RECT 449.250 273.150 450.450 281.400 ;
        RECT 482.550 275.400 484.350 287.250 ;
        RECT 487.050 275.550 488.850 287.250 ;
        RECT 490.050 276.900 491.850 287.250 ;
        RECT 529.650 281.400 531.450 287.250 ;
        RECT 532.650 281.400 534.450 287.250 ;
        RECT 535.650 281.400 537.450 287.250 ;
        RECT 572.400 281.400 574.200 287.250 ;
        RECT 490.050 275.550 492.450 276.900 ;
        RECT 482.550 274.200 483.750 275.400 ;
        RECT 487.950 274.200 489.750 274.650 ;
        RECT 445.950 269.850 448.050 271.950 ;
        RECT 448.950 271.050 451.050 273.150 ;
        RECT 482.550 273.000 489.750 274.200 ;
        RECT 487.950 272.850 489.750 273.000 ;
        RECT 404.100 267.150 405.900 268.950 ;
        RECT 364.950 265.050 367.050 267.150 ;
        RECT 403.950 265.050 406.050 267.150 ;
        RECT 406.950 266.850 409.050 268.950 ;
        RECT 446.100 268.050 447.900 269.850 ;
        RECT 326.550 262.800 330.150 263.700 ;
        RECT 323.850 255.750 325.650 261.600 ;
        RECT 328.350 255.750 330.150 262.800 ;
        RECT 366.000 258.600 367.050 265.050 ;
        RECT 407.400 258.600 408.600 266.850 ;
        RECT 449.250 263.700 450.450 271.050 ;
        RECT 451.950 269.850 454.050 271.950 ;
        RECT 485.100 270.150 486.900 271.950 ;
        RECT 452.100 268.050 453.900 269.850 ;
        RECT 482.100 267.150 483.900 268.950 ;
        RECT 484.950 268.050 487.050 270.150 ;
        RECT 481.950 265.050 484.050 267.150 ;
        RECT 488.700 264.600 489.600 272.850 ;
        RECT 491.100 268.950 492.450 275.550 ;
        RECT 533.250 273.150 534.450 281.400 ;
        RECT 575.700 275.400 577.500 287.250 ;
        RECT 579.900 275.400 581.700 287.250 ;
        RECT 585.150 275.400 586.950 287.250 ;
        RECT 588.150 281.400 589.950 287.250 ;
        RECT 593.250 281.400 595.050 287.250 ;
        RECT 598.050 281.400 599.850 287.250 ;
        RECT 593.550 280.500 594.750 281.400 ;
        RECT 601.050 280.500 602.850 287.250 ;
        RECT 604.950 281.400 606.750 287.250 ;
        RECT 609.150 281.400 610.950 287.250 ;
        RECT 613.650 284.400 615.450 287.250 ;
        RECT 589.950 278.400 594.750 280.500 ;
        RECT 597.150 278.700 604.050 280.500 ;
        RECT 609.150 279.300 613.050 281.400 ;
        RECT 593.550 277.500 594.750 278.400 ;
        RECT 606.450 277.800 608.250 278.400 ;
        RECT 593.550 276.300 601.050 277.500 ;
        RECT 599.250 275.700 601.050 276.300 ;
        RECT 601.950 276.900 608.250 277.800 ;
        RECT 572.250 273.150 574.050 274.950 ;
        RECT 529.950 269.850 532.050 271.950 ;
        RECT 532.950 271.050 535.050 273.150 ;
        RECT 490.950 266.850 493.050 268.950 ;
        RECT 530.100 268.050 531.900 269.850 ;
        RECT 487.950 263.700 489.750 264.600 ;
        RECT 446.850 262.800 450.450 263.700 ;
        RECT 486.450 262.800 489.750 263.700 ;
        RECT 362.550 255.750 364.350 258.600 ;
        RECT 365.550 255.750 367.350 258.600 ;
        RECT 368.550 255.750 370.350 258.600 ;
        RECT 404.550 255.750 406.350 258.600 ;
        RECT 407.550 255.750 409.350 258.600 ;
        RECT 446.850 255.750 448.650 262.800 ;
        RECT 451.350 255.750 453.150 261.600 ;
        RECT 486.450 258.600 487.350 262.800 ;
        RECT 492.000 261.600 493.050 266.850 ;
        RECT 533.250 263.700 534.450 271.050 ;
        RECT 535.950 269.850 538.050 271.950 ;
        RECT 571.950 271.050 574.050 273.150 ;
        RECT 575.850 270.150 577.050 275.400 ;
        RECT 585.150 274.800 596.250 275.400 ;
        RECT 601.950 274.800 602.850 276.900 ;
        RECT 606.450 276.600 608.250 276.900 ;
        RECT 609.150 276.600 611.850 278.400 ;
        RECT 609.150 275.700 610.050 276.600 ;
        RECT 585.150 274.200 602.850 274.800 ;
        RECT 581.100 270.150 582.900 271.950 ;
        RECT 536.100 268.050 537.900 269.850 ;
        RECT 574.950 268.050 577.050 270.150 ;
        RECT 574.950 264.750 576.150 268.050 ;
        RECT 577.950 266.850 580.050 268.950 ;
        RECT 580.950 268.050 583.050 270.150 ;
        RECT 578.100 265.050 579.900 266.850 ;
        RECT 530.850 262.800 534.450 263.700 ;
        RECT 572.250 263.700 576.000 264.750 ;
        RECT 482.550 255.750 484.350 258.600 ;
        RECT 485.550 255.750 487.350 258.600 ;
        RECT 488.550 255.750 490.350 258.600 ;
        RECT 491.550 255.750 493.350 261.600 ;
        RECT 530.850 255.750 532.650 262.800 ;
        RECT 572.250 261.600 573.450 263.700 ;
        RECT 535.350 255.750 537.150 261.600 ;
        RECT 571.650 255.750 573.450 261.600 ;
        RECT 574.650 260.700 582.450 262.050 ;
        RECT 574.650 255.750 576.450 260.700 ;
        RECT 577.650 255.750 579.450 259.800 ;
        RECT 580.650 255.750 582.450 260.700 ;
        RECT 585.150 261.600 586.050 274.200 ;
        RECT 594.450 273.900 602.850 274.200 ;
        RECT 604.050 274.800 610.050 275.700 ;
        RECT 610.950 274.800 613.050 275.700 ;
        RECT 616.650 275.400 618.450 287.250 ;
        RECT 651.300 275.400 653.100 287.250 ;
        RECT 655.500 275.400 657.300 287.250 ;
        RECT 658.800 281.400 660.600 287.250 ;
        RECT 697.650 281.400 699.450 287.250 ;
        RECT 700.650 281.400 702.450 287.250 ;
        RECT 703.650 281.400 705.450 287.250 ;
        RECT 594.450 273.600 596.250 273.900 ;
        RECT 604.050 270.150 604.950 274.800 ;
        RECT 610.950 273.600 615.150 274.800 ;
        RECT 614.250 271.800 616.050 273.600 ;
        RECT 595.950 269.100 598.050 270.150 ;
        RECT 587.100 267.150 588.900 268.950 ;
        RECT 590.100 268.050 598.050 269.100 ;
        RECT 601.950 268.050 604.950 270.150 ;
        RECT 590.100 267.300 591.900 268.050 ;
        RECT 588.000 266.400 588.900 267.150 ;
        RECT 593.100 266.400 594.900 267.000 ;
        RECT 588.000 265.200 594.900 266.400 ;
        RECT 593.850 264.000 594.900 265.200 ;
        RECT 604.050 264.000 604.950 268.050 ;
        RECT 613.950 267.750 616.050 268.050 ;
        RECT 612.150 265.950 616.050 267.750 ;
        RECT 617.250 265.950 618.450 275.400 ;
        RECT 650.100 270.150 651.900 271.950 ;
        RECT 655.950 270.150 657.150 275.400 ;
        RECT 658.950 273.150 660.750 274.950 ;
        RECT 701.250 273.150 702.450 281.400 ;
        RECT 708.150 275.400 709.950 287.250 ;
        RECT 711.150 281.400 712.950 287.250 ;
        RECT 716.250 281.400 718.050 287.250 ;
        RECT 721.050 281.400 722.850 287.250 ;
        RECT 716.550 280.500 717.750 281.400 ;
        RECT 724.050 280.500 725.850 287.250 ;
        RECT 727.950 281.400 729.750 287.250 ;
        RECT 732.150 281.400 733.950 287.250 ;
        RECT 736.650 284.400 738.450 287.250 ;
        RECT 712.950 278.400 717.750 280.500 ;
        RECT 720.150 278.700 727.050 280.500 ;
        RECT 732.150 279.300 736.050 281.400 ;
        RECT 716.550 277.500 717.750 278.400 ;
        RECT 729.450 277.800 731.250 278.400 ;
        RECT 716.550 276.300 724.050 277.500 ;
        RECT 722.250 275.700 724.050 276.300 ;
        RECT 724.950 276.900 731.250 277.800 ;
        RECT 708.150 274.800 719.250 275.400 ;
        RECT 724.950 274.800 725.850 276.900 ;
        RECT 729.450 276.600 731.250 276.900 ;
        RECT 732.150 276.600 734.850 278.400 ;
        RECT 732.150 275.700 733.050 276.600 ;
        RECT 708.150 274.200 725.850 274.800 ;
        RECT 658.950 271.050 661.050 273.150 ;
        RECT 649.950 268.050 652.050 270.150 ;
        RECT 652.950 266.850 655.050 268.950 ;
        RECT 655.950 268.050 658.050 270.150 ;
        RECT 697.950 269.850 700.050 271.950 ;
        RECT 700.950 271.050 703.050 273.150 ;
        RECT 698.100 268.050 699.900 269.850 ;
        RECT 593.850 263.100 604.950 264.000 ;
        RECT 613.950 263.850 618.450 265.950 ;
        RECT 653.100 265.050 654.900 266.850 ;
        RECT 656.850 264.750 658.050 268.050 ;
        RECT 593.850 262.200 594.900 263.100 ;
        RECT 604.050 262.800 604.950 263.100 ;
        RECT 585.150 255.750 586.950 261.600 ;
        RECT 589.950 259.500 592.050 261.600 ;
        RECT 593.550 260.400 595.350 262.200 ;
        RECT 596.850 261.450 598.650 262.200 ;
        RECT 596.850 260.400 601.800 261.450 ;
        RECT 604.050 261.000 605.850 262.800 ;
        RECT 617.250 261.600 618.450 263.850 ;
        RECT 657.000 263.700 660.750 264.750 ;
        RECT 701.250 263.700 702.450 271.050 ;
        RECT 703.950 269.850 706.050 271.950 ;
        RECT 704.100 268.050 705.900 269.850 ;
        RECT 610.950 260.700 613.050 261.600 ;
        RECT 591.000 258.600 592.050 259.500 ;
        RECT 600.750 258.600 601.800 260.400 ;
        RECT 609.300 259.500 613.050 260.700 ;
        RECT 609.300 258.600 610.350 259.500 ;
        RECT 588.150 255.750 589.950 258.600 ;
        RECT 591.000 257.700 594.750 258.600 ;
        RECT 592.950 255.750 594.750 257.700 ;
        RECT 597.450 255.750 599.250 258.600 ;
        RECT 600.750 255.750 602.550 258.600 ;
        RECT 604.650 255.750 606.450 258.600 ;
        RECT 608.850 255.750 610.650 258.600 ;
        RECT 613.350 255.750 615.150 258.600 ;
        RECT 616.650 255.750 618.450 261.600 ;
        RECT 650.550 260.700 658.350 262.050 ;
        RECT 650.550 255.750 652.350 260.700 ;
        RECT 653.550 255.750 655.350 259.800 ;
        RECT 656.550 255.750 658.350 260.700 ;
        RECT 659.550 261.600 660.750 263.700 ;
        RECT 698.850 262.800 702.450 263.700 ;
        RECT 659.550 255.750 661.350 261.600 ;
        RECT 698.850 255.750 700.650 262.800 ;
        RECT 708.150 261.600 709.050 274.200 ;
        RECT 717.450 273.900 725.850 274.200 ;
        RECT 727.050 274.800 733.050 275.700 ;
        RECT 733.950 274.800 736.050 275.700 ;
        RECT 739.650 275.400 741.450 287.250 ;
        RECT 717.450 273.600 719.250 273.900 ;
        RECT 727.050 270.150 727.950 274.800 ;
        RECT 733.950 273.600 738.150 274.800 ;
        RECT 737.250 271.800 739.050 273.600 ;
        RECT 718.950 269.100 721.050 270.150 ;
        RECT 710.100 267.150 711.900 268.950 ;
        RECT 713.100 268.050 721.050 269.100 ;
        RECT 724.950 268.050 727.950 270.150 ;
        RECT 713.100 267.300 714.900 268.050 ;
        RECT 711.000 266.400 711.900 267.150 ;
        RECT 716.100 266.400 717.900 267.000 ;
        RECT 711.000 265.200 717.900 266.400 ;
        RECT 716.850 264.000 717.900 265.200 ;
        RECT 727.050 264.000 727.950 268.050 ;
        RECT 736.950 267.750 739.050 268.050 ;
        RECT 735.150 265.950 739.050 267.750 ;
        RECT 740.250 265.950 741.450 275.400 ;
        RECT 716.850 263.100 727.950 264.000 ;
        RECT 736.950 263.850 741.450 265.950 ;
        RECT 716.850 262.200 717.900 263.100 ;
        RECT 727.050 262.800 727.950 263.100 ;
        RECT 703.350 255.750 705.150 261.600 ;
        RECT 708.150 255.750 709.950 261.600 ;
        RECT 712.950 259.500 715.050 261.600 ;
        RECT 716.550 260.400 718.350 262.200 ;
        RECT 719.850 261.450 721.650 262.200 ;
        RECT 719.850 260.400 724.800 261.450 ;
        RECT 727.050 261.000 728.850 262.800 ;
        RECT 740.250 261.600 741.450 263.850 ;
        RECT 733.950 260.700 736.050 261.600 ;
        RECT 714.000 258.600 715.050 259.500 ;
        RECT 723.750 258.600 724.800 260.400 ;
        RECT 732.300 259.500 736.050 260.700 ;
        RECT 732.300 258.600 733.350 259.500 ;
        RECT 711.150 255.750 712.950 258.600 ;
        RECT 714.000 257.700 717.750 258.600 ;
        RECT 715.950 255.750 717.750 257.700 ;
        RECT 720.450 255.750 722.250 258.600 ;
        RECT 723.750 255.750 725.550 258.600 ;
        RECT 727.650 255.750 729.450 258.600 ;
        RECT 731.850 255.750 733.650 258.600 ;
        RECT 736.350 255.750 738.150 258.600 ;
        RECT 739.650 255.750 741.450 261.600 ;
        RECT 34.650 245.400 36.450 251.250 ;
        RECT 35.250 243.300 36.450 245.400 ;
        RECT 37.650 246.300 39.450 251.250 ;
        RECT 40.650 247.200 42.450 251.250 ;
        RECT 43.650 246.300 45.450 251.250 ;
        RECT 37.650 244.950 45.450 246.300 ;
        RECT 79.650 245.400 81.450 251.250 ;
        RECT 80.250 243.300 81.450 245.400 ;
        RECT 82.650 246.300 84.450 251.250 ;
        RECT 85.650 247.200 87.450 251.250 ;
        RECT 88.650 246.300 90.450 251.250 ;
        RECT 82.650 244.950 90.450 246.300 ;
        RECT 125.850 244.200 127.650 251.250 ;
        RECT 130.350 245.400 132.150 251.250 ;
        RECT 163.650 248.400 165.450 251.250 ;
        RECT 166.650 248.400 168.450 251.250 ;
        RECT 125.850 243.300 129.450 244.200 ;
        RECT 35.250 242.250 39.000 243.300 ;
        RECT 80.250 242.250 84.000 243.300 ;
        RECT 37.950 238.950 39.150 242.250 ;
        RECT 41.100 240.150 42.900 241.950 ;
        RECT 37.950 236.850 40.050 238.950 ;
        RECT 40.950 238.050 43.050 240.150 ;
        RECT 82.950 238.950 84.150 242.250 ;
        RECT 86.100 240.150 87.900 241.950 ;
        RECT 43.950 236.850 46.050 238.950 ;
        RECT 82.950 236.850 85.050 238.950 ;
        RECT 85.950 238.050 88.050 240.150 ;
        RECT 88.950 236.850 91.050 238.950 ;
        RECT 125.100 237.150 126.900 238.950 ;
        RECT 34.950 233.850 37.050 235.950 ;
        RECT 35.250 232.050 37.050 233.850 ;
        RECT 38.850 231.600 40.050 236.850 ;
        RECT 44.100 235.050 45.900 236.850 ;
        RECT 79.950 233.850 82.050 235.950 ;
        RECT 80.250 232.050 82.050 233.850 ;
        RECT 83.850 231.600 85.050 236.850 ;
        RECT 89.100 235.050 90.900 236.850 ;
        RECT 124.950 235.050 127.050 237.150 ;
        RECT 128.250 235.950 129.450 243.300 ;
        RECT 164.400 240.150 165.600 248.400 ;
        RECT 206.100 243.000 207.900 251.250 ;
        RECT 131.100 237.150 132.900 238.950 ;
        RECT 163.950 238.050 166.050 240.150 ;
        RECT 166.950 239.850 169.050 241.950 ;
        RECT 203.400 241.350 207.900 243.000 ;
        RECT 211.500 242.400 213.300 251.250 ;
        RECT 248.100 243.000 249.900 251.250 ;
        RECT 245.400 241.350 249.900 243.000 ;
        RECT 253.500 242.400 255.300 251.250 ;
        RECT 287.550 248.400 289.350 251.250 ;
        RECT 288.150 244.500 289.350 248.400 ;
        RECT 290.850 245.400 292.650 251.250 ;
        RECT 293.850 245.400 295.650 251.250 ;
        RECT 330.150 246.900 331.950 251.250 ;
        RECT 328.650 245.400 331.950 246.900 ;
        RECT 333.150 245.400 334.950 251.250 ;
        RECT 288.150 243.600 293.250 244.500 ;
        RECT 291.000 242.700 293.250 243.600 ;
        RECT 167.100 238.050 168.900 239.850 ;
        RECT 127.950 233.850 130.050 235.950 ;
        RECT 130.950 235.050 133.050 237.150 ;
        RECT 35.400 219.750 37.200 225.600 ;
        RECT 38.700 219.750 40.500 231.600 ;
        RECT 42.900 219.750 44.700 231.600 ;
        RECT 80.400 219.750 82.200 225.600 ;
        RECT 83.700 219.750 85.500 231.600 ;
        RECT 87.900 219.750 89.700 231.600 ;
        RECT 128.250 225.600 129.450 233.850 ;
        RECT 164.400 225.600 165.600 238.050 ;
        RECT 203.400 237.150 204.600 241.350 ;
        RECT 245.400 237.150 246.600 241.350 ;
        RECT 202.950 235.050 205.050 237.150 ;
        RECT 203.250 226.800 204.300 235.050 ;
        RECT 205.950 233.850 208.050 235.950 ;
        RECT 211.950 233.850 214.050 235.950 ;
        RECT 244.950 235.050 247.050 237.150 ;
        RECT 286.950 236.850 289.050 238.950 ;
        RECT 205.950 232.050 207.750 233.850 ;
        RECT 208.950 230.850 211.050 232.950 ;
        RECT 212.100 232.050 213.900 233.850 ;
        RECT 209.100 229.050 210.900 230.850 ;
        RECT 245.250 226.800 246.300 235.050 ;
        RECT 247.950 233.850 250.050 235.950 ;
        RECT 253.950 233.850 256.050 235.950 ;
        RECT 287.100 235.050 288.900 236.850 ;
        RECT 291.000 234.300 292.050 242.700 ;
        RECT 294.150 238.950 295.350 245.400 ;
        RECT 292.950 236.850 295.350 238.950 ;
        RECT 247.950 232.050 249.750 233.850 ;
        RECT 250.950 230.850 253.050 232.950 ;
        RECT 254.100 232.050 255.900 233.850 ;
        RECT 291.000 233.400 293.250 234.300 ;
        RECT 287.550 232.500 293.250 233.400 ;
        RECT 251.100 229.050 252.900 230.850 ;
        RECT 203.250 225.900 210.300 226.800 ;
        RECT 203.250 225.600 204.450 225.900 ;
        RECT 124.650 219.750 126.450 225.600 ;
        RECT 127.650 219.750 129.450 225.600 ;
        RECT 130.650 219.750 132.450 225.600 ;
        RECT 163.650 219.750 165.450 225.600 ;
        RECT 166.650 219.750 168.450 225.600 ;
        RECT 202.650 219.750 204.450 225.600 ;
        RECT 208.650 225.600 210.300 225.900 ;
        RECT 245.250 225.900 252.300 226.800 ;
        RECT 245.250 225.600 246.450 225.900 ;
        RECT 205.650 219.750 207.450 225.000 ;
        RECT 208.650 219.750 210.450 225.600 ;
        RECT 211.650 219.750 213.450 225.600 ;
        RECT 244.650 219.750 246.450 225.600 ;
        RECT 250.650 225.600 252.300 225.900 ;
        RECT 287.550 225.600 288.750 232.500 ;
        RECT 294.150 231.600 295.350 236.850 ;
        RECT 328.650 238.950 329.850 245.400 ;
        RECT 331.950 243.900 333.750 244.500 ;
        RECT 337.650 243.900 339.450 251.250 ;
        RECT 371.550 246.300 373.350 251.250 ;
        RECT 374.550 247.200 376.350 251.250 ;
        RECT 377.550 246.300 379.350 251.250 ;
        RECT 371.550 244.950 379.350 246.300 ;
        RECT 380.550 245.400 382.350 251.250 ;
        RECT 418.650 245.400 420.450 251.250 ;
        RECT 331.950 242.700 339.450 243.900 ;
        RECT 380.550 243.300 381.750 245.400 ;
        RECT 328.650 236.850 331.050 238.950 ;
        RECT 332.100 237.150 333.900 238.950 ;
        RECT 328.650 231.600 329.850 236.850 ;
        RECT 331.950 235.050 334.050 237.150 ;
        RECT 247.650 219.750 249.450 225.000 ;
        RECT 250.650 219.750 252.450 225.600 ;
        RECT 253.650 219.750 255.450 225.600 ;
        RECT 287.550 219.750 289.350 225.600 ;
        RECT 290.850 219.750 292.650 231.600 ;
        RECT 293.850 219.750 295.650 231.600 ;
        RECT 328.050 219.750 329.850 231.600 ;
        RECT 331.050 219.750 332.850 231.600 ;
        RECT 335.100 225.600 336.300 242.700 ;
        RECT 378.000 242.250 381.750 243.300 ;
        RECT 419.250 243.300 420.450 245.400 ;
        RECT 421.650 246.300 423.450 251.250 ;
        RECT 424.650 247.200 426.450 251.250 ;
        RECT 427.650 246.300 429.450 251.250 ;
        RECT 461.550 248.400 463.350 251.250 ;
        RECT 464.550 248.400 466.350 251.250 ;
        RECT 467.550 248.400 469.350 251.250 ;
        RECT 421.650 244.950 429.450 246.300 ;
        RECT 465.450 244.200 466.350 248.400 ;
        RECT 470.550 245.400 472.350 251.250 ;
        RECT 465.450 243.300 468.750 244.200 ;
        RECT 419.250 242.250 423.000 243.300 ;
        RECT 466.950 242.400 468.750 243.300 ;
        RECT 374.100 240.150 375.900 241.950 ;
        RECT 337.950 236.850 340.050 238.950 ;
        RECT 370.950 236.850 373.050 238.950 ;
        RECT 373.950 238.050 376.050 240.150 ;
        RECT 377.850 238.950 379.050 242.250 ;
        RECT 379.950 240.450 382.050 241.050 ;
        RECT 412.950 240.450 415.050 241.050 ;
        RECT 379.950 239.550 415.050 240.450 ;
        RECT 379.950 238.950 382.050 239.550 ;
        RECT 412.950 238.950 415.050 239.550 ;
        RECT 421.950 238.950 423.150 242.250 ;
        RECT 425.100 240.150 426.900 241.950 ;
        RECT 376.950 236.850 379.050 238.950 ;
        RECT 421.950 236.850 424.050 238.950 ;
        RECT 424.950 238.050 427.050 240.150 ;
        RECT 460.950 239.850 463.050 241.950 ;
        RECT 427.950 236.850 430.050 238.950 ;
        RECT 461.100 238.050 462.900 239.850 ;
        RECT 463.950 236.850 466.050 238.950 ;
        RECT 338.100 235.050 339.900 236.850 ;
        RECT 371.100 235.050 372.900 236.850 ;
        RECT 376.950 231.600 378.150 236.850 ;
        RECT 379.950 233.850 382.050 235.950 ;
        RECT 418.950 233.850 421.050 235.950 ;
        RECT 379.950 232.050 381.750 233.850 ;
        RECT 419.250 232.050 421.050 233.850 ;
        RECT 422.850 231.600 424.050 236.850 ;
        RECT 428.100 235.050 429.900 236.850 ;
        RECT 464.100 235.050 465.900 236.850 ;
        RECT 467.700 234.150 468.600 242.400 ;
        RECT 471.000 240.150 472.050 245.400 ;
        RECT 509.850 244.200 511.650 251.250 ;
        RECT 514.350 245.400 516.150 251.250 ;
        RECT 548.550 248.400 550.350 251.250 ;
        RECT 551.550 248.400 553.350 251.250 ;
        RECT 509.850 243.300 513.450 244.200 ;
        RECT 469.950 238.050 472.050 240.150 ;
        RECT 466.950 234.000 468.750 234.150 ;
        RECT 461.550 232.800 468.750 234.000 ;
        RECT 461.550 231.600 462.750 232.800 ;
        RECT 466.950 232.350 468.750 232.800 ;
        RECT 334.650 219.750 336.450 225.600 ;
        RECT 337.650 219.750 339.450 225.600 ;
        RECT 372.300 219.750 374.100 231.600 ;
        RECT 376.500 219.750 378.300 231.600 ;
        RECT 379.800 219.750 381.600 225.600 ;
        RECT 419.400 219.750 421.200 225.600 ;
        RECT 422.700 219.750 424.500 231.600 ;
        RECT 426.900 219.750 428.700 231.600 ;
        RECT 461.550 219.750 463.350 231.600 ;
        RECT 470.100 231.450 471.450 238.050 ;
        RECT 509.100 237.150 510.900 238.950 ;
        RECT 508.950 235.050 511.050 237.150 ;
        RECT 512.250 235.950 513.450 243.300 ;
        RECT 547.950 239.850 550.050 241.950 ;
        RECT 551.400 240.150 552.600 248.400 ;
        RECT 587.550 246.300 589.350 251.250 ;
        RECT 590.550 247.200 592.350 251.250 ;
        RECT 593.550 246.300 595.350 251.250 ;
        RECT 587.550 244.950 595.350 246.300 ;
        RECT 596.550 245.400 598.350 251.250 ;
        RECT 596.550 243.300 597.750 245.400 ;
        RECT 632.850 244.200 634.650 251.250 ;
        RECT 637.350 245.400 639.150 251.250 ;
        RECT 642.150 245.400 643.950 251.250 ;
        RECT 645.150 248.400 646.950 251.250 ;
        RECT 649.950 249.300 651.750 251.250 ;
        RECT 648.000 248.400 651.750 249.300 ;
        RECT 654.450 248.400 656.250 251.250 ;
        RECT 657.750 248.400 659.550 251.250 ;
        RECT 661.650 248.400 663.450 251.250 ;
        RECT 665.850 248.400 667.650 251.250 ;
        RECT 670.350 248.400 672.150 251.250 ;
        RECT 648.000 247.500 649.050 248.400 ;
        RECT 646.950 245.400 649.050 247.500 ;
        RECT 657.750 246.600 658.800 248.400 ;
        RECT 632.850 243.300 636.450 244.200 ;
        RECT 594.000 242.250 597.750 243.300 ;
        RECT 590.100 240.150 591.900 241.950 ;
        RECT 515.100 237.150 516.900 238.950 ;
        RECT 548.100 238.050 549.900 239.850 ;
        RECT 550.950 238.050 553.050 240.150 ;
        RECT 511.950 233.850 514.050 235.950 ;
        RECT 514.950 235.050 517.050 237.150 ;
        RECT 466.050 219.750 467.850 231.450 ;
        RECT 469.050 230.100 471.450 231.450 ;
        RECT 469.050 219.750 470.850 230.100 ;
        RECT 512.250 225.600 513.450 233.850 ;
        RECT 551.400 225.600 552.600 238.050 ;
        RECT 586.950 236.850 589.050 238.950 ;
        RECT 589.950 238.050 592.050 240.150 ;
        RECT 593.850 238.950 595.050 242.250 ;
        RECT 592.950 236.850 595.050 238.950 ;
        RECT 632.100 237.150 633.900 238.950 ;
        RECT 587.100 235.050 588.900 236.850 ;
        RECT 592.950 231.600 594.150 236.850 ;
        RECT 595.950 233.850 598.050 235.950 ;
        RECT 631.950 235.050 634.050 237.150 ;
        RECT 635.250 235.950 636.450 243.300 ;
        RECT 638.100 237.150 639.900 238.950 ;
        RECT 634.950 233.850 637.050 235.950 ;
        RECT 637.950 235.050 640.050 237.150 ;
        RECT 595.950 232.050 597.750 233.850 ;
        RECT 508.650 219.750 510.450 225.600 ;
        RECT 511.650 219.750 513.450 225.600 ;
        RECT 514.650 219.750 516.450 225.600 ;
        RECT 548.550 219.750 550.350 225.600 ;
        RECT 551.550 219.750 553.350 225.600 ;
        RECT 588.300 219.750 590.100 231.600 ;
        RECT 592.500 219.750 594.300 231.600 ;
        RECT 635.250 225.600 636.450 233.850 ;
        RECT 642.150 232.800 643.050 245.400 ;
        RECT 650.550 244.800 652.350 246.600 ;
        RECT 653.850 245.550 658.800 246.600 ;
        RECT 666.300 247.500 667.350 248.400 ;
        RECT 666.300 246.300 670.050 247.500 ;
        RECT 653.850 244.800 655.650 245.550 ;
        RECT 650.850 243.900 651.900 244.800 ;
        RECT 661.050 244.200 662.850 246.000 ;
        RECT 667.950 245.400 670.050 246.300 ;
        RECT 673.650 245.400 675.450 251.250 ;
        RECT 661.050 243.900 661.950 244.200 ;
        RECT 650.850 243.000 661.950 243.900 ;
        RECT 674.250 243.150 675.450 245.400 ;
        RECT 707.550 246.300 709.350 251.250 ;
        RECT 710.550 247.200 712.350 251.250 ;
        RECT 713.550 246.300 715.350 251.250 ;
        RECT 707.550 244.950 715.350 246.300 ;
        RECT 716.550 245.400 718.350 251.250 ;
        RECT 749.850 245.400 751.650 251.250 ;
        RECT 716.550 243.300 717.750 245.400 ;
        RECT 754.350 244.200 756.150 251.250 ;
        RECT 650.850 241.800 651.900 243.000 ;
        RECT 645.000 240.600 651.900 241.800 ;
        RECT 645.000 239.850 645.900 240.600 ;
        RECT 650.100 240.000 651.900 240.600 ;
        RECT 644.100 238.050 645.900 239.850 ;
        RECT 647.100 238.950 648.900 239.700 ;
        RECT 661.050 238.950 661.950 243.000 ;
        RECT 670.950 241.050 675.450 243.150 ;
        RECT 714.000 242.250 717.750 243.300 ;
        RECT 752.550 243.300 756.150 244.200 ;
        RECT 669.150 239.250 673.050 241.050 ;
        RECT 670.950 238.950 673.050 239.250 ;
        RECT 647.100 237.900 655.050 238.950 ;
        RECT 652.950 236.850 655.050 237.900 ;
        RECT 658.950 236.850 661.950 238.950 ;
        RECT 651.450 233.100 653.250 233.400 ;
        RECT 651.450 232.800 659.850 233.100 ;
        RECT 642.150 232.200 659.850 232.800 ;
        RECT 642.150 231.600 653.250 232.200 ;
        RECT 595.800 219.750 597.600 225.600 ;
        RECT 631.650 219.750 633.450 225.600 ;
        RECT 634.650 219.750 636.450 225.600 ;
        RECT 637.650 219.750 639.450 225.600 ;
        RECT 642.150 219.750 643.950 231.600 ;
        RECT 656.250 230.700 658.050 231.300 ;
        RECT 650.550 229.500 658.050 230.700 ;
        RECT 658.950 230.100 659.850 232.200 ;
        RECT 661.050 232.200 661.950 236.850 ;
        RECT 671.250 233.400 673.050 235.200 ;
        RECT 667.950 232.200 672.150 233.400 ;
        RECT 661.050 231.300 667.050 232.200 ;
        RECT 667.950 231.300 670.050 232.200 ;
        RECT 674.250 231.600 675.450 241.050 ;
        RECT 710.100 240.150 711.900 241.950 ;
        RECT 706.950 236.850 709.050 238.950 ;
        RECT 709.950 238.050 712.050 240.150 ;
        RECT 713.850 238.950 715.050 242.250 ;
        RECT 712.950 236.850 715.050 238.950 ;
        RECT 749.100 237.150 750.900 238.950 ;
        RECT 707.100 235.050 708.900 236.850 ;
        RECT 712.950 231.600 714.150 236.850 ;
        RECT 715.950 233.850 718.050 235.950 ;
        RECT 748.950 235.050 751.050 237.150 ;
        RECT 752.550 235.950 753.750 243.300 ;
        RECT 755.100 237.150 756.900 238.950 ;
        RECT 751.950 233.850 754.050 235.950 ;
        RECT 754.950 235.050 757.050 237.150 ;
        RECT 715.950 232.050 717.750 233.850 ;
        RECT 666.150 230.400 667.050 231.300 ;
        RECT 663.450 230.100 665.250 230.400 ;
        RECT 650.550 228.600 651.750 229.500 ;
        RECT 658.950 229.200 665.250 230.100 ;
        RECT 663.450 228.600 665.250 229.200 ;
        RECT 666.150 228.600 668.850 230.400 ;
        RECT 646.950 226.500 651.750 228.600 ;
        RECT 654.150 226.500 661.050 228.300 ;
        RECT 650.550 225.600 651.750 226.500 ;
        RECT 645.150 219.750 646.950 225.600 ;
        RECT 650.250 219.750 652.050 225.600 ;
        RECT 655.050 219.750 656.850 225.600 ;
        RECT 658.050 219.750 659.850 226.500 ;
        RECT 666.150 225.600 670.050 227.700 ;
        RECT 661.950 219.750 663.750 225.600 ;
        RECT 666.150 219.750 667.950 225.600 ;
        RECT 670.650 219.750 672.450 222.600 ;
        RECT 673.650 219.750 675.450 231.600 ;
        RECT 708.300 219.750 710.100 231.600 ;
        RECT 712.500 219.750 714.300 231.600 ;
        RECT 752.550 225.600 753.750 233.850 ;
        RECT 715.800 219.750 717.600 225.600 ;
        RECT 749.550 219.750 751.350 225.600 ;
        RECT 752.550 219.750 754.350 225.600 ;
        RECT 755.550 219.750 757.350 225.600 ;
        RECT 34.650 203.400 36.450 215.250 ;
        RECT 37.650 202.500 39.450 215.250 ;
        RECT 40.650 203.400 42.450 215.250 ;
        RECT 43.650 202.500 45.450 215.250 ;
        RECT 46.650 203.400 48.450 215.250 ;
        RECT 49.650 202.500 51.450 215.250 ;
        RECT 52.650 203.400 54.450 215.250 ;
        RECT 55.650 202.500 57.450 215.250 ;
        RECT 58.650 203.400 60.450 215.250 ;
        RECT 94.650 209.400 96.450 215.250 ;
        RECT 97.650 209.400 99.450 215.250 ;
        RECT 100.650 209.400 102.450 215.250 ;
        RECT 36.750 201.300 39.450 202.500 ;
        RECT 41.700 201.300 45.450 202.500 ;
        RECT 47.700 201.300 51.450 202.500 ;
        RECT 53.550 201.300 57.450 202.500 ;
        RECT 36.750 196.950 37.800 201.300 ;
        RECT 34.950 194.850 37.800 196.950 ;
        RECT 36.750 191.700 37.800 194.850 ;
        RECT 41.700 194.400 42.900 201.300 ;
        RECT 47.700 194.400 48.900 201.300 ;
        RECT 53.550 194.400 54.750 201.300 ;
        RECT 98.250 201.150 99.450 209.400 ;
        RECT 105.150 203.400 106.950 215.250 ;
        RECT 108.150 209.400 109.950 215.250 ;
        RECT 113.250 209.400 115.050 215.250 ;
        RECT 118.050 209.400 119.850 215.250 ;
        RECT 113.550 208.500 114.750 209.400 ;
        RECT 121.050 208.500 122.850 215.250 ;
        RECT 124.950 209.400 126.750 215.250 ;
        RECT 129.150 209.400 130.950 215.250 ;
        RECT 133.650 212.400 135.450 215.250 ;
        RECT 109.950 206.400 114.750 208.500 ;
        RECT 117.150 206.700 124.050 208.500 ;
        RECT 129.150 207.300 133.050 209.400 ;
        RECT 113.550 205.500 114.750 206.400 ;
        RECT 126.450 205.800 128.250 206.400 ;
        RECT 113.550 204.300 121.050 205.500 ;
        RECT 119.250 203.700 121.050 204.300 ;
        RECT 121.950 204.900 128.250 205.800 ;
        RECT 105.150 202.800 116.250 203.400 ;
        RECT 121.950 202.800 122.850 204.900 ;
        RECT 126.450 204.600 128.250 204.900 ;
        RECT 129.150 204.600 131.850 206.400 ;
        RECT 129.150 203.700 130.050 204.600 ;
        RECT 105.150 202.200 122.850 202.800 ;
        RECT 94.950 197.850 97.050 199.950 ;
        RECT 97.950 199.050 100.050 201.150 ;
        RECT 55.950 194.850 58.050 196.950 ;
        RECT 95.100 196.050 96.900 197.850 ;
        RECT 38.700 192.600 42.900 194.400 ;
        RECT 44.700 192.600 48.900 194.400 ;
        RECT 50.700 192.600 54.750 194.400 ;
        RECT 56.100 193.050 57.900 194.850 ;
        RECT 41.700 191.700 42.900 192.600 ;
        RECT 47.700 191.700 48.900 192.600 ;
        RECT 53.550 191.700 54.750 192.600 ;
        RECT 98.250 191.700 99.450 199.050 ;
        RECT 100.950 197.850 103.050 199.950 ;
        RECT 101.100 196.050 102.900 197.850 ;
        RECT 36.750 190.650 39.600 191.700 ;
        RECT 36.900 190.500 39.600 190.650 ;
        RECT 41.700 190.500 45.600 191.700 ;
        RECT 47.700 190.500 51.450 191.700 ;
        RECT 53.550 190.500 57.600 191.700 ;
        RECT 37.800 189.600 39.600 190.500 ;
        RECT 43.800 189.600 45.600 190.500 ;
        RECT 34.650 183.750 36.450 189.600 ;
        RECT 37.650 183.750 39.450 189.600 ;
        RECT 40.650 183.750 42.450 189.600 ;
        RECT 43.650 183.750 45.450 189.600 ;
        RECT 46.650 183.750 48.450 189.600 ;
        RECT 49.650 183.750 51.450 190.500 ;
        RECT 55.800 189.600 57.600 190.500 ;
        RECT 95.850 190.800 99.450 191.700 ;
        RECT 52.650 183.750 54.450 189.600 ;
        RECT 55.650 183.750 57.450 189.600 ;
        RECT 58.650 183.750 60.450 189.600 ;
        RECT 95.850 183.750 97.650 190.800 ;
        RECT 105.150 189.600 106.050 202.200 ;
        RECT 114.450 201.900 122.850 202.200 ;
        RECT 124.050 202.800 130.050 203.700 ;
        RECT 130.950 202.800 133.050 203.700 ;
        RECT 136.650 203.400 138.450 215.250 ;
        RECT 173.400 209.400 175.200 215.250 ;
        RECT 176.700 203.400 178.500 215.250 ;
        RECT 180.900 203.400 182.700 215.250 ;
        RECT 215.550 209.400 217.350 215.250 ;
        RECT 218.550 209.400 220.350 215.250 ;
        RECT 221.550 210.000 223.350 215.250 ;
        RECT 218.700 209.100 220.350 209.400 ;
        RECT 224.550 209.400 226.350 215.250 ;
        RECT 260.550 209.400 262.350 215.250 ;
        RECT 263.550 209.400 265.350 215.250 ;
        RECT 266.550 209.400 268.350 215.250 ;
        RECT 302.550 209.400 304.350 215.250 ;
        RECT 224.550 209.100 225.750 209.400 ;
        RECT 218.700 208.200 225.750 209.100 ;
        RECT 218.100 204.150 219.900 205.950 ;
        RECT 114.450 201.600 116.250 201.900 ;
        RECT 124.050 198.150 124.950 202.800 ;
        RECT 130.950 201.600 135.150 202.800 ;
        RECT 134.250 199.800 136.050 201.600 ;
        RECT 115.950 197.100 118.050 198.150 ;
        RECT 107.100 195.150 108.900 196.950 ;
        RECT 110.100 196.050 118.050 197.100 ;
        RECT 121.950 196.050 124.950 198.150 ;
        RECT 110.100 195.300 111.900 196.050 ;
        RECT 108.000 194.400 108.900 195.150 ;
        RECT 113.100 194.400 114.900 195.000 ;
        RECT 108.000 193.200 114.900 194.400 ;
        RECT 113.850 192.000 114.900 193.200 ;
        RECT 124.050 192.000 124.950 196.050 ;
        RECT 133.950 195.750 136.050 196.050 ;
        RECT 132.150 193.950 136.050 195.750 ;
        RECT 137.250 193.950 138.450 203.400 ;
        RECT 173.250 201.150 175.050 202.950 ;
        RECT 172.950 199.050 175.050 201.150 ;
        RECT 176.850 198.150 178.050 203.400 ;
        RECT 215.100 201.150 216.900 202.950 ;
        RECT 217.950 202.050 220.050 204.150 ;
        RECT 221.250 201.150 223.050 202.950 ;
        RECT 182.100 198.150 183.900 199.950 ;
        RECT 214.950 199.050 217.050 201.150 ;
        RECT 220.950 199.050 223.050 201.150 ;
        RECT 224.700 199.950 225.750 208.200 ;
        RECT 263.550 201.150 264.750 209.400 ;
        RECT 302.550 202.500 303.750 209.400 ;
        RECT 305.850 203.400 307.650 215.250 ;
        RECT 308.850 203.400 310.650 215.250 ;
        RECT 344.550 209.400 346.350 215.250 ;
        RECT 347.550 209.400 349.350 215.250 ;
        RECT 350.550 209.400 352.350 215.250 ;
        RECT 383.550 209.400 385.350 215.250 ;
        RECT 302.550 201.600 308.250 202.500 ;
        RECT 113.850 191.100 124.950 192.000 ;
        RECT 133.950 191.850 138.450 193.950 ;
        RECT 175.950 196.050 178.050 198.150 ;
        RECT 175.950 192.750 177.150 196.050 ;
        RECT 178.950 194.850 181.050 196.950 ;
        RECT 181.950 196.050 184.050 198.150 ;
        RECT 223.950 197.850 226.050 199.950 ;
        RECT 259.950 197.850 262.050 199.950 ;
        RECT 262.950 199.050 265.050 201.150 ;
        RECT 306.000 200.700 308.250 201.600 ;
        RECT 179.100 193.050 180.900 194.850 ;
        RECT 224.400 193.650 225.600 197.850 ;
        RECT 260.100 196.050 261.900 197.850 ;
        RECT 113.850 190.200 114.900 191.100 ;
        RECT 124.050 190.800 124.950 191.100 ;
        RECT 100.350 183.750 102.150 189.600 ;
        RECT 105.150 183.750 106.950 189.600 ;
        RECT 109.950 187.500 112.050 189.600 ;
        RECT 113.550 188.400 115.350 190.200 ;
        RECT 116.850 189.450 118.650 190.200 ;
        RECT 116.850 188.400 121.800 189.450 ;
        RECT 124.050 189.000 125.850 190.800 ;
        RECT 137.250 189.600 138.450 191.850 ;
        RECT 173.250 191.700 177.000 192.750 ;
        RECT 173.250 189.600 174.450 191.700 ;
        RECT 130.950 188.700 133.050 189.600 ;
        RECT 111.000 186.600 112.050 187.500 ;
        RECT 120.750 186.600 121.800 188.400 ;
        RECT 129.300 187.500 133.050 188.700 ;
        RECT 129.300 186.600 130.350 187.500 ;
        RECT 108.150 183.750 109.950 186.600 ;
        RECT 111.000 185.700 114.750 186.600 ;
        RECT 112.950 183.750 114.750 185.700 ;
        RECT 117.450 183.750 119.250 186.600 ;
        RECT 120.750 183.750 122.550 186.600 ;
        RECT 124.650 183.750 126.450 186.600 ;
        RECT 128.850 183.750 130.650 186.600 ;
        RECT 133.350 183.750 135.150 186.600 ;
        RECT 136.650 183.750 138.450 189.600 ;
        RECT 172.650 183.750 174.450 189.600 ;
        RECT 175.650 188.700 183.450 190.050 ;
        RECT 175.650 183.750 177.450 188.700 ;
        RECT 178.650 183.750 180.450 187.800 ;
        RECT 181.650 183.750 183.450 188.700 ;
        RECT 215.700 183.750 217.500 192.600 ;
        RECT 221.100 192.000 225.600 193.650 ;
        RECT 221.100 183.750 222.900 192.000 ;
        RECT 263.550 191.700 264.750 199.050 ;
        RECT 265.950 197.850 268.050 199.950 ;
        RECT 302.100 198.150 303.900 199.950 ;
        RECT 266.100 196.050 267.900 197.850 ;
        RECT 301.950 196.050 304.050 198.150 ;
        RECT 306.000 192.300 307.050 200.700 ;
        RECT 309.150 198.150 310.350 203.400 ;
        RECT 347.550 201.150 348.750 209.400 ;
        RECT 383.550 202.500 384.750 209.400 ;
        RECT 386.850 203.400 388.650 215.250 ;
        RECT 389.850 203.400 391.650 215.250 ;
        RECT 426.450 203.400 428.250 215.250 ;
        RECT 430.650 203.400 432.450 215.250 ;
        RECT 467.400 209.400 469.200 215.250 ;
        RECT 470.700 203.400 472.500 215.250 ;
        RECT 474.900 203.400 476.700 215.250 ;
        RECT 511.650 209.400 513.450 215.250 ;
        RECT 514.650 209.400 516.450 215.250 ;
        RECT 517.650 209.400 519.450 215.250 ;
        RECT 551.550 209.400 553.350 215.250 ;
        RECT 554.550 209.400 556.350 215.250 ;
        RECT 557.550 210.000 559.350 215.250 ;
        RECT 383.550 201.600 389.250 202.500 ;
        RECT 307.950 196.050 310.350 198.150 ;
        RECT 343.950 197.850 346.050 199.950 ;
        RECT 346.950 199.050 349.050 201.150 ;
        RECT 387.000 200.700 389.250 201.600 ;
        RECT 344.100 196.050 345.900 197.850 ;
        RECT 263.550 190.800 267.150 191.700 ;
        RECT 306.000 191.400 308.250 192.300 ;
        RECT 260.850 183.750 262.650 189.600 ;
        RECT 265.350 183.750 267.150 190.800 ;
        RECT 303.150 190.500 308.250 191.400 ;
        RECT 303.150 186.600 304.350 190.500 ;
        RECT 309.150 189.600 310.350 196.050 ;
        RECT 347.550 191.700 348.750 199.050 ;
        RECT 349.950 197.850 352.050 199.950 ;
        RECT 383.100 198.150 384.900 199.950 ;
        RECT 350.100 196.050 351.900 197.850 ;
        RECT 382.950 196.050 385.050 198.150 ;
        RECT 387.000 192.300 388.050 200.700 ;
        RECT 390.150 198.150 391.350 203.400 ;
        RECT 426.450 202.350 429.000 203.400 ;
        RECT 425.100 198.150 426.900 199.950 ;
        RECT 388.950 196.050 391.350 198.150 ;
        RECT 424.950 196.050 427.050 198.150 ;
        RECT 347.550 190.800 351.150 191.700 ;
        RECT 387.000 191.400 389.250 192.300 ;
        RECT 302.550 183.750 304.350 186.600 ;
        RECT 305.850 183.750 307.650 189.600 ;
        RECT 308.850 183.750 310.650 189.600 ;
        RECT 344.850 183.750 346.650 189.600 ;
        RECT 349.350 183.750 351.150 190.800 ;
        RECT 384.150 190.500 389.250 191.400 ;
        RECT 384.150 186.600 385.350 190.500 ;
        RECT 390.150 189.600 391.350 196.050 ;
        RECT 427.950 195.150 429.000 202.350 ;
        RECT 467.250 201.150 469.050 202.950 ;
        RECT 431.100 198.150 432.900 199.950 ;
        RECT 466.950 199.050 469.050 201.150 ;
        RECT 470.850 198.150 472.050 203.400 ;
        RECT 515.250 201.150 516.450 209.400 ;
        RECT 554.700 209.100 556.350 209.400 ;
        RECT 560.550 209.400 562.350 215.250 ;
        RECT 560.550 209.100 561.750 209.400 ;
        RECT 554.700 208.200 561.750 209.100 ;
        RECT 554.100 204.150 555.900 205.950 ;
        RECT 551.100 201.150 552.900 202.950 ;
        RECT 553.950 202.050 556.050 204.150 ;
        RECT 557.250 201.150 559.050 202.950 ;
        RECT 476.100 198.150 477.900 199.950 ;
        RECT 430.950 196.050 433.050 198.150 ;
        RECT 469.950 196.050 472.050 198.150 ;
        RECT 427.950 193.050 430.050 195.150 ;
        RECT 383.550 183.750 385.350 186.600 ;
        RECT 386.850 183.750 388.650 189.600 ;
        RECT 389.850 183.750 391.650 189.600 ;
        RECT 427.950 186.600 429.000 193.050 ;
        RECT 469.950 192.750 471.150 196.050 ;
        RECT 472.950 194.850 475.050 196.950 ;
        RECT 475.950 196.050 478.050 198.150 ;
        RECT 511.950 197.850 514.050 199.950 ;
        RECT 514.950 199.050 517.050 201.150 ;
        RECT 512.100 196.050 513.900 197.850 ;
        RECT 473.100 193.050 474.900 194.850 ;
        RECT 467.250 191.700 471.000 192.750 ;
        RECT 515.250 191.700 516.450 199.050 ;
        RECT 517.950 197.850 520.050 199.950 ;
        RECT 550.950 199.050 553.050 201.150 ;
        RECT 556.950 199.050 559.050 201.150 ;
        RECT 560.700 199.950 561.750 208.200 ;
        RECT 566.550 203.400 568.350 215.250 ;
        RECT 569.550 212.400 571.350 215.250 ;
        RECT 574.050 209.400 575.850 215.250 ;
        RECT 578.250 209.400 580.050 215.250 ;
        RECT 571.950 207.300 575.850 209.400 ;
        RECT 582.150 208.500 583.950 215.250 ;
        RECT 585.150 209.400 586.950 215.250 ;
        RECT 589.950 209.400 591.750 215.250 ;
        RECT 595.050 209.400 596.850 215.250 ;
        RECT 590.250 208.500 591.450 209.400 ;
        RECT 580.950 206.700 587.850 208.500 ;
        RECT 590.250 206.400 595.050 208.500 ;
        RECT 573.150 204.600 575.850 206.400 ;
        RECT 576.750 205.800 578.550 206.400 ;
        RECT 576.750 204.900 583.050 205.800 ;
        RECT 590.250 205.500 591.450 206.400 ;
        RECT 576.750 204.600 578.550 204.900 ;
        RECT 574.950 203.700 575.850 204.600 ;
        RECT 559.950 197.850 562.050 199.950 ;
        RECT 518.100 196.050 519.900 197.850 ;
        RECT 560.400 193.650 561.600 197.850 ;
        RECT 467.250 189.600 468.450 191.700 ;
        RECT 512.850 190.800 516.450 191.700 ;
        RECT 424.650 183.750 426.450 186.600 ;
        RECT 427.650 183.750 429.450 186.600 ;
        RECT 430.650 183.750 432.450 186.600 ;
        RECT 466.650 183.750 468.450 189.600 ;
        RECT 469.650 188.700 477.450 190.050 ;
        RECT 469.650 183.750 471.450 188.700 ;
        RECT 472.650 183.750 474.450 187.800 ;
        RECT 475.650 183.750 477.450 188.700 ;
        RECT 512.850 183.750 514.650 190.800 ;
        RECT 517.350 183.750 519.150 189.600 ;
        RECT 551.700 183.750 553.500 192.600 ;
        RECT 557.100 192.000 561.600 193.650 ;
        RECT 566.550 193.950 567.750 203.400 ;
        RECT 571.950 202.800 574.050 203.700 ;
        RECT 574.950 202.800 580.950 203.700 ;
        RECT 569.850 201.600 574.050 202.800 ;
        RECT 568.950 199.800 570.750 201.600 ;
        RECT 580.050 198.150 580.950 202.800 ;
        RECT 582.150 202.800 583.050 204.900 ;
        RECT 583.950 204.300 591.450 205.500 ;
        RECT 583.950 203.700 585.750 204.300 ;
        RECT 598.050 203.400 599.850 215.250 ;
        RECT 632.550 209.400 634.350 215.250 ;
        RECT 635.550 209.400 637.350 215.250 ;
        RECT 638.550 209.400 640.350 215.250 ;
        RECT 588.750 202.800 599.850 203.400 ;
        RECT 582.150 202.200 599.850 202.800 ;
        RECT 582.150 201.900 590.550 202.200 ;
        RECT 588.750 201.600 590.550 201.900 ;
        RECT 580.050 196.050 583.050 198.150 ;
        RECT 586.950 197.100 589.050 198.150 ;
        RECT 586.950 196.050 594.900 197.100 ;
        RECT 568.950 195.750 571.050 196.050 ;
        RECT 568.950 193.950 572.850 195.750 ;
        RECT 557.100 183.750 558.900 192.000 ;
        RECT 566.550 191.850 571.050 193.950 ;
        RECT 580.050 192.000 580.950 196.050 ;
        RECT 593.100 195.300 594.900 196.050 ;
        RECT 596.100 195.150 597.900 196.950 ;
        RECT 590.100 194.400 591.900 195.000 ;
        RECT 596.100 194.400 597.000 195.150 ;
        RECT 590.100 193.200 597.000 194.400 ;
        RECT 590.100 192.000 591.150 193.200 ;
        RECT 566.550 189.600 567.750 191.850 ;
        RECT 580.050 191.100 591.150 192.000 ;
        RECT 580.050 190.800 580.950 191.100 ;
        RECT 566.550 183.750 568.350 189.600 ;
        RECT 571.950 188.700 574.050 189.600 ;
        RECT 579.150 189.000 580.950 190.800 ;
        RECT 590.100 190.200 591.150 191.100 ;
        RECT 586.350 189.450 588.150 190.200 ;
        RECT 571.950 187.500 575.700 188.700 ;
        RECT 574.650 186.600 575.700 187.500 ;
        RECT 583.200 188.400 588.150 189.450 ;
        RECT 589.650 188.400 591.450 190.200 ;
        RECT 598.950 189.600 599.850 202.200 ;
        RECT 635.550 201.150 636.750 209.400 ;
        RECT 645.150 203.400 646.950 215.250 ;
        RECT 648.150 209.400 649.950 215.250 ;
        RECT 653.250 209.400 655.050 215.250 ;
        RECT 658.050 209.400 659.850 215.250 ;
        RECT 653.550 208.500 654.750 209.400 ;
        RECT 661.050 208.500 662.850 215.250 ;
        RECT 664.950 209.400 666.750 215.250 ;
        RECT 669.150 209.400 670.950 215.250 ;
        RECT 673.650 212.400 675.450 215.250 ;
        RECT 649.950 206.400 654.750 208.500 ;
        RECT 657.150 206.700 664.050 208.500 ;
        RECT 669.150 207.300 673.050 209.400 ;
        RECT 653.550 205.500 654.750 206.400 ;
        RECT 666.450 205.800 668.250 206.400 ;
        RECT 653.550 204.300 661.050 205.500 ;
        RECT 659.250 203.700 661.050 204.300 ;
        RECT 661.950 204.900 668.250 205.800 ;
        RECT 645.150 202.800 656.250 203.400 ;
        RECT 661.950 202.800 662.850 204.900 ;
        RECT 666.450 204.600 668.250 204.900 ;
        RECT 669.150 204.600 671.850 206.400 ;
        RECT 669.150 203.700 670.050 204.600 ;
        RECT 645.150 202.200 662.850 202.800 ;
        RECT 631.950 197.850 634.050 199.950 ;
        RECT 634.950 199.050 637.050 201.150 ;
        RECT 632.100 196.050 633.900 197.850 ;
        RECT 635.550 191.700 636.750 199.050 ;
        RECT 637.950 197.850 640.050 199.950 ;
        RECT 638.100 196.050 639.900 197.850 ;
        RECT 635.550 190.800 639.150 191.700 ;
        RECT 583.200 186.600 584.250 188.400 ;
        RECT 592.950 187.500 595.050 189.600 ;
        RECT 592.950 186.600 594.000 187.500 ;
        RECT 569.850 183.750 571.650 186.600 ;
        RECT 574.350 183.750 576.150 186.600 ;
        RECT 578.550 183.750 580.350 186.600 ;
        RECT 582.450 183.750 584.250 186.600 ;
        RECT 585.750 183.750 587.550 186.600 ;
        RECT 590.250 185.700 594.000 186.600 ;
        RECT 590.250 183.750 592.050 185.700 ;
        RECT 595.050 183.750 596.850 186.600 ;
        RECT 598.050 183.750 599.850 189.600 ;
        RECT 632.850 183.750 634.650 189.600 ;
        RECT 637.350 183.750 639.150 190.800 ;
        RECT 645.150 189.600 646.050 202.200 ;
        RECT 654.450 201.900 662.850 202.200 ;
        RECT 664.050 202.800 670.050 203.700 ;
        RECT 670.950 202.800 673.050 203.700 ;
        RECT 676.650 203.400 678.450 215.250 ;
        RECT 708.300 203.400 710.100 215.250 ;
        RECT 712.500 203.400 714.300 215.250 ;
        RECT 715.800 209.400 717.600 215.250 ;
        RECT 723.150 203.400 724.950 215.250 ;
        RECT 726.150 209.400 727.950 215.250 ;
        RECT 731.250 209.400 733.050 215.250 ;
        RECT 736.050 209.400 737.850 215.250 ;
        RECT 731.550 208.500 732.750 209.400 ;
        RECT 739.050 208.500 740.850 215.250 ;
        RECT 742.950 209.400 744.750 215.250 ;
        RECT 747.150 209.400 748.950 215.250 ;
        RECT 751.650 212.400 753.450 215.250 ;
        RECT 727.950 206.400 732.750 208.500 ;
        RECT 735.150 206.700 742.050 208.500 ;
        RECT 747.150 207.300 751.050 209.400 ;
        RECT 731.550 205.500 732.750 206.400 ;
        RECT 744.450 205.800 746.250 206.400 ;
        RECT 731.550 204.300 739.050 205.500 ;
        RECT 737.250 203.700 739.050 204.300 ;
        RECT 739.950 204.900 746.250 205.800 ;
        RECT 654.450 201.600 656.250 201.900 ;
        RECT 664.050 198.150 664.950 202.800 ;
        RECT 670.950 201.600 675.150 202.800 ;
        RECT 674.250 199.800 676.050 201.600 ;
        RECT 655.950 197.100 658.050 198.150 ;
        RECT 647.100 195.150 648.900 196.950 ;
        RECT 650.100 196.050 658.050 197.100 ;
        RECT 661.950 196.050 664.950 198.150 ;
        RECT 650.100 195.300 651.900 196.050 ;
        RECT 648.000 194.400 648.900 195.150 ;
        RECT 653.100 194.400 654.900 195.000 ;
        RECT 648.000 193.200 654.900 194.400 ;
        RECT 653.850 192.000 654.900 193.200 ;
        RECT 664.050 192.000 664.950 196.050 ;
        RECT 673.950 195.750 676.050 196.050 ;
        RECT 672.150 193.950 676.050 195.750 ;
        RECT 677.250 193.950 678.450 203.400 ;
        RECT 707.100 198.150 708.900 199.950 ;
        RECT 712.950 198.150 714.150 203.400 ;
        RECT 715.950 201.150 717.750 202.950 ;
        RECT 723.150 202.800 734.250 203.400 ;
        RECT 739.950 202.800 740.850 204.900 ;
        RECT 744.450 204.600 746.250 204.900 ;
        RECT 747.150 204.600 749.850 206.400 ;
        RECT 747.150 203.700 748.050 204.600 ;
        RECT 723.150 202.200 740.850 202.800 ;
        RECT 715.950 199.050 718.050 201.150 ;
        RECT 706.950 196.050 709.050 198.150 ;
        RECT 709.950 194.850 712.050 196.950 ;
        RECT 712.950 196.050 715.050 198.150 ;
        RECT 653.850 191.100 664.950 192.000 ;
        RECT 673.950 191.850 678.450 193.950 ;
        RECT 710.100 193.050 711.900 194.850 ;
        RECT 713.850 192.750 715.050 196.050 ;
        RECT 653.850 190.200 654.900 191.100 ;
        RECT 664.050 190.800 664.950 191.100 ;
        RECT 645.150 183.750 646.950 189.600 ;
        RECT 649.950 187.500 652.050 189.600 ;
        RECT 653.550 188.400 655.350 190.200 ;
        RECT 656.850 189.450 658.650 190.200 ;
        RECT 656.850 188.400 661.800 189.450 ;
        RECT 664.050 189.000 665.850 190.800 ;
        RECT 677.250 189.600 678.450 191.850 ;
        RECT 714.000 191.700 717.750 192.750 ;
        RECT 670.950 188.700 673.050 189.600 ;
        RECT 651.000 186.600 652.050 187.500 ;
        RECT 660.750 186.600 661.800 188.400 ;
        RECT 669.300 187.500 673.050 188.700 ;
        RECT 669.300 186.600 670.350 187.500 ;
        RECT 648.150 183.750 649.950 186.600 ;
        RECT 651.000 185.700 654.750 186.600 ;
        RECT 652.950 183.750 654.750 185.700 ;
        RECT 657.450 183.750 659.250 186.600 ;
        RECT 660.750 183.750 662.550 186.600 ;
        RECT 664.650 183.750 666.450 186.600 ;
        RECT 668.850 183.750 670.650 186.600 ;
        RECT 673.350 183.750 675.150 186.600 ;
        RECT 676.650 183.750 678.450 189.600 ;
        RECT 707.550 188.700 715.350 190.050 ;
        RECT 707.550 183.750 709.350 188.700 ;
        RECT 710.550 183.750 712.350 187.800 ;
        RECT 713.550 183.750 715.350 188.700 ;
        RECT 716.550 189.600 717.750 191.700 ;
        RECT 723.150 189.600 724.050 202.200 ;
        RECT 732.450 201.900 740.850 202.200 ;
        RECT 742.050 202.800 748.050 203.700 ;
        RECT 748.950 202.800 751.050 203.700 ;
        RECT 754.650 203.400 756.450 215.250 ;
        RECT 732.450 201.600 734.250 201.900 ;
        RECT 742.050 198.150 742.950 202.800 ;
        RECT 748.950 201.600 753.150 202.800 ;
        RECT 752.250 199.800 754.050 201.600 ;
        RECT 733.950 197.100 736.050 198.150 ;
        RECT 725.100 195.150 726.900 196.950 ;
        RECT 728.100 196.050 736.050 197.100 ;
        RECT 739.950 196.050 742.950 198.150 ;
        RECT 728.100 195.300 729.900 196.050 ;
        RECT 726.000 194.400 726.900 195.150 ;
        RECT 731.100 194.400 732.900 195.000 ;
        RECT 726.000 193.200 732.900 194.400 ;
        RECT 731.850 192.000 732.900 193.200 ;
        RECT 742.050 192.000 742.950 196.050 ;
        RECT 751.950 195.750 754.050 196.050 ;
        RECT 750.150 193.950 754.050 195.750 ;
        RECT 755.250 193.950 756.450 203.400 ;
        RECT 731.850 191.100 742.950 192.000 ;
        RECT 751.950 191.850 756.450 193.950 ;
        RECT 731.850 190.200 732.900 191.100 ;
        RECT 742.050 190.800 742.950 191.100 ;
        RECT 716.550 183.750 718.350 189.600 ;
        RECT 723.150 183.750 724.950 189.600 ;
        RECT 727.950 187.500 730.050 189.600 ;
        RECT 731.550 188.400 733.350 190.200 ;
        RECT 734.850 189.450 736.650 190.200 ;
        RECT 734.850 188.400 739.800 189.450 ;
        RECT 742.050 189.000 743.850 190.800 ;
        RECT 755.250 189.600 756.450 191.850 ;
        RECT 748.950 188.700 751.050 189.600 ;
        RECT 729.000 186.600 730.050 187.500 ;
        RECT 738.750 186.600 739.800 188.400 ;
        RECT 747.300 187.500 751.050 188.700 ;
        RECT 747.300 186.600 748.350 187.500 ;
        RECT 726.150 183.750 727.950 186.600 ;
        RECT 729.000 185.700 732.750 186.600 ;
        RECT 730.950 183.750 732.750 185.700 ;
        RECT 735.450 183.750 737.250 186.600 ;
        RECT 738.750 183.750 740.550 186.600 ;
        RECT 742.650 183.750 744.450 186.600 ;
        RECT 746.850 183.750 748.650 186.600 ;
        RECT 751.350 183.750 753.150 186.600 ;
        RECT 754.650 183.750 756.450 189.600 ;
        RECT 32.550 173.400 34.350 179.250 ;
        RECT 35.550 173.400 37.350 179.250 ;
        RECT 68.550 174.300 70.350 179.250 ;
        RECT 71.550 175.200 73.350 179.250 ;
        RECT 74.550 174.300 76.350 179.250 ;
        RECT 32.100 168.150 33.900 169.950 ;
        RECT 31.950 166.050 34.050 168.150 ;
        RECT 35.400 166.950 36.600 173.400 ;
        RECT 68.550 172.950 76.350 174.300 ;
        RECT 77.550 173.400 79.350 179.250 ;
        RECT 84.150 173.400 85.950 179.250 ;
        RECT 87.150 176.400 88.950 179.250 ;
        RECT 91.950 177.300 93.750 179.250 ;
        RECT 90.000 176.400 93.750 177.300 ;
        RECT 96.450 176.400 98.250 179.250 ;
        RECT 99.750 176.400 101.550 179.250 ;
        RECT 103.650 176.400 105.450 179.250 ;
        RECT 107.850 176.400 109.650 179.250 ;
        RECT 112.350 176.400 114.150 179.250 ;
        RECT 90.000 175.500 91.050 176.400 ;
        RECT 88.950 173.400 91.050 175.500 ;
        RECT 99.750 174.600 100.800 176.400 ;
        RECT 77.550 171.300 78.750 173.400 ;
        RECT 75.000 170.250 78.750 171.300 ;
        RECT 71.100 168.150 72.900 169.950 ;
        RECT 34.950 164.850 37.050 166.950 ;
        RECT 67.950 164.850 70.050 166.950 ;
        RECT 70.950 166.050 73.050 168.150 ;
        RECT 74.850 166.950 76.050 170.250 ;
        RECT 73.950 164.850 76.050 166.950 ;
        RECT 35.400 159.600 36.600 164.850 ;
        RECT 68.100 163.050 69.900 164.850 ;
        RECT 73.950 159.600 75.150 164.850 ;
        RECT 76.950 161.850 79.050 163.950 ;
        RECT 76.950 160.050 78.750 161.850 ;
        RECT 84.150 160.800 85.050 173.400 ;
        RECT 92.550 172.800 94.350 174.600 ;
        RECT 95.850 173.550 100.800 174.600 ;
        RECT 108.300 175.500 109.350 176.400 ;
        RECT 108.300 174.300 112.050 175.500 ;
        RECT 95.850 172.800 97.650 173.550 ;
        RECT 92.850 171.900 93.900 172.800 ;
        RECT 103.050 172.200 104.850 174.000 ;
        RECT 109.950 173.400 112.050 174.300 ;
        RECT 115.650 173.400 117.450 179.250 ;
        RECT 103.050 171.900 103.950 172.200 ;
        RECT 92.850 171.000 103.950 171.900 ;
        RECT 116.250 171.150 117.450 173.400 ;
        RECT 152.850 172.200 154.650 179.250 ;
        RECT 157.350 173.400 159.150 179.250 ;
        RECT 190.650 176.400 192.450 179.250 ;
        RECT 193.650 176.400 195.450 179.250 ;
        RECT 152.850 171.300 156.450 172.200 ;
        RECT 92.850 169.800 93.900 171.000 ;
        RECT 87.000 168.600 93.900 169.800 ;
        RECT 87.000 167.850 87.900 168.600 ;
        RECT 92.100 168.000 93.900 168.600 ;
        RECT 86.100 166.050 87.900 167.850 ;
        RECT 89.100 166.950 90.900 167.700 ;
        RECT 103.050 166.950 103.950 171.000 ;
        RECT 112.950 169.050 117.450 171.150 ;
        RECT 111.150 167.250 115.050 169.050 ;
        RECT 112.950 166.950 115.050 167.250 ;
        RECT 89.100 165.900 97.050 166.950 ;
        RECT 94.950 164.850 97.050 165.900 ;
        RECT 100.950 164.850 103.950 166.950 ;
        RECT 93.450 161.100 95.250 161.400 ;
        RECT 93.450 160.800 101.850 161.100 ;
        RECT 84.150 160.200 101.850 160.800 ;
        RECT 84.150 159.600 95.250 160.200 ;
        RECT 32.550 147.750 34.350 159.600 ;
        RECT 35.550 147.750 37.350 159.600 ;
        RECT 69.300 147.750 71.100 159.600 ;
        RECT 73.500 147.750 75.300 159.600 ;
        RECT 76.800 147.750 78.600 153.600 ;
        RECT 84.150 147.750 85.950 159.600 ;
        RECT 98.250 158.700 100.050 159.300 ;
        RECT 92.550 157.500 100.050 158.700 ;
        RECT 100.950 158.100 101.850 160.200 ;
        RECT 103.050 160.200 103.950 164.850 ;
        RECT 113.250 161.400 115.050 163.200 ;
        RECT 109.950 160.200 114.150 161.400 ;
        RECT 103.050 159.300 109.050 160.200 ;
        RECT 109.950 159.300 112.050 160.200 ;
        RECT 116.250 159.600 117.450 169.050 ;
        RECT 152.100 165.150 153.900 166.950 ;
        RECT 151.950 163.050 154.050 165.150 ;
        RECT 155.250 163.950 156.450 171.300 ;
        RECT 191.400 168.150 192.600 176.400 ;
        RECT 229.650 173.400 231.450 179.250 ;
        RECT 230.250 171.300 231.450 173.400 ;
        RECT 232.650 174.300 234.450 179.250 ;
        RECT 235.650 175.200 237.450 179.250 ;
        RECT 238.650 174.300 240.450 179.250 ;
        RECT 232.650 172.950 240.450 174.300 ;
        RECT 230.250 170.250 234.000 171.300 ;
        RECT 269.700 170.400 271.500 179.250 ;
        RECT 275.100 171.000 276.900 179.250 ;
        RECT 314.550 174.300 316.350 179.250 ;
        RECT 317.550 175.200 319.350 179.250 ;
        RECT 320.550 174.300 322.350 179.250 ;
        RECT 314.550 172.950 322.350 174.300 ;
        RECT 323.550 173.400 325.350 179.250 ;
        RECT 323.550 171.300 324.750 173.400 ;
        RECT 362.850 172.200 364.650 179.250 ;
        RECT 367.350 173.400 369.150 179.250 ;
        RECT 362.850 171.300 366.450 172.200 ;
        RECT 158.100 165.150 159.900 166.950 ;
        RECT 190.950 166.050 193.050 168.150 ;
        RECT 193.950 167.850 196.050 169.950 ;
        RECT 194.100 166.050 195.900 167.850 ;
        RECT 232.950 166.950 234.150 170.250 ;
        RECT 236.100 168.150 237.900 169.950 ;
        RECT 275.100 169.350 279.600 171.000 ;
        RECT 321.000 170.250 324.750 171.300 ;
        RECT 154.950 161.850 157.050 163.950 ;
        RECT 157.950 163.050 160.050 165.150 ;
        RECT 108.150 158.400 109.050 159.300 ;
        RECT 105.450 158.100 107.250 158.400 ;
        RECT 92.550 156.600 93.750 157.500 ;
        RECT 100.950 157.200 107.250 158.100 ;
        RECT 105.450 156.600 107.250 157.200 ;
        RECT 108.150 156.600 110.850 158.400 ;
        RECT 88.950 154.500 93.750 156.600 ;
        RECT 96.150 154.500 103.050 156.300 ;
        RECT 92.550 153.600 93.750 154.500 ;
        RECT 87.150 147.750 88.950 153.600 ;
        RECT 92.250 147.750 94.050 153.600 ;
        RECT 97.050 147.750 98.850 153.600 ;
        RECT 100.050 147.750 101.850 154.500 ;
        RECT 108.150 153.600 112.050 155.700 ;
        RECT 103.950 147.750 105.750 153.600 ;
        RECT 108.150 147.750 109.950 153.600 ;
        RECT 112.650 147.750 114.450 150.600 ;
        RECT 115.650 147.750 117.450 159.600 ;
        RECT 155.250 153.600 156.450 161.850 ;
        RECT 191.400 153.600 192.600 166.050 ;
        RECT 232.950 164.850 235.050 166.950 ;
        RECT 235.950 166.050 238.050 168.150 ;
        RECT 238.950 164.850 241.050 166.950 ;
        RECT 278.400 165.150 279.600 169.350 ;
        RECT 317.100 168.150 318.900 169.950 ;
        RECT 229.950 161.850 232.050 163.950 ;
        RECT 230.250 160.050 232.050 161.850 ;
        RECT 233.850 159.600 235.050 164.850 ;
        RECT 239.100 163.050 240.900 164.850 ;
        RECT 268.950 161.850 271.050 163.950 ;
        RECT 274.950 161.850 277.050 163.950 ;
        RECT 277.950 163.050 280.050 165.150 ;
        RECT 313.950 164.850 316.050 166.950 ;
        RECT 316.950 166.050 319.050 168.150 ;
        RECT 320.850 166.950 322.050 170.250 ;
        RECT 319.950 164.850 322.050 166.950 ;
        RECT 362.100 165.150 363.900 166.950 ;
        RECT 314.100 163.050 315.900 164.850 ;
        RECT 269.100 160.050 270.900 161.850 ;
        RECT 151.650 147.750 153.450 153.600 ;
        RECT 154.650 147.750 156.450 153.600 ;
        RECT 157.650 147.750 159.450 153.600 ;
        RECT 190.650 147.750 192.450 153.600 ;
        RECT 193.650 147.750 195.450 153.600 ;
        RECT 230.400 147.750 232.200 153.600 ;
        RECT 233.700 147.750 235.500 159.600 ;
        RECT 237.900 147.750 239.700 159.600 ;
        RECT 271.950 158.850 274.050 160.950 ;
        RECT 275.250 160.050 277.050 161.850 ;
        RECT 272.100 157.050 273.900 158.850 ;
        RECT 278.700 154.800 279.750 163.050 ;
        RECT 319.950 159.600 321.150 164.850 ;
        RECT 322.950 161.850 325.050 163.950 ;
        RECT 361.950 163.050 364.050 165.150 ;
        RECT 365.250 163.950 366.450 171.300 ;
        RECT 401.700 170.400 403.500 179.250 ;
        RECT 407.100 171.000 408.900 179.250 ;
        RECT 446.550 174.300 448.350 179.250 ;
        RECT 449.550 175.200 451.350 179.250 ;
        RECT 452.550 174.300 454.350 179.250 ;
        RECT 446.550 172.950 454.350 174.300 ;
        RECT 455.550 173.400 457.350 179.250 ;
        RECT 455.550 171.300 456.750 173.400 ;
        RECT 407.100 169.350 411.600 171.000 ;
        RECT 453.000 170.250 456.750 171.300 ;
        RECT 491.700 170.400 493.500 179.250 ;
        RECT 497.100 171.000 498.900 179.250 ;
        RECT 536.850 172.200 538.650 179.250 ;
        RECT 541.350 173.400 543.150 179.250 ;
        RECT 577.650 173.400 579.450 179.250 ;
        RECT 536.850 171.300 540.450 172.200 ;
        RECT 368.100 165.150 369.900 166.950 ;
        RECT 410.400 165.150 411.600 169.350 ;
        RECT 449.100 168.150 450.900 169.950 ;
        RECT 364.950 161.850 367.050 163.950 ;
        RECT 367.950 163.050 370.050 165.150 ;
        RECT 400.950 161.850 403.050 163.950 ;
        RECT 406.950 161.850 409.050 163.950 ;
        RECT 409.950 163.050 412.050 165.150 ;
        RECT 445.950 164.850 448.050 166.950 ;
        RECT 448.950 166.050 451.050 168.150 ;
        RECT 452.850 166.950 454.050 170.250 ;
        RECT 497.100 169.350 501.600 171.000 ;
        RECT 451.950 164.850 454.050 166.950 ;
        RECT 500.400 165.150 501.600 169.350 ;
        RECT 536.100 165.150 537.900 166.950 ;
        RECT 446.100 163.050 447.900 164.850 ;
        RECT 322.950 160.050 324.750 161.850 ;
        RECT 272.700 153.900 279.750 154.800 ;
        RECT 272.700 153.600 274.350 153.900 ;
        RECT 269.550 147.750 271.350 153.600 ;
        RECT 272.550 147.750 274.350 153.600 ;
        RECT 278.550 153.600 279.750 153.900 ;
        RECT 275.550 147.750 277.350 153.000 ;
        RECT 278.550 147.750 280.350 153.600 ;
        RECT 315.300 147.750 317.100 159.600 ;
        RECT 319.500 147.750 321.300 159.600 ;
        RECT 365.250 153.600 366.450 161.850 ;
        RECT 401.100 160.050 402.900 161.850 ;
        RECT 403.950 158.850 406.050 160.950 ;
        RECT 407.250 160.050 409.050 161.850 ;
        RECT 404.100 157.050 405.900 158.850 ;
        RECT 410.700 154.800 411.750 163.050 ;
        RECT 451.950 159.600 453.150 164.850 ;
        RECT 454.950 161.850 457.050 163.950 ;
        RECT 490.950 161.850 493.050 163.950 ;
        RECT 496.950 161.850 499.050 163.950 ;
        RECT 499.950 163.050 502.050 165.150 ;
        RECT 535.950 163.050 538.050 165.150 ;
        RECT 539.250 163.950 540.450 171.300 ;
        RECT 578.250 171.300 579.450 173.400 ;
        RECT 580.650 174.300 582.450 179.250 ;
        RECT 583.650 175.200 585.450 179.250 ;
        RECT 586.650 174.300 588.450 179.250 ;
        RECT 580.650 172.950 588.450 174.300 ;
        RECT 620.550 174.300 622.350 179.250 ;
        RECT 623.550 175.200 625.350 179.250 ;
        RECT 626.550 174.300 628.350 179.250 ;
        RECT 620.550 172.950 628.350 174.300 ;
        RECT 629.550 173.400 631.350 179.250 ;
        RECT 629.550 171.300 630.750 173.400 ;
        RECT 665.850 172.200 667.650 179.250 ;
        RECT 670.350 173.400 672.150 179.250 ;
        RECT 704.850 173.400 706.650 179.250 ;
        RECT 709.350 172.200 711.150 179.250 ;
        RECT 665.850 171.300 669.450 172.200 ;
        RECT 578.250 170.250 582.000 171.300 ;
        RECT 627.000 170.250 630.750 171.300 ;
        RECT 580.950 166.950 582.150 170.250 ;
        RECT 584.100 168.150 585.900 169.950 ;
        RECT 623.100 168.150 624.900 169.950 ;
        RECT 542.100 165.150 543.900 166.950 ;
        RECT 454.950 160.050 456.750 161.850 ;
        RECT 491.100 160.050 492.900 161.850 ;
        RECT 404.700 153.900 411.750 154.800 ;
        RECT 404.700 153.600 406.350 153.900 ;
        RECT 322.800 147.750 324.600 153.600 ;
        RECT 361.650 147.750 363.450 153.600 ;
        RECT 364.650 147.750 366.450 153.600 ;
        RECT 367.650 147.750 369.450 153.600 ;
        RECT 401.550 147.750 403.350 153.600 ;
        RECT 404.550 147.750 406.350 153.600 ;
        RECT 410.550 153.600 411.750 153.900 ;
        RECT 407.550 147.750 409.350 153.000 ;
        RECT 410.550 147.750 412.350 153.600 ;
        RECT 447.300 147.750 449.100 159.600 ;
        RECT 451.500 147.750 453.300 159.600 ;
        RECT 493.950 158.850 496.050 160.950 ;
        RECT 497.250 160.050 499.050 161.850 ;
        RECT 494.100 157.050 495.900 158.850 ;
        RECT 500.700 154.800 501.750 163.050 ;
        RECT 538.950 161.850 541.050 163.950 ;
        RECT 541.950 163.050 544.050 165.150 ;
        RECT 580.950 164.850 583.050 166.950 ;
        RECT 583.950 166.050 586.050 168.150 ;
        RECT 586.950 164.850 589.050 166.950 ;
        RECT 619.950 164.850 622.050 166.950 ;
        RECT 622.950 166.050 625.050 168.150 ;
        RECT 626.850 166.950 628.050 170.250 ;
        RECT 625.950 164.850 628.050 166.950 ;
        RECT 665.100 165.150 666.900 166.950 ;
        RECT 577.950 161.850 580.050 163.950 ;
        RECT 494.700 153.900 501.750 154.800 ;
        RECT 494.700 153.600 496.350 153.900 ;
        RECT 454.800 147.750 456.600 153.600 ;
        RECT 491.550 147.750 493.350 153.600 ;
        RECT 494.550 147.750 496.350 153.600 ;
        RECT 500.550 153.600 501.750 153.900 ;
        RECT 539.250 153.600 540.450 161.850 ;
        RECT 578.250 160.050 580.050 161.850 ;
        RECT 581.850 159.600 583.050 164.850 ;
        RECT 587.100 163.050 588.900 164.850 ;
        RECT 620.100 163.050 621.900 164.850 ;
        RECT 625.950 159.600 627.150 164.850 ;
        RECT 628.950 161.850 631.050 163.950 ;
        RECT 664.950 163.050 667.050 165.150 ;
        RECT 668.250 163.950 669.450 171.300 ;
        RECT 707.550 171.300 711.150 172.200 ;
        RECT 749.850 172.200 751.650 179.250 ;
        RECT 754.350 173.400 756.150 179.250 ;
        RECT 749.850 171.300 753.450 172.200 ;
        RECT 671.100 165.150 672.900 166.950 ;
        RECT 704.100 165.150 705.900 166.950 ;
        RECT 667.950 161.850 670.050 163.950 ;
        RECT 670.950 163.050 673.050 165.150 ;
        RECT 703.950 163.050 706.050 165.150 ;
        RECT 707.550 163.950 708.750 171.300 ;
        RECT 710.100 165.150 711.900 166.950 ;
        RECT 749.100 165.150 750.900 166.950 ;
        RECT 706.950 161.850 709.050 163.950 ;
        RECT 709.950 163.050 712.050 165.150 ;
        RECT 748.950 163.050 751.050 165.150 ;
        RECT 752.250 163.950 753.450 171.300 ;
        RECT 755.100 165.150 756.900 166.950 ;
        RECT 751.950 161.850 754.050 163.950 ;
        RECT 754.950 163.050 757.050 165.150 ;
        RECT 628.950 160.050 630.750 161.850 ;
        RECT 497.550 147.750 499.350 153.000 ;
        RECT 500.550 147.750 502.350 153.600 ;
        RECT 535.650 147.750 537.450 153.600 ;
        RECT 538.650 147.750 540.450 153.600 ;
        RECT 541.650 147.750 543.450 153.600 ;
        RECT 578.400 147.750 580.200 153.600 ;
        RECT 581.700 147.750 583.500 159.600 ;
        RECT 585.900 147.750 587.700 159.600 ;
        RECT 621.300 147.750 623.100 159.600 ;
        RECT 625.500 147.750 627.300 159.600 ;
        RECT 668.250 153.600 669.450 161.850 ;
        RECT 707.550 153.600 708.750 161.850 ;
        RECT 752.250 153.600 753.450 161.850 ;
        RECT 628.800 147.750 630.600 153.600 ;
        RECT 664.650 147.750 666.450 153.600 ;
        RECT 667.650 147.750 669.450 153.600 ;
        RECT 670.650 147.750 672.450 153.600 ;
        RECT 704.550 147.750 706.350 153.600 ;
        RECT 707.550 147.750 709.350 153.600 ;
        RECT 710.550 147.750 712.350 153.600 ;
        RECT 748.650 147.750 750.450 153.600 ;
        RECT 751.650 147.750 753.450 153.600 ;
        RECT 754.650 147.750 756.450 153.600 ;
        RECT 2.550 131.400 4.350 143.250 ;
        RECT 5.550 140.400 7.350 143.250 ;
        RECT 10.050 137.400 11.850 143.250 ;
        RECT 14.250 137.400 16.050 143.250 ;
        RECT 7.950 135.300 11.850 137.400 ;
        RECT 18.150 136.500 19.950 143.250 ;
        RECT 21.150 137.400 22.950 143.250 ;
        RECT 25.950 137.400 27.750 143.250 ;
        RECT 31.050 137.400 32.850 143.250 ;
        RECT 26.250 136.500 27.450 137.400 ;
        RECT 16.950 134.700 23.850 136.500 ;
        RECT 26.250 134.400 31.050 136.500 ;
        RECT 9.150 132.600 11.850 134.400 ;
        RECT 12.750 133.800 14.550 134.400 ;
        RECT 12.750 132.900 19.050 133.800 ;
        RECT 26.250 133.500 27.450 134.400 ;
        RECT 12.750 132.600 14.550 132.900 ;
        RECT 10.950 131.700 11.850 132.600 ;
        RECT 2.550 121.950 3.750 131.400 ;
        RECT 7.950 130.800 10.050 131.700 ;
        RECT 10.950 130.800 16.950 131.700 ;
        RECT 5.850 129.600 10.050 130.800 ;
        RECT 4.950 127.800 6.750 129.600 ;
        RECT 16.050 126.150 16.950 130.800 ;
        RECT 18.150 130.800 19.050 132.900 ;
        RECT 19.950 132.300 27.450 133.500 ;
        RECT 19.950 131.700 21.750 132.300 ;
        RECT 34.050 131.400 35.850 143.250 ;
        RECT 70.650 131.400 72.450 143.250 ;
        RECT 24.750 130.800 35.850 131.400 ;
        RECT 18.150 130.200 35.850 130.800 ;
        RECT 73.650 130.500 75.450 143.250 ;
        RECT 76.650 131.400 78.450 143.250 ;
        RECT 79.650 130.500 81.450 143.250 ;
        RECT 82.650 131.400 84.450 143.250 ;
        RECT 85.650 130.500 87.450 143.250 ;
        RECT 88.650 131.400 90.450 143.250 ;
        RECT 91.650 130.500 93.450 143.250 ;
        RECT 94.650 131.400 96.450 143.250 ;
        RECT 99.150 131.400 100.950 143.250 ;
        RECT 102.150 137.400 103.950 143.250 ;
        RECT 107.250 137.400 109.050 143.250 ;
        RECT 112.050 137.400 113.850 143.250 ;
        RECT 107.550 136.500 108.750 137.400 ;
        RECT 115.050 136.500 116.850 143.250 ;
        RECT 118.950 137.400 120.750 143.250 ;
        RECT 123.150 137.400 124.950 143.250 ;
        RECT 127.650 140.400 129.450 143.250 ;
        RECT 103.950 134.400 108.750 136.500 ;
        RECT 111.150 134.700 118.050 136.500 ;
        RECT 123.150 135.300 127.050 137.400 ;
        RECT 107.550 133.500 108.750 134.400 ;
        RECT 120.450 133.800 122.250 134.400 ;
        RECT 107.550 132.300 115.050 133.500 ;
        RECT 113.250 131.700 115.050 132.300 ;
        RECT 115.950 132.900 122.250 133.800 ;
        RECT 18.150 129.900 26.550 130.200 ;
        RECT 24.750 129.600 26.550 129.900 ;
        RECT 16.050 124.050 19.050 126.150 ;
        RECT 22.950 125.100 25.050 126.150 ;
        RECT 22.950 124.050 30.900 125.100 ;
        RECT 4.950 123.750 7.050 124.050 ;
        RECT 4.950 121.950 8.850 123.750 ;
        RECT 2.550 119.850 7.050 121.950 ;
        RECT 16.050 120.000 16.950 124.050 ;
        RECT 29.100 123.300 30.900 124.050 ;
        RECT 32.100 123.150 33.900 124.950 ;
        RECT 26.100 122.400 27.900 123.000 ;
        RECT 32.100 122.400 33.000 123.150 ;
        RECT 26.100 121.200 33.000 122.400 ;
        RECT 26.100 120.000 27.150 121.200 ;
        RECT 2.550 117.600 3.750 119.850 ;
        RECT 16.050 119.100 27.150 120.000 ;
        RECT 16.050 118.800 16.950 119.100 ;
        RECT 2.550 111.750 4.350 117.600 ;
        RECT 7.950 116.700 10.050 117.600 ;
        RECT 15.150 117.000 16.950 118.800 ;
        RECT 26.100 118.200 27.150 119.100 ;
        RECT 22.350 117.450 24.150 118.200 ;
        RECT 7.950 115.500 11.700 116.700 ;
        RECT 10.650 114.600 11.700 115.500 ;
        RECT 19.200 116.400 24.150 117.450 ;
        RECT 25.650 116.400 27.450 118.200 ;
        RECT 34.950 117.600 35.850 130.200 ;
        RECT 72.750 129.300 75.450 130.500 ;
        RECT 77.700 129.300 81.450 130.500 ;
        RECT 83.700 129.300 87.450 130.500 ;
        RECT 89.550 129.300 93.450 130.500 ;
        RECT 99.150 130.800 110.250 131.400 ;
        RECT 115.950 130.800 116.850 132.900 ;
        RECT 120.450 132.600 122.250 132.900 ;
        RECT 123.150 132.600 125.850 134.400 ;
        RECT 123.150 131.700 124.050 132.600 ;
        RECT 99.150 130.200 116.850 130.800 ;
        RECT 72.750 124.950 73.800 129.300 ;
        RECT 70.950 122.850 73.800 124.950 ;
        RECT 72.750 119.700 73.800 122.850 ;
        RECT 77.700 122.400 78.900 129.300 ;
        RECT 83.700 122.400 84.900 129.300 ;
        RECT 89.550 122.400 90.750 129.300 ;
        RECT 91.950 122.850 94.050 124.950 ;
        RECT 74.700 120.600 78.900 122.400 ;
        RECT 80.700 120.600 84.900 122.400 ;
        RECT 86.700 120.600 90.750 122.400 ;
        RECT 92.100 121.050 93.900 122.850 ;
        RECT 77.700 119.700 78.900 120.600 ;
        RECT 83.700 119.700 84.900 120.600 ;
        RECT 89.550 119.700 90.750 120.600 ;
        RECT 72.750 118.650 75.600 119.700 ;
        RECT 72.900 118.500 75.600 118.650 ;
        RECT 77.700 118.500 81.600 119.700 ;
        RECT 83.700 118.500 87.450 119.700 ;
        RECT 89.550 118.500 93.600 119.700 ;
        RECT 73.800 117.600 75.600 118.500 ;
        RECT 79.800 117.600 81.600 118.500 ;
        RECT 19.200 114.600 20.250 116.400 ;
        RECT 28.950 115.500 31.050 117.600 ;
        RECT 28.950 114.600 30.000 115.500 ;
        RECT 5.850 111.750 7.650 114.600 ;
        RECT 10.350 111.750 12.150 114.600 ;
        RECT 14.550 111.750 16.350 114.600 ;
        RECT 18.450 111.750 20.250 114.600 ;
        RECT 21.750 111.750 23.550 114.600 ;
        RECT 26.250 113.700 30.000 114.600 ;
        RECT 26.250 111.750 28.050 113.700 ;
        RECT 31.050 111.750 32.850 114.600 ;
        RECT 34.050 111.750 35.850 117.600 ;
        RECT 70.650 111.750 72.450 117.600 ;
        RECT 73.650 111.750 75.450 117.600 ;
        RECT 76.650 111.750 78.450 117.600 ;
        RECT 79.650 111.750 81.450 117.600 ;
        RECT 82.650 111.750 84.450 117.600 ;
        RECT 85.650 111.750 87.450 118.500 ;
        RECT 91.800 117.600 93.600 118.500 ;
        RECT 99.150 117.600 100.050 130.200 ;
        RECT 108.450 129.900 116.850 130.200 ;
        RECT 118.050 130.800 124.050 131.700 ;
        RECT 124.950 130.800 127.050 131.700 ;
        RECT 130.650 131.400 132.450 143.250 ;
        RECT 165.300 131.400 167.100 143.250 ;
        RECT 169.500 131.400 171.300 143.250 ;
        RECT 172.800 137.400 174.600 143.250 ;
        RECT 209.550 137.400 211.350 143.250 ;
        RECT 212.550 137.400 214.350 143.250 ;
        RECT 215.550 137.400 217.350 143.250 ;
        RECT 108.450 129.600 110.250 129.900 ;
        RECT 118.050 126.150 118.950 130.800 ;
        RECT 124.950 129.600 129.150 130.800 ;
        RECT 128.250 127.800 130.050 129.600 ;
        RECT 109.950 125.100 112.050 126.150 ;
        RECT 101.100 123.150 102.900 124.950 ;
        RECT 104.100 124.050 112.050 125.100 ;
        RECT 115.950 124.050 118.950 126.150 ;
        RECT 104.100 123.300 105.900 124.050 ;
        RECT 102.000 122.400 102.900 123.150 ;
        RECT 107.100 122.400 108.900 123.000 ;
        RECT 102.000 121.200 108.900 122.400 ;
        RECT 107.850 120.000 108.900 121.200 ;
        RECT 118.050 120.000 118.950 124.050 ;
        RECT 127.950 123.750 130.050 124.050 ;
        RECT 126.150 121.950 130.050 123.750 ;
        RECT 131.250 121.950 132.450 131.400 ;
        RECT 164.100 126.150 165.900 127.950 ;
        RECT 169.950 126.150 171.150 131.400 ;
        RECT 172.950 129.150 174.750 130.950 ;
        RECT 212.550 129.150 213.750 137.400 ;
        RECT 251.550 131.400 253.350 143.250 ;
        RECT 255.750 131.400 257.550 143.250 ;
        RECT 293.550 137.400 295.350 143.250 ;
        RECT 296.550 137.400 298.350 143.250 ;
        RECT 299.550 138.000 301.350 143.250 ;
        RECT 296.700 137.100 298.350 137.400 ;
        RECT 302.550 137.400 304.350 143.250 ;
        RECT 338.550 137.400 340.350 143.250 ;
        RECT 341.550 137.400 343.350 143.250 ;
        RECT 344.550 137.400 346.350 143.250 ;
        RECT 380.550 137.400 382.350 143.250 ;
        RECT 383.550 137.400 385.350 143.250 ;
        RECT 386.550 137.400 388.350 143.250 ;
        RECT 422.550 137.400 424.350 143.250 ;
        RECT 425.550 137.400 427.350 143.250 ;
        RECT 428.550 138.000 430.350 143.250 ;
        RECT 302.550 137.100 303.750 137.400 ;
        RECT 296.700 136.200 303.750 137.100 ;
        RECT 296.100 132.150 297.900 133.950 ;
        RECT 255.000 130.350 257.550 131.400 ;
        RECT 172.950 127.050 175.050 129.150 ;
        RECT 163.950 124.050 166.050 126.150 ;
        RECT 166.950 122.850 169.050 124.950 ;
        RECT 169.950 124.050 172.050 126.150 ;
        RECT 208.950 125.850 211.050 127.950 ;
        RECT 211.950 127.050 214.050 129.150 ;
        RECT 209.100 124.050 210.900 125.850 ;
        RECT 107.850 119.100 118.950 120.000 ;
        RECT 127.950 119.850 132.450 121.950 ;
        RECT 167.100 121.050 168.900 122.850 ;
        RECT 170.850 120.750 172.050 124.050 ;
        RECT 107.850 118.200 108.900 119.100 ;
        RECT 118.050 118.800 118.950 119.100 ;
        RECT 88.650 111.750 90.450 117.600 ;
        RECT 91.650 111.750 93.450 117.600 ;
        RECT 94.650 111.750 96.450 117.600 ;
        RECT 99.150 111.750 100.950 117.600 ;
        RECT 103.950 115.500 106.050 117.600 ;
        RECT 107.550 116.400 109.350 118.200 ;
        RECT 110.850 117.450 112.650 118.200 ;
        RECT 110.850 116.400 115.800 117.450 ;
        RECT 118.050 117.000 119.850 118.800 ;
        RECT 131.250 117.600 132.450 119.850 ;
        RECT 171.000 119.700 174.750 120.750 ;
        RECT 124.950 116.700 127.050 117.600 ;
        RECT 105.000 114.600 106.050 115.500 ;
        RECT 114.750 114.600 115.800 116.400 ;
        RECT 123.300 115.500 127.050 116.700 ;
        RECT 123.300 114.600 124.350 115.500 ;
        RECT 102.150 111.750 103.950 114.600 ;
        RECT 105.000 113.700 108.750 114.600 ;
        RECT 106.950 111.750 108.750 113.700 ;
        RECT 111.450 111.750 113.250 114.600 ;
        RECT 114.750 111.750 116.550 114.600 ;
        RECT 118.650 111.750 120.450 114.600 ;
        RECT 122.850 111.750 124.650 114.600 ;
        RECT 127.350 111.750 129.150 114.600 ;
        RECT 130.650 111.750 132.450 117.600 ;
        RECT 164.550 116.700 172.350 118.050 ;
        RECT 164.550 111.750 166.350 116.700 ;
        RECT 167.550 111.750 169.350 115.800 ;
        RECT 170.550 111.750 172.350 116.700 ;
        RECT 173.550 117.600 174.750 119.700 ;
        RECT 212.550 119.700 213.750 127.050 ;
        RECT 214.950 125.850 217.050 127.950 ;
        RECT 251.100 126.150 252.900 127.950 ;
        RECT 215.100 124.050 216.900 125.850 ;
        RECT 250.950 124.050 253.050 126.150 ;
        RECT 255.000 123.150 256.050 130.350 ;
        RECT 293.100 129.150 294.900 130.950 ;
        RECT 295.950 130.050 298.050 132.150 ;
        RECT 299.250 129.150 301.050 130.950 ;
        RECT 257.100 126.150 258.900 127.950 ;
        RECT 292.950 127.050 295.050 129.150 ;
        RECT 298.950 127.050 301.050 129.150 ;
        RECT 302.700 127.950 303.750 136.200 ;
        RECT 341.550 129.150 342.750 137.400 ;
        RECT 383.550 129.150 384.750 137.400 ;
        RECT 425.700 137.100 427.350 137.400 ;
        RECT 431.550 137.400 433.350 143.250 ;
        RECT 466.650 137.400 468.450 143.250 ;
        RECT 469.650 138.000 471.450 143.250 ;
        RECT 431.550 137.100 432.750 137.400 ;
        RECT 425.700 136.200 432.750 137.100 ;
        RECT 425.100 132.150 426.900 133.950 ;
        RECT 422.100 129.150 423.900 130.950 ;
        RECT 424.950 130.050 427.050 132.150 ;
        RECT 428.250 129.150 430.050 130.950 ;
        RECT 256.950 124.050 259.050 126.150 ;
        RECT 301.950 125.850 304.050 127.950 ;
        RECT 337.950 125.850 340.050 127.950 ;
        RECT 340.950 127.050 343.050 129.150 ;
        RECT 253.950 121.050 256.050 123.150 ;
        RECT 302.400 121.650 303.600 125.850 ;
        RECT 338.100 124.050 339.900 125.850 ;
        RECT 212.550 118.800 216.150 119.700 ;
        RECT 173.550 111.750 175.350 117.600 ;
        RECT 209.850 111.750 211.650 117.600 ;
        RECT 214.350 111.750 216.150 118.800 ;
        RECT 255.000 114.600 256.050 121.050 ;
        RECT 251.550 111.750 253.350 114.600 ;
        RECT 254.550 111.750 256.350 114.600 ;
        RECT 257.550 111.750 259.350 114.600 ;
        RECT 293.700 111.750 295.500 120.600 ;
        RECT 299.100 120.000 303.600 121.650 ;
        RECT 299.100 111.750 300.900 120.000 ;
        RECT 341.550 119.700 342.750 127.050 ;
        RECT 343.950 125.850 346.050 127.950 ;
        RECT 379.950 125.850 382.050 127.950 ;
        RECT 382.950 127.050 385.050 129.150 ;
        RECT 344.100 124.050 345.900 125.850 ;
        RECT 380.100 124.050 381.900 125.850 ;
        RECT 383.550 119.700 384.750 127.050 ;
        RECT 385.950 125.850 388.050 127.950 ;
        RECT 421.950 127.050 424.050 129.150 ;
        RECT 427.950 127.050 430.050 129.150 ;
        RECT 431.700 127.950 432.750 136.200 ;
        RECT 467.250 137.100 468.450 137.400 ;
        RECT 472.650 137.400 474.450 143.250 ;
        RECT 475.650 137.400 477.450 143.250 ;
        RECT 472.650 137.100 474.300 137.400 ;
        RECT 467.250 136.200 474.300 137.100 ;
        RECT 467.250 127.950 468.300 136.200 ;
        RECT 473.100 132.150 474.900 133.950 ;
        RECT 469.950 129.150 471.750 130.950 ;
        RECT 472.950 130.050 475.050 132.150 ;
        RECT 510.300 131.400 512.100 143.250 ;
        RECT 514.500 131.400 516.300 143.250 ;
        RECT 517.800 137.400 519.600 143.250 ;
        RECT 551.550 137.400 553.350 143.250 ;
        RECT 554.550 137.400 556.350 143.250 ;
        RECT 590.550 137.400 592.350 143.250 ;
        RECT 593.550 137.400 595.350 143.250 ;
        RECT 596.550 137.400 598.350 143.250 ;
        RECT 476.100 129.150 477.900 130.950 ;
        RECT 430.950 125.850 433.050 127.950 ;
        RECT 466.950 125.850 469.050 127.950 ;
        RECT 469.950 127.050 472.050 129.150 ;
        RECT 475.950 127.050 478.050 129.150 ;
        RECT 509.100 126.150 510.900 127.950 ;
        RECT 514.950 126.150 516.150 131.400 ;
        RECT 517.950 129.150 519.750 130.950 ;
        RECT 517.950 127.050 520.050 129.150 ;
        RECT 386.100 124.050 387.900 125.850 ;
        RECT 431.400 121.650 432.600 125.850 ;
        RECT 341.550 118.800 345.150 119.700 ;
        RECT 383.550 118.800 387.150 119.700 ;
        RECT 338.850 111.750 340.650 117.600 ;
        RECT 343.350 111.750 345.150 118.800 ;
        RECT 380.850 111.750 382.650 117.600 ;
        RECT 385.350 111.750 387.150 118.800 ;
        RECT 422.700 111.750 424.500 120.600 ;
        RECT 428.100 120.000 432.600 121.650 ;
        RECT 467.400 121.650 468.600 125.850 ;
        RECT 508.950 124.050 511.050 126.150 ;
        RECT 511.950 122.850 514.050 124.950 ;
        RECT 514.950 124.050 517.050 126.150 ;
        RECT 554.400 124.950 555.600 137.400 ;
        RECT 593.550 129.150 594.750 137.400 ;
        RECT 629.550 131.400 631.350 143.250 ;
        RECT 634.050 131.550 635.850 143.250 ;
        RECT 637.050 132.900 638.850 143.250 ;
        RECT 674.550 137.400 676.350 143.250 ;
        RECT 677.550 137.400 679.350 143.250 ;
        RECT 680.550 137.400 682.350 143.250 ;
        RECT 718.650 137.400 720.450 143.250 ;
        RECT 721.650 137.400 723.450 143.250 ;
        RECT 724.650 137.400 726.450 143.250 ;
        RECT 637.050 131.550 639.450 132.900 ;
        RECT 629.550 130.200 630.750 131.400 ;
        RECT 634.950 130.200 636.750 130.650 ;
        RECT 589.950 125.850 592.050 127.950 ;
        RECT 592.950 127.050 595.050 129.150 ;
        RECT 629.550 129.000 636.750 130.200 ;
        RECT 634.950 128.850 636.750 129.000 ;
        RECT 467.400 120.000 471.900 121.650 ;
        RECT 512.100 121.050 513.900 122.850 ;
        RECT 515.850 120.750 517.050 124.050 ;
        RECT 551.100 123.150 552.900 124.950 ;
        RECT 550.950 121.050 553.050 123.150 ;
        RECT 553.950 122.850 556.050 124.950 ;
        RECT 590.100 124.050 591.900 125.850 ;
        RECT 428.100 111.750 429.900 120.000 ;
        RECT 470.100 111.750 471.900 120.000 ;
        RECT 475.500 111.750 477.300 120.600 ;
        RECT 516.000 119.700 519.750 120.750 ;
        RECT 509.550 116.700 517.350 118.050 ;
        RECT 509.550 111.750 511.350 116.700 ;
        RECT 512.550 111.750 514.350 115.800 ;
        RECT 515.550 111.750 517.350 116.700 ;
        RECT 518.550 117.600 519.750 119.700 ;
        RECT 518.550 111.750 520.350 117.600 ;
        RECT 554.400 114.600 555.600 122.850 ;
        RECT 593.550 119.700 594.750 127.050 ;
        RECT 595.950 125.850 598.050 127.950 ;
        RECT 632.100 126.150 633.900 127.950 ;
        RECT 596.100 124.050 597.900 125.850 ;
        RECT 629.100 123.150 630.900 124.950 ;
        RECT 631.950 124.050 634.050 126.150 ;
        RECT 628.950 121.050 631.050 123.150 ;
        RECT 635.700 120.600 636.600 128.850 ;
        RECT 638.100 124.950 639.450 131.550 ;
        RECT 677.550 129.150 678.750 137.400 ;
        RECT 722.250 129.150 723.450 137.400 ;
        RECT 673.950 125.850 676.050 127.950 ;
        RECT 676.950 127.050 679.050 129.150 ;
        RECT 637.950 122.850 640.050 124.950 ;
        RECT 674.100 124.050 675.900 125.850 ;
        RECT 634.950 119.700 636.750 120.600 ;
        RECT 593.550 118.800 597.150 119.700 ;
        RECT 551.550 111.750 553.350 114.600 ;
        RECT 554.550 111.750 556.350 114.600 ;
        RECT 590.850 111.750 592.650 117.600 ;
        RECT 595.350 111.750 597.150 118.800 ;
        RECT 633.450 118.800 636.750 119.700 ;
        RECT 633.450 114.600 634.350 118.800 ;
        RECT 639.000 117.600 640.050 122.850 ;
        RECT 677.550 119.700 678.750 127.050 ;
        RECT 679.950 125.850 682.050 127.950 ;
        RECT 718.950 125.850 721.050 127.950 ;
        RECT 721.950 127.050 724.050 129.150 ;
        RECT 680.100 124.050 681.900 125.850 ;
        RECT 719.100 124.050 720.900 125.850 ;
        RECT 722.250 119.700 723.450 127.050 ;
        RECT 724.950 125.850 727.050 127.950 ;
        RECT 725.100 124.050 726.900 125.850 ;
        RECT 677.550 118.800 681.150 119.700 ;
        RECT 629.550 111.750 631.350 114.600 ;
        RECT 632.550 111.750 634.350 114.600 ;
        RECT 635.550 111.750 637.350 114.600 ;
        RECT 638.550 111.750 640.350 117.600 ;
        RECT 674.850 111.750 676.650 117.600 ;
        RECT 679.350 111.750 681.150 118.800 ;
        RECT 719.850 118.800 723.450 119.700 ;
        RECT 719.850 111.750 721.650 118.800 ;
        RECT 724.350 111.750 726.150 117.600 ;
        RECT 34.650 104.400 36.450 107.250 ;
        RECT 37.650 104.400 39.450 107.250 ;
        RECT 40.650 104.400 42.450 107.250 ;
        RECT 37.950 97.950 39.000 104.400 ;
        RECT 77.850 100.200 79.650 107.250 ;
        RECT 82.350 101.400 84.150 107.250 ;
        RECT 116.550 102.300 118.350 107.250 ;
        RECT 119.550 103.200 121.350 107.250 ;
        RECT 122.550 102.300 124.350 107.250 ;
        RECT 116.550 100.950 124.350 102.300 ;
        RECT 125.550 101.400 127.350 107.250 ;
        RECT 132.150 101.400 133.950 107.250 ;
        RECT 135.150 104.400 136.950 107.250 ;
        RECT 139.950 105.300 141.750 107.250 ;
        RECT 138.000 104.400 141.750 105.300 ;
        RECT 144.450 104.400 146.250 107.250 ;
        RECT 147.750 104.400 149.550 107.250 ;
        RECT 151.650 104.400 153.450 107.250 ;
        RECT 155.850 104.400 157.650 107.250 ;
        RECT 160.350 104.400 162.150 107.250 ;
        RECT 138.000 103.500 139.050 104.400 ;
        RECT 136.950 101.400 139.050 103.500 ;
        RECT 147.750 102.600 148.800 104.400 ;
        RECT 77.850 99.300 81.450 100.200 ;
        RECT 125.550 99.300 126.750 101.400 ;
        RECT 37.950 95.850 40.050 97.950 ;
        RECT 34.950 92.850 37.050 94.950 ;
        RECT 35.100 91.050 36.900 92.850 ;
        RECT 37.950 88.650 39.000 95.850 ;
        RECT 40.950 92.850 43.050 94.950 ;
        RECT 77.100 93.150 78.900 94.950 ;
        RECT 41.100 91.050 42.900 92.850 ;
        RECT 76.950 91.050 79.050 93.150 ;
        RECT 80.250 91.950 81.450 99.300 ;
        RECT 123.000 98.250 126.750 99.300 ;
        RECT 119.100 96.150 120.900 97.950 ;
        RECT 83.100 93.150 84.900 94.950 ;
        RECT 79.950 89.850 82.050 91.950 ;
        RECT 82.950 91.050 85.050 93.150 ;
        RECT 115.950 92.850 118.050 94.950 ;
        RECT 118.950 94.050 121.050 96.150 ;
        RECT 122.850 94.950 124.050 98.250 ;
        RECT 121.950 92.850 124.050 94.950 ;
        RECT 116.100 91.050 117.900 92.850 ;
        RECT 36.450 87.600 39.000 88.650 ;
        RECT 36.450 75.750 38.250 87.600 ;
        RECT 40.650 75.750 42.450 87.600 ;
        RECT 80.250 81.600 81.450 89.850 ;
        RECT 121.950 87.600 123.150 92.850 ;
        RECT 124.950 89.850 127.050 91.950 ;
        RECT 124.950 88.050 126.750 89.850 ;
        RECT 132.150 88.800 133.050 101.400 ;
        RECT 140.550 100.800 142.350 102.600 ;
        RECT 143.850 101.550 148.800 102.600 ;
        RECT 156.300 103.500 157.350 104.400 ;
        RECT 156.300 102.300 160.050 103.500 ;
        RECT 143.850 100.800 145.650 101.550 ;
        RECT 140.850 99.900 141.900 100.800 ;
        RECT 151.050 100.200 152.850 102.000 ;
        RECT 157.950 101.400 160.050 102.300 ;
        RECT 163.650 101.400 165.450 107.250 ;
        RECT 151.050 99.900 151.950 100.200 ;
        RECT 140.850 99.000 151.950 99.900 ;
        RECT 164.250 99.150 165.450 101.400 ;
        RECT 140.850 97.800 141.900 99.000 ;
        RECT 135.000 96.600 141.900 97.800 ;
        RECT 135.000 95.850 135.900 96.600 ;
        RECT 140.100 96.000 141.900 96.600 ;
        RECT 134.100 94.050 135.900 95.850 ;
        RECT 137.100 94.950 138.900 95.700 ;
        RECT 151.050 94.950 151.950 99.000 ;
        RECT 160.950 97.050 165.450 99.150 ;
        RECT 159.150 95.250 163.050 97.050 ;
        RECT 160.950 94.950 163.050 95.250 ;
        RECT 137.100 93.900 145.050 94.950 ;
        RECT 142.950 92.850 145.050 93.900 ;
        RECT 148.950 92.850 151.950 94.950 ;
        RECT 141.450 89.100 143.250 89.400 ;
        RECT 141.450 88.800 149.850 89.100 ;
        RECT 132.150 88.200 149.850 88.800 ;
        RECT 132.150 87.600 143.250 88.200 ;
        RECT 76.650 75.750 78.450 81.600 ;
        RECT 79.650 75.750 81.450 81.600 ;
        RECT 82.650 75.750 84.450 81.600 ;
        RECT 117.300 75.750 119.100 87.600 ;
        RECT 121.500 75.750 123.300 87.600 ;
        RECT 124.800 75.750 126.600 81.600 ;
        RECT 132.150 75.750 133.950 87.600 ;
        RECT 146.250 86.700 148.050 87.300 ;
        RECT 140.550 85.500 148.050 86.700 ;
        RECT 148.950 86.100 149.850 88.200 ;
        RECT 151.050 88.200 151.950 92.850 ;
        RECT 161.250 89.400 163.050 91.200 ;
        RECT 157.950 88.200 162.150 89.400 ;
        RECT 151.050 87.300 157.050 88.200 ;
        RECT 157.950 87.300 160.050 88.200 ;
        RECT 164.250 87.600 165.450 97.050 ;
        RECT 156.150 86.400 157.050 87.300 ;
        RECT 153.450 86.100 155.250 86.400 ;
        RECT 140.550 84.600 141.750 85.500 ;
        RECT 148.950 85.200 155.250 86.100 ;
        RECT 153.450 84.600 155.250 85.200 ;
        RECT 156.150 84.600 158.850 86.400 ;
        RECT 136.950 82.500 141.750 84.600 ;
        RECT 144.150 82.500 151.050 84.300 ;
        RECT 140.550 81.600 141.750 82.500 ;
        RECT 135.150 75.750 136.950 81.600 ;
        RECT 140.250 75.750 142.050 81.600 ;
        RECT 145.050 75.750 146.850 81.600 ;
        RECT 148.050 75.750 149.850 82.500 ;
        RECT 156.150 81.600 160.050 83.700 ;
        RECT 151.950 75.750 153.750 81.600 ;
        RECT 156.150 75.750 157.950 81.600 ;
        RECT 160.650 75.750 162.450 78.600 ;
        RECT 163.650 75.750 165.450 87.600 ;
        RECT 167.550 101.400 169.350 107.250 ;
        RECT 170.850 104.400 172.650 107.250 ;
        RECT 175.350 104.400 177.150 107.250 ;
        RECT 179.550 104.400 181.350 107.250 ;
        RECT 183.450 104.400 185.250 107.250 ;
        RECT 186.750 104.400 188.550 107.250 ;
        RECT 191.250 105.300 193.050 107.250 ;
        RECT 191.250 104.400 195.000 105.300 ;
        RECT 196.050 104.400 197.850 107.250 ;
        RECT 175.650 103.500 176.700 104.400 ;
        RECT 172.950 102.300 176.700 103.500 ;
        RECT 184.200 102.600 185.250 104.400 ;
        RECT 193.950 103.500 195.000 104.400 ;
        RECT 172.950 101.400 175.050 102.300 ;
        RECT 167.550 99.150 168.750 101.400 ;
        RECT 180.150 100.200 181.950 102.000 ;
        RECT 184.200 101.550 189.150 102.600 ;
        RECT 187.350 100.800 189.150 101.550 ;
        RECT 190.650 100.800 192.450 102.600 ;
        RECT 193.950 101.400 196.050 103.500 ;
        RECT 199.050 101.400 200.850 107.250 ;
        RECT 230.550 104.400 232.350 107.250 ;
        RECT 233.550 104.400 235.350 107.250 ;
        RECT 236.550 104.400 238.350 107.250 ;
        RECT 181.050 99.900 181.950 100.200 ;
        RECT 191.100 99.900 192.150 100.800 ;
        RECT 167.550 97.050 172.050 99.150 ;
        RECT 181.050 99.000 192.150 99.900 ;
        RECT 167.550 87.600 168.750 97.050 ;
        RECT 169.950 95.250 173.850 97.050 ;
        RECT 169.950 94.950 172.050 95.250 ;
        RECT 181.050 94.950 181.950 99.000 ;
        RECT 191.100 97.800 192.150 99.000 ;
        RECT 191.100 96.600 198.000 97.800 ;
        RECT 191.100 96.000 192.900 96.600 ;
        RECT 197.100 95.850 198.000 96.600 ;
        RECT 194.100 94.950 195.900 95.700 ;
        RECT 181.050 92.850 184.050 94.950 ;
        RECT 187.950 93.900 195.900 94.950 ;
        RECT 197.100 94.050 198.900 95.850 ;
        RECT 187.950 92.850 190.050 93.900 ;
        RECT 169.950 89.400 171.750 91.200 ;
        RECT 170.850 88.200 175.050 89.400 ;
        RECT 181.050 88.200 181.950 92.850 ;
        RECT 189.750 89.100 191.550 89.400 ;
        RECT 167.550 75.750 169.350 87.600 ;
        RECT 172.950 87.300 175.050 88.200 ;
        RECT 175.950 87.300 181.950 88.200 ;
        RECT 183.150 88.800 191.550 89.100 ;
        RECT 199.950 88.800 200.850 101.400 ;
        RECT 217.950 99.450 220.050 100.050 ;
        RECT 229.950 99.450 232.050 100.050 ;
        RECT 217.950 98.550 232.050 99.450 ;
        RECT 217.950 97.950 220.050 98.550 ;
        RECT 229.950 97.950 232.050 98.550 ;
        RECT 234.000 97.950 235.050 104.400 ;
        RECT 273.150 102.900 274.950 107.250 ;
        RECT 232.950 95.850 235.050 97.950 ;
        RECT 229.950 92.850 232.050 94.950 ;
        RECT 230.100 91.050 231.900 92.850 ;
        RECT 183.150 88.200 200.850 88.800 ;
        RECT 175.950 86.400 176.850 87.300 ;
        RECT 174.150 84.600 176.850 86.400 ;
        RECT 177.750 86.100 179.550 86.400 ;
        RECT 183.150 86.100 184.050 88.200 ;
        RECT 189.750 87.600 200.850 88.200 ;
        RECT 234.000 88.650 235.050 95.850 ;
        RECT 271.650 101.400 274.950 102.900 ;
        RECT 276.150 101.400 277.950 107.250 ;
        RECT 271.650 94.950 272.850 101.400 ;
        RECT 274.950 99.900 276.750 100.500 ;
        RECT 280.650 99.900 282.450 107.250 ;
        RECT 314.850 101.400 316.650 107.250 ;
        RECT 319.350 100.200 321.150 107.250 ;
        RECT 356.850 101.400 358.650 107.250 ;
        RECT 361.350 100.200 363.150 107.250 ;
        RECT 274.950 98.700 282.450 99.900 ;
        RECT 317.550 99.300 321.150 100.200 ;
        RECT 359.550 99.300 363.150 100.200 ;
        RECT 235.950 92.850 238.050 94.950 ;
        RECT 271.650 92.850 274.050 94.950 ;
        RECT 275.100 93.150 276.900 94.950 ;
        RECT 236.100 91.050 237.900 92.850 ;
        RECT 234.000 87.600 236.550 88.650 ;
        RECT 271.650 87.600 272.850 92.850 ;
        RECT 274.950 91.050 277.050 93.150 ;
        RECT 177.750 85.200 184.050 86.100 ;
        RECT 184.950 86.700 186.750 87.300 ;
        RECT 184.950 85.500 192.450 86.700 ;
        RECT 177.750 84.600 179.550 85.200 ;
        RECT 191.250 84.600 192.450 85.500 ;
        RECT 172.950 81.600 176.850 83.700 ;
        RECT 181.950 82.500 188.850 84.300 ;
        RECT 191.250 82.500 196.050 84.600 ;
        RECT 170.550 75.750 172.350 78.600 ;
        RECT 175.050 75.750 176.850 81.600 ;
        RECT 179.250 75.750 181.050 81.600 ;
        RECT 183.150 75.750 184.950 82.500 ;
        RECT 191.250 81.600 192.450 82.500 ;
        RECT 186.150 75.750 187.950 81.600 ;
        RECT 190.950 75.750 192.750 81.600 ;
        RECT 196.050 75.750 197.850 81.600 ;
        RECT 199.050 75.750 200.850 87.600 ;
        RECT 230.550 75.750 232.350 87.600 ;
        RECT 234.750 75.750 236.550 87.600 ;
        RECT 271.050 75.750 272.850 87.600 ;
        RECT 274.050 75.750 275.850 87.600 ;
        RECT 278.100 81.600 279.300 98.700 ;
        RECT 280.950 92.850 283.050 94.950 ;
        RECT 314.100 93.150 315.900 94.950 ;
        RECT 281.100 91.050 282.900 92.850 ;
        RECT 313.950 91.050 316.050 93.150 ;
        RECT 317.550 91.950 318.750 99.300 ;
        RECT 320.100 93.150 321.900 94.950 ;
        RECT 356.100 93.150 357.900 94.950 ;
        RECT 316.950 89.850 319.050 91.950 ;
        RECT 319.950 91.050 322.050 93.150 ;
        RECT 355.950 91.050 358.050 93.150 ;
        RECT 359.550 91.950 360.750 99.300 ;
        RECT 398.700 98.400 400.500 107.250 ;
        RECT 404.100 99.000 405.900 107.250 ;
        RECT 443.550 104.400 445.350 107.250 ;
        RECT 446.550 104.400 448.350 107.250 ;
        RECT 479.550 104.400 481.350 107.250 ;
        RECT 482.550 104.400 484.350 107.250 ;
        RECT 404.100 97.350 408.600 99.000 ;
        RECT 362.100 93.150 363.900 94.950 ;
        RECT 407.400 93.150 408.600 97.350 ;
        RECT 442.950 95.850 445.050 97.950 ;
        RECT 446.400 96.150 447.600 104.400 ;
        RECT 443.100 94.050 444.900 95.850 ;
        RECT 445.950 94.050 448.050 96.150 ;
        RECT 478.950 95.850 481.050 97.950 ;
        RECT 482.400 96.150 483.600 104.400 ;
        RECT 488.550 101.400 490.350 107.250 ;
        RECT 491.850 104.400 493.650 107.250 ;
        RECT 496.350 104.400 498.150 107.250 ;
        RECT 500.550 104.400 502.350 107.250 ;
        RECT 504.450 104.400 506.250 107.250 ;
        RECT 507.750 104.400 509.550 107.250 ;
        RECT 512.250 105.300 514.050 107.250 ;
        RECT 512.250 104.400 516.000 105.300 ;
        RECT 517.050 104.400 518.850 107.250 ;
        RECT 496.650 103.500 497.700 104.400 ;
        RECT 493.950 102.300 497.700 103.500 ;
        RECT 505.200 102.600 506.250 104.400 ;
        RECT 514.950 103.500 516.000 104.400 ;
        RECT 493.950 101.400 496.050 102.300 ;
        RECT 488.550 99.150 489.750 101.400 ;
        RECT 501.150 100.200 502.950 102.000 ;
        RECT 505.200 101.550 510.150 102.600 ;
        RECT 508.350 100.800 510.150 101.550 ;
        RECT 511.650 100.800 513.450 102.600 ;
        RECT 514.950 101.400 517.050 103.500 ;
        RECT 520.050 101.400 521.850 107.250 ;
        RECT 502.050 99.900 502.950 100.200 ;
        RECT 512.100 99.900 513.150 100.800 ;
        RECT 488.550 97.050 493.050 99.150 ;
        RECT 502.050 99.000 513.150 99.900 ;
        RECT 479.100 94.050 480.900 95.850 ;
        RECT 481.950 94.050 484.050 96.150 ;
        RECT 358.950 89.850 361.050 91.950 ;
        RECT 361.950 91.050 364.050 93.150 ;
        RECT 397.950 89.850 400.050 91.950 ;
        RECT 403.950 89.850 406.050 91.950 ;
        RECT 406.950 91.050 409.050 93.150 ;
        RECT 317.550 81.600 318.750 89.850 ;
        RECT 359.550 81.600 360.750 89.850 ;
        RECT 398.100 88.050 399.900 89.850 ;
        RECT 400.950 86.850 403.050 88.950 ;
        RECT 404.250 88.050 406.050 89.850 ;
        RECT 401.100 85.050 402.900 86.850 ;
        RECT 407.700 82.800 408.750 91.050 ;
        RECT 401.700 81.900 408.750 82.800 ;
        RECT 401.700 81.600 403.350 81.900 ;
        RECT 277.650 75.750 279.450 81.600 ;
        RECT 280.650 75.750 282.450 81.600 ;
        RECT 314.550 75.750 316.350 81.600 ;
        RECT 317.550 75.750 319.350 81.600 ;
        RECT 320.550 75.750 322.350 81.600 ;
        RECT 356.550 75.750 358.350 81.600 ;
        RECT 359.550 75.750 361.350 81.600 ;
        RECT 362.550 75.750 364.350 81.600 ;
        RECT 398.550 75.750 400.350 81.600 ;
        RECT 401.550 75.750 403.350 81.600 ;
        RECT 407.550 81.600 408.750 81.900 ;
        RECT 446.400 81.600 447.600 94.050 ;
        RECT 482.400 81.600 483.600 94.050 ;
        RECT 488.550 87.600 489.750 97.050 ;
        RECT 490.950 95.250 494.850 97.050 ;
        RECT 490.950 94.950 493.050 95.250 ;
        RECT 502.050 94.950 502.950 99.000 ;
        RECT 512.100 97.800 513.150 99.000 ;
        RECT 512.100 96.600 519.000 97.800 ;
        RECT 512.100 96.000 513.900 96.600 ;
        RECT 518.100 95.850 519.000 96.600 ;
        RECT 515.100 94.950 516.900 95.700 ;
        RECT 502.050 92.850 505.050 94.950 ;
        RECT 508.950 93.900 516.900 94.950 ;
        RECT 518.100 94.050 519.900 95.850 ;
        RECT 508.950 92.850 511.050 93.900 ;
        RECT 490.950 89.400 492.750 91.200 ;
        RECT 491.850 88.200 496.050 89.400 ;
        RECT 502.050 88.200 502.950 92.850 ;
        RECT 510.750 89.100 512.550 89.400 ;
        RECT 404.550 75.750 406.350 81.000 ;
        RECT 407.550 75.750 409.350 81.600 ;
        RECT 443.550 75.750 445.350 81.600 ;
        RECT 446.550 75.750 448.350 81.600 ;
        RECT 479.550 75.750 481.350 81.600 ;
        RECT 482.550 75.750 484.350 81.600 ;
        RECT 488.550 75.750 490.350 87.600 ;
        RECT 493.950 87.300 496.050 88.200 ;
        RECT 496.950 87.300 502.950 88.200 ;
        RECT 504.150 88.800 512.550 89.100 ;
        RECT 520.950 88.800 521.850 101.400 ;
        RECT 554.550 102.300 556.350 107.250 ;
        RECT 557.550 103.200 559.350 107.250 ;
        RECT 560.550 102.300 562.350 107.250 ;
        RECT 554.550 100.950 562.350 102.300 ;
        RECT 563.550 101.400 565.350 107.250 ;
        RECT 563.550 99.300 564.750 101.400 ;
        RECT 602.850 100.200 604.650 107.250 ;
        RECT 607.350 101.400 609.150 107.250 ;
        RECT 641.550 101.400 643.350 107.250 ;
        RECT 644.550 101.400 646.350 107.250 ;
        RECT 647.550 101.400 649.350 107.250 ;
        RECT 644.400 100.500 646.200 101.400 ;
        RECT 650.550 100.500 652.350 107.250 ;
        RECT 653.550 101.400 655.350 107.250 ;
        RECT 656.550 101.400 658.350 107.250 ;
        RECT 659.550 101.400 661.350 107.250 ;
        RECT 662.550 101.400 664.350 107.250 ;
        RECT 665.550 101.400 667.350 107.250 ;
        RECT 701.550 104.400 703.350 107.250 ;
        RECT 704.550 104.400 706.350 107.250 ;
        RECT 656.400 100.500 658.200 101.400 ;
        RECT 662.400 100.500 664.200 101.400 ;
        RECT 602.850 99.300 606.450 100.200 ;
        RECT 644.400 99.300 648.450 100.500 ;
        RECT 650.550 99.300 654.300 100.500 ;
        RECT 656.400 99.300 660.300 100.500 ;
        RECT 662.400 100.350 665.100 100.500 ;
        RECT 662.400 99.300 665.250 100.350 ;
        RECT 561.000 98.250 564.750 99.300 ;
        RECT 557.100 96.150 558.900 97.950 ;
        RECT 553.950 92.850 556.050 94.950 ;
        RECT 556.950 94.050 559.050 96.150 ;
        RECT 560.850 94.950 562.050 98.250 ;
        RECT 559.950 92.850 562.050 94.950 ;
        RECT 602.100 93.150 603.900 94.950 ;
        RECT 554.100 91.050 555.900 92.850 ;
        RECT 504.150 88.200 521.850 88.800 ;
        RECT 496.950 86.400 497.850 87.300 ;
        RECT 495.150 84.600 497.850 86.400 ;
        RECT 498.750 86.100 500.550 86.400 ;
        RECT 504.150 86.100 505.050 88.200 ;
        RECT 510.750 87.600 521.850 88.200 ;
        RECT 559.950 87.600 561.150 92.850 ;
        RECT 562.950 89.850 565.050 91.950 ;
        RECT 601.950 91.050 604.050 93.150 ;
        RECT 605.250 91.950 606.450 99.300 ;
        RECT 647.250 98.400 648.450 99.300 ;
        RECT 653.100 98.400 654.300 99.300 ;
        RECT 659.100 98.400 660.300 99.300 ;
        RECT 644.100 96.150 645.900 97.950 ;
        RECT 647.250 96.600 651.300 98.400 ;
        RECT 653.100 96.600 657.300 98.400 ;
        RECT 659.100 96.600 663.300 98.400 ;
        RECT 608.100 93.150 609.900 94.950 ;
        RECT 643.950 94.050 646.050 96.150 ;
        RECT 604.950 89.850 607.050 91.950 ;
        RECT 607.950 91.050 610.050 93.150 ;
        RECT 562.950 88.050 564.750 89.850 ;
        RECT 498.750 85.200 505.050 86.100 ;
        RECT 505.950 86.700 507.750 87.300 ;
        RECT 505.950 85.500 513.450 86.700 ;
        RECT 498.750 84.600 500.550 85.200 ;
        RECT 512.250 84.600 513.450 85.500 ;
        RECT 493.950 81.600 497.850 83.700 ;
        RECT 502.950 82.500 509.850 84.300 ;
        RECT 512.250 82.500 517.050 84.600 ;
        RECT 491.550 75.750 493.350 78.600 ;
        RECT 496.050 75.750 497.850 81.600 ;
        RECT 500.250 75.750 502.050 81.600 ;
        RECT 504.150 75.750 505.950 82.500 ;
        RECT 512.250 81.600 513.450 82.500 ;
        RECT 507.150 75.750 508.950 81.600 ;
        RECT 511.950 75.750 513.750 81.600 ;
        RECT 517.050 75.750 518.850 81.600 ;
        RECT 520.050 75.750 521.850 87.600 ;
        RECT 555.300 75.750 557.100 87.600 ;
        RECT 559.500 75.750 561.300 87.600 ;
        RECT 605.250 81.600 606.450 89.850 ;
        RECT 647.250 89.700 648.450 96.600 ;
        RECT 653.100 89.700 654.300 96.600 ;
        RECT 659.100 89.700 660.300 96.600 ;
        RECT 664.200 96.150 665.250 99.300 ;
        RECT 664.200 94.050 667.050 96.150 ;
        RECT 700.950 95.850 703.050 97.950 ;
        RECT 704.400 96.150 705.600 104.400 ;
        RECT 743.850 100.200 745.650 107.250 ;
        RECT 748.350 101.400 750.150 107.250 ;
        RECT 743.850 99.300 747.450 100.200 ;
        RECT 701.100 94.050 702.900 95.850 ;
        RECT 703.950 94.050 706.050 96.150 ;
        RECT 664.200 89.700 665.250 94.050 ;
        RECT 644.550 88.500 648.450 89.700 ;
        RECT 650.550 88.500 654.300 89.700 ;
        RECT 656.550 88.500 660.300 89.700 ;
        RECT 662.550 88.500 665.250 89.700 ;
        RECT 562.800 75.750 564.600 81.600 ;
        RECT 601.650 75.750 603.450 81.600 ;
        RECT 604.650 75.750 606.450 81.600 ;
        RECT 607.650 75.750 609.450 81.600 ;
        RECT 641.550 75.750 643.350 87.600 ;
        RECT 644.550 75.750 646.350 88.500 ;
        RECT 647.550 75.750 649.350 87.600 ;
        RECT 650.550 75.750 652.350 88.500 ;
        RECT 653.550 75.750 655.350 87.600 ;
        RECT 656.550 75.750 658.350 88.500 ;
        RECT 659.550 75.750 661.350 87.600 ;
        RECT 662.550 75.750 664.350 88.500 ;
        RECT 665.550 75.750 667.350 87.600 ;
        RECT 704.400 81.600 705.600 94.050 ;
        RECT 743.100 93.150 744.900 94.950 ;
        RECT 742.950 91.050 745.050 93.150 ;
        RECT 746.250 91.950 747.450 99.300 ;
        RECT 749.100 93.150 750.900 94.950 ;
        RECT 745.950 89.850 748.050 91.950 ;
        RECT 748.950 91.050 751.050 93.150 ;
        RECT 746.250 81.600 747.450 89.850 ;
        RECT 701.550 75.750 703.350 81.600 ;
        RECT 704.550 75.750 706.350 81.600 ;
        RECT 742.650 75.750 744.450 81.600 ;
        RECT 745.650 75.750 747.450 81.600 ;
        RECT 748.650 75.750 750.450 81.600 ;
        RECT 3.150 59.400 4.950 71.250 ;
        RECT 6.150 65.400 7.950 71.250 ;
        RECT 11.250 65.400 13.050 71.250 ;
        RECT 16.050 65.400 17.850 71.250 ;
        RECT 11.550 64.500 12.750 65.400 ;
        RECT 19.050 64.500 20.850 71.250 ;
        RECT 22.950 65.400 24.750 71.250 ;
        RECT 27.150 65.400 28.950 71.250 ;
        RECT 31.650 68.400 33.450 71.250 ;
        RECT 7.950 62.400 12.750 64.500 ;
        RECT 15.150 62.700 22.050 64.500 ;
        RECT 27.150 63.300 31.050 65.400 ;
        RECT 11.550 61.500 12.750 62.400 ;
        RECT 24.450 61.800 26.250 62.400 ;
        RECT 11.550 60.300 19.050 61.500 ;
        RECT 17.250 59.700 19.050 60.300 ;
        RECT 19.950 60.900 26.250 61.800 ;
        RECT 3.150 58.800 14.250 59.400 ;
        RECT 19.950 58.800 20.850 60.900 ;
        RECT 24.450 60.600 26.250 60.900 ;
        RECT 27.150 60.600 29.850 62.400 ;
        RECT 27.150 59.700 28.050 60.600 ;
        RECT 3.150 58.200 20.850 58.800 ;
        RECT 3.150 45.600 4.050 58.200 ;
        RECT 12.450 57.900 20.850 58.200 ;
        RECT 22.050 58.800 28.050 59.700 ;
        RECT 28.950 58.800 31.050 59.700 ;
        RECT 34.650 59.400 36.450 71.250 ;
        RECT 70.650 65.400 72.450 71.250 ;
        RECT 73.650 66.000 75.450 71.250 ;
        RECT 12.450 57.600 14.250 57.900 ;
        RECT 22.050 54.150 22.950 58.800 ;
        RECT 28.950 57.600 33.150 58.800 ;
        RECT 32.250 55.800 34.050 57.600 ;
        RECT 13.950 53.100 16.050 54.150 ;
        RECT 5.100 51.150 6.900 52.950 ;
        RECT 8.100 52.050 16.050 53.100 ;
        RECT 19.950 52.050 22.950 54.150 ;
        RECT 8.100 51.300 9.900 52.050 ;
        RECT 6.000 50.400 6.900 51.150 ;
        RECT 11.100 50.400 12.900 51.000 ;
        RECT 6.000 49.200 12.900 50.400 ;
        RECT 11.850 48.000 12.900 49.200 ;
        RECT 22.050 48.000 22.950 52.050 ;
        RECT 31.950 51.750 34.050 52.050 ;
        RECT 30.150 49.950 34.050 51.750 ;
        RECT 35.250 49.950 36.450 59.400 ;
        RECT 71.250 65.100 72.450 65.400 ;
        RECT 76.650 65.400 78.450 71.250 ;
        RECT 79.650 65.400 81.450 71.250 ;
        RECT 76.650 65.100 78.300 65.400 ;
        RECT 71.250 64.200 78.300 65.100 ;
        RECT 71.250 55.950 72.300 64.200 ;
        RECT 77.100 60.150 78.900 61.950 ;
        RECT 73.950 57.150 75.750 58.950 ;
        RECT 76.950 58.050 79.050 60.150 ;
        RECT 113.550 59.400 115.350 71.250 ;
        RECT 117.750 59.400 119.550 71.250 ;
        RECT 152.550 65.400 154.350 71.250 ;
        RECT 155.550 65.400 157.350 71.250 ;
        RECT 80.100 57.150 81.900 58.950 ;
        RECT 117.000 58.350 119.550 59.400 ;
        RECT 70.950 53.850 73.050 55.950 ;
        RECT 73.950 55.050 76.050 57.150 ;
        RECT 79.950 55.050 82.050 57.150 ;
        RECT 113.100 54.150 114.900 55.950 ;
        RECT 11.850 47.100 22.950 48.000 ;
        RECT 31.950 47.850 36.450 49.950 ;
        RECT 71.400 49.650 72.600 53.850 ;
        RECT 112.950 52.050 115.050 54.150 ;
        RECT 117.000 51.150 118.050 58.350 ;
        RECT 119.100 54.150 120.900 55.950 ;
        RECT 152.100 54.150 153.900 55.950 ;
        RECT 118.950 52.050 121.050 54.150 ;
        RECT 151.950 52.050 154.050 54.150 ;
        RECT 71.400 48.000 75.900 49.650 ;
        RECT 115.950 49.050 118.050 51.150 ;
        RECT 11.850 46.200 12.900 47.100 ;
        RECT 22.050 46.800 22.950 47.100 ;
        RECT 3.150 39.750 4.950 45.600 ;
        RECT 7.950 43.500 10.050 45.600 ;
        RECT 11.550 44.400 13.350 46.200 ;
        RECT 14.850 45.450 16.650 46.200 ;
        RECT 14.850 44.400 19.800 45.450 ;
        RECT 22.050 45.000 23.850 46.800 ;
        RECT 35.250 45.600 36.450 47.850 ;
        RECT 28.950 44.700 31.050 45.600 ;
        RECT 9.000 42.600 10.050 43.500 ;
        RECT 18.750 42.600 19.800 44.400 ;
        RECT 27.300 43.500 31.050 44.700 ;
        RECT 27.300 42.600 28.350 43.500 ;
        RECT 6.150 39.750 7.950 42.600 ;
        RECT 9.000 41.700 12.750 42.600 ;
        RECT 10.950 39.750 12.750 41.700 ;
        RECT 15.450 39.750 17.250 42.600 ;
        RECT 18.750 39.750 20.550 42.600 ;
        RECT 22.650 39.750 24.450 42.600 ;
        RECT 26.850 39.750 28.650 42.600 ;
        RECT 31.350 39.750 33.150 42.600 ;
        RECT 34.650 39.750 36.450 45.600 ;
        RECT 74.100 39.750 75.900 48.000 ;
        RECT 79.500 39.750 81.300 48.600 ;
        RECT 117.000 42.600 118.050 49.050 ;
        RECT 155.700 48.300 156.900 65.400 ;
        RECT 159.150 59.400 160.950 71.250 ;
        RECT 162.150 59.400 163.950 71.250 ;
        RECT 197.550 65.400 199.350 71.250 ;
        RECT 200.550 65.400 202.350 71.250 ;
        RECT 203.550 65.400 205.350 71.250 ;
        RECT 239.550 65.400 241.350 71.250 ;
        RECT 242.550 65.400 244.350 71.250 ;
        RECT 245.550 65.400 247.350 71.250 ;
        RECT 157.950 53.850 160.050 55.950 ;
        RECT 162.150 54.150 163.350 59.400 ;
        RECT 200.550 57.150 201.750 65.400 ;
        RECT 242.550 57.150 243.750 65.400 ;
        RECT 281.550 59.400 283.350 71.250 ;
        RECT 285.750 59.400 287.550 71.250 ;
        RECT 322.650 65.400 324.450 71.250 ;
        RECT 325.650 65.400 327.450 71.250 ;
        RECT 285.000 58.350 287.550 59.400 ;
        RECT 158.100 52.050 159.900 53.850 ;
        RECT 160.950 52.050 163.350 54.150 ;
        RECT 196.950 53.850 199.050 55.950 ;
        RECT 199.950 55.050 202.050 57.150 ;
        RECT 197.100 52.050 198.900 53.850 ;
        RECT 152.550 47.100 160.050 48.300 ;
        RECT 113.550 39.750 115.350 42.600 ;
        RECT 116.550 39.750 118.350 42.600 ;
        RECT 119.550 39.750 121.350 42.600 ;
        RECT 152.550 39.750 154.350 47.100 ;
        RECT 158.250 46.500 160.050 47.100 ;
        RECT 162.150 45.600 163.350 52.050 ;
        RECT 200.550 47.700 201.750 55.050 ;
        RECT 202.950 53.850 205.050 55.950 ;
        RECT 238.950 53.850 241.050 55.950 ;
        RECT 241.950 55.050 244.050 57.150 ;
        RECT 203.100 52.050 204.900 53.850 ;
        RECT 239.100 52.050 240.900 53.850 ;
        RECT 242.550 47.700 243.750 55.050 ;
        RECT 244.950 53.850 247.050 55.950 ;
        RECT 281.100 54.150 282.900 55.950 ;
        RECT 245.100 52.050 246.900 53.850 ;
        RECT 280.950 52.050 283.050 54.150 ;
        RECT 285.000 51.150 286.050 58.350 ;
        RECT 287.100 54.150 288.900 55.950 ;
        RECT 286.950 52.050 289.050 54.150 ;
        RECT 323.400 52.950 324.600 65.400 ;
        RECT 363.450 59.400 365.250 71.250 ;
        RECT 367.650 59.400 369.450 71.250 ;
        RECT 400.650 65.400 402.450 71.250 ;
        RECT 403.650 65.400 405.450 71.250 ;
        RECT 363.450 58.350 366.000 59.400 ;
        RECT 362.100 54.150 363.900 55.950 ;
        RECT 283.950 49.050 286.050 51.150 ;
        RECT 322.950 50.850 325.050 52.950 ;
        RECT 326.100 51.150 327.900 52.950 ;
        RECT 361.950 52.050 364.050 54.150 ;
        RECT 364.950 51.150 366.000 58.350 ;
        RECT 368.100 54.150 369.900 55.950 ;
        RECT 367.950 52.050 370.050 54.150 ;
        RECT 401.400 52.950 402.600 65.400 ;
        RECT 408.150 59.400 409.950 71.250 ;
        RECT 411.150 65.400 412.950 71.250 ;
        RECT 416.250 65.400 418.050 71.250 ;
        RECT 421.050 65.400 422.850 71.250 ;
        RECT 416.550 64.500 417.750 65.400 ;
        RECT 424.050 64.500 425.850 71.250 ;
        RECT 427.950 65.400 429.750 71.250 ;
        RECT 432.150 65.400 433.950 71.250 ;
        RECT 436.650 68.400 438.450 71.250 ;
        RECT 412.950 62.400 417.750 64.500 ;
        RECT 420.150 62.700 427.050 64.500 ;
        RECT 432.150 63.300 436.050 65.400 ;
        RECT 416.550 61.500 417.750 62.400 ;
        RECT 429.450 61.800 431.250 62.400 ;
        RECT 416.550 60.300 424.050 61.500 ;
        RECT 422.250 59.700 424.050 60.300 ;
        RECT 424.950 60.900 431.250 61.800 ;
        RECT 408.150 58.800 419.250 59.400 ;
        RECT 424.950 58.800 425.850 60.900 ;
        RECT 429.450 60.600 431.250 60.900 ;
        RECT 432.150 60.600 434.850 62.400 ;
        RECT 432.150 59.700 433.050 60.600 ;
        RECT 408.150 58.200 425.850 58.800 ;
        RECT 200.550 46.800 204.150 47.700 ;
        RECT 242.550 46.800 246.150 47.700 ;
        RECT 157.050 39.750 158.850 45.600 ;
        RECT 160.050 44.100 163.350 45.600 ;
        RECT 160.050 39.750 161.850 44.100 ;
        RECT 197.850 39.750 199.650 45.600 ;
        RECT 202.350 39.750 204.150 46.800 ;
        RECT 239.850 39.750 241.650 45.600 ;
        RECT 244.350 39.750 246.150 46.800 ;
        RECT 285.000 42.600 286.050 49.050 ;
        RECT 323.400 42.600 324.600 50.850 ;
        RECT 325.950 49.050 328.050 51.150 ;
        RECT 364.950 49.050 367.050 51.150 ;
        RECT 400.950 50.850 403.050 52.950 ;
        RECT 404.100 51.150 405.900 52.950 ;
        RECT 364.950 42.600 366.000 49.050 ;
        RECT 401.400 42.600 402.600 50.850 ;
        RECT 403.950 49.050 406.050 51.150 ;
        RECT 408.150 45.600 409.050 58.200 ;
        RECT 417.450 57.900 425.850 58.200 ;
        RECT 427.050 58.800 433.050 59.700 ;
        RECT 433.950 58.800 436.050 59.700 ;
        RECT 439.650 59.400 441.450 71.250 ;
        RECT 417.450 57.600 419.250 57.900 ;
        RECT 427.050 54.150 427.950 58.800 ;
        RECT 433.950 57.600 438.150 58.800 ;
        RECT 437.250 55.800 439.050 57.600 ;
        RECT 418.950 53.100 421.050 54.150 ;
        RECT 410.100 51.150 411.900 52.950 ;
        RECT 413.100 52.050 421.050 53.100 ;
        RECT 424.950 52.050 427.950 54.150 ;
        RECT 413.100 51.300 414.900 52.050 ;
        RECT 411.000 50.400 411.900 51.150 ;
        RECT 416.100 50.400 417.900 51.000 ;
        RECT 411.000 49.200 417.900 50.400 ;
        RECT 416.850 48.000 417.900 49.200 ;
        RECT 427.050 48.000 427.950 52.050 ;
        RECT 436.950 51.750 439.050 52.050 ;
        RECT 435.150 49.950 439.050 51.750 ;
        RECT 440.250 49.950 441.450 59.400 ;
        RECT 416.850 47.100 427.950 48.000 ;
        RECT 436.950 47.850 441.450 49.950 ;
        RECT 416.850 46.200 417.900 47.100 ;
        RECT 427.050 46.800 427.950 47.100 ;
        RECT 281.550 39.750 283.350 42.600 ;
        RECT 284.550 39.750 286.350 42.600 ;
        RECT 287.550 39.750 289.350 42.600 ;
        RECT 322.650 39.750 324.450 42.600 ;
        RECT 325.650 39.750 327.450 42.600 ;
        RECT 361.650 39.750 363.450 42.600 ;
        RECT 364.650 39.750 366.450 42.600 ;
        RECT 367.650 39.750 369.450 42.600 ;
        RECT 400.650 39.750 402.450 42.600 ;
        RECT 403.650 39.750 405.450 42.600 ;
        RECT 408.150 39.750 409.950 45.600 ;
        RECT 412.950 43.500 415.050 45.600 ;
        RECT 416.550 44.400 418.350 46.200 ;
        RECT 419.850 45.450 421.650 46.200 ;
        RECT 419.850 44.400 424.800 45.450 ;
        RECT 427.050 45.000 428.850 46.800 ;
        RECT 440.250 45.600 441.450 47.850 ;
        RECT 433.950 44.700 436.050 45.600 ;
        RECT 414.000 42.600 415.050 43.500 ;
        RECT 423.750 42.600 424.800 44.400 ;
        RECT 432.300 43.500 436.050 44.700 ;
        RECT 432.300 42.600 433.350 43.500 ;
        RECT 411.150 39.750 412.950 42.600 ;
        RECT 414.000 41.700 417.750 42.600 ;
        RECT 415.950 39.750 417.750 41.700 ;
        RECT 420.450 39.750 422.250 42.600 ;
        RECT 423.750 39.750 425.550 42.600 ;
        RECT 427.650 39.750 429.450 42.600 ;
        RECT 431.850 39.750 433.650 42.600 ;
        RECT 436.350 39.750 438.150 42.600 ;
        RECT 439.650 39.750 441.450 45.600 ;
        RECT 443.550 59.400 445.350 71.250 ;
        RECT 446.550 68.400 448.350 71.250 ;
        RECT 451.050 65.400 452.850 71.250 ;
        RECT 455.250 65.400 457.050 71.250 ;
        RECT 448.950 63.300 452.850 65.400 ;
        RECT 459.150 64.500 460.950 71.250 ;
        RECT 462.150 65.400 463.950 71.250 ;
        RECT 466.950 65.400 468.750 71.250 ;
        RECT 472.050 65.400 473.850 71.250 ;
        RECT 467.250 64.500 468.450 65.400 ;
        RECT 457.950 62.700 464.850 64.500 ;
        RECT 467.250 62.400 472.050 64.500 ;
        RECT 450.150 60.600 452.850 62.400 ;
        RECT 453.750 61.800 455.550 62.400 ;
        RECT 453.750 60.900 460.050 61.800 ;
        RECT 467.250 61.500 468.450 62.400 ;
        RECT 453.750 60.600 455.550 60.900 ;
        RECT 451.950 59.700 452.850 60.600 ;
        RECT 443.550 49.950 444.750 59.400 ;
        RECT 448.950 58.800 451.050 59.700 ;
        RECT 451.950 58.800 457.950 59.700 ;
        RECT 446.850 57.600 451.050 58.800 ;
        RECT 445.950 55.800 447.750 57.600 ;
        RECT 457.050 54.150 457.950 58.800 ;
        RECT 459.150 58.800 460.050 60.900 ;
        RECT 460.950 60.300 468.450 61.500 ;
        RECT 460.950 59.700 462.750 60.300 ;
        RECT 475.050 59.400 476.850 71.250 ;
        RECT 509.550 65.400 511.350 71.250 ;
        RECT 512.550 65.400 514.350 71.250 ;
        RECT 550.650 65.400 552.450 71.250 ;
        RECT 553.650 65.400 555.450 71.250 ;
        RECT 556.650 65.400 558.450 71.250 ;
        RECT 593.400 65.400 595.200 71.250 ;
        RECT 465.750 58.800 476.850 59.400 ;
        RECT 459.150 58.200 476.850 58.800 ;
        RECT 459.150 57.900 467.550 58.200 ;
        RECT 465.750 57.600 467.550 57.900 ;
        RECT 457.050 52.050 460.050 54.150 ;
        RECT 463.950 53.100 466.050 54.150 ;
        RECT 463.950 52.050 471.900 53.100 ;
        RECT 445.950 51.750 448.050 52.050 ;
        RECT 445.950 49.950 449.850 51.750 ;
        RECT 443.550 47.850 448.050 49.950 ;
        RECT 457.050 48.000 457.950 52.050 ;
        RECT 470.100 51.300 471.900 52.050 ;
        RECT 473.100 51.150 474.900 52.950 ;
        RECT 467.100 50.400 468.900 51.000 ;
        RECT 473.100 50.400 474.000 51.150 ;
        RECT 467.100 49.200 474.000 50.400 ;
        RECT 467.100 48.000 468.150 49.200 ;
        RECT 443.550 45.600 444.750 47.850 ;
        RECT 457.050 47.100 468.150 48.000 ;
        RECT 457.050 46.800 457.950 47.100 ;
        RECT 443.550 39.750 445.350 45.600 ;
        RECT 448.950 44.700 451.050 45.600 ;
        RECT 456.150 45.000 457.950 46.800 ;
        RECT 467.100 46.200 468.150 47.100 ;
        RECT 463.350 45.450 465.150 46.200 ;
        RECT 448.950 43.500 452.700 44.700 ;
        RECT 451.650 42.600 452.700 43.500 ;
        RECT 460.200 44.400 465.150 45.450 ;
        RECT 466.650 44.400 468.450 46.200 ;
        RECT 475.950 45.600 476.850 58.200 ;
        RECT 512.400 52.950 513.600 65.400 ;
        RECT 554.250 57.150 555.450 65.400 ;
        RECT 596.700 59.400 598.500 71.250 ;
        RECT 600.900 59.400 602.700 71.250 ;
        RECT 606.150 59.400 607.950 71.250 ;
        RECT 609.150 65.400 610.950 71.250 ;
        RECT 614.250 65.400 616.050 71.250 ;
        RECT 619.050 65.400 620.850 71.250 ;
        RECT 614.550 64.500 615.750 65.400 ;
        RECT 622.050 64.500 623.850 71.250 ;
        RECT 625.950 65.400 627.750 71.250 ;
        RECT 630.150 65.400 631.950 71.250 ;
        RECT 634.650 68.400 636.450 71.250 ;
        RECT 610.950 62.400 615.750 64.500 ;
        RECT 618.150 62.700 625.050 64.500 ;
        RECT 630.150 63.300 634.050 65.400 ;
        RECT 614.550 61.500 615.750 62.400 ;
        RECT 627.450 61.800 629.250 62.400 ;
        RECT 614.550 60.300 622.050 61.500 ;
        RECT 620.250 59.700 622.050 60.300 ;
        RECT 622.950 60.900 629.250 61.800 ;
        RECT 593.250 57.150 595.050 58.950 ;
        RECT 550.950 53.850 553.050 55.950 ;
        RECT 553.950 55.050 556.050 57.150 ;
        RECT 509.100 51.150 510.900 52.950 ;
        RECT 508.950 49.050 511.050 51.150 ;
        RECT 511.950 50.850 514.050 52.950 ;
        RECT 551.100 52.050 552.900 53.850 ;
        RECT 460.200 42.600 461.250 44.400 ;
        RECT 469.950 43.500 472.050 45.600 ;
        RECT 469.950 42.600 471.000 43.500 ;
        RECT 446.850 39.750 448.650 42.600 ;
        RECT 451.350 39.750 453.150 42.600 ;
        RECT 455.550 39.750 457.350 42.600 ;
        RECT 459.450 39.750 461.250 42.600 ;
        RECT 462.750 39.750 464.550 42.600 ;
        RECT 467.250 41.700 471.000 42.600 ;
        RECT 467.250 39.750 469.050 41.700 ;
        RECT 472.050 39.750 473.850 42.600 ;
        RECT 475.050 39.750 476.850 45.600 ;
        RECT 512.400 42.600 513.600 50.850 ;
        RECT 554.250 47.700 555.450 55.050 ;
        RECT 556.950 53.850 559.050 55.950 ;
        RECT 592.950 55.050 595.050 57.150 ;
        RECT 596.850 54.150 598.050 59.400 ;
        RECT 606.150 58.800 617.250 59.400 ;
        RECT 622.950 58.800 623.850 60.900 ;
        RECT 627.450 60.600 629.250 60.900 ;
        RECT 630.150 60.600 632.850 62.400 ;
        RECT 630.150 59.700 631.050 60.600 ;
        RECT 606.150 58.200 623.850 58.800 ;
        RECT 602.100 54.150 603.900 55.950 ;
        RECT 557.100 52.050 558.900 53.850 ;
        RECT 595.950 52.050 598.050 54.150 ;
        RECT 595.950 48.750 597.150 52.050 ;
        RECT 598.950 50.850 601.050 52.950 ;
        RECT 601.950 52.050 604.050 54.150 ;
        RECT 599.100 49.050 600.900 50.850 ;
        RECT 551.850 46.800 555.450 47.700 ;
        RECT 593.250 47.700 597.000 48.750 ;
        RECT 509.550 39.750 511.350 42.600 ;
        RECT 512.550 39.750 514.350 42.600 ;
        RECT 551.850 39.750 553.650 46.800 ;
        RECT 593.250 45.600 594.450 47.700 ;
        RECT 556.350 39.750 558.150 45.600 ;
        RECT 592.650 39.750 594.450 45.600 ;
        RECT 595.650 44.700 603.450 46.050 ;
        RECT 595.650 39.750 597.450 44.700 ;
        RECT 598.650 39.750 600.450 43.800 ;
        RECT 601.650 39.750 603.450 44.700 ;
        RECT 606.150 45.600 607.050 58.200 ;
        RECT 615.450 57.900 623.850 58.200 ;
        RECT 625.050 58.800 631.050 59.700 ;
        RECT 631.950 58.800 634.050 59.700 ;
        RECT 637.650 59.400 639.450 71.250 ;
        RECT 671.550 65.400 673.350 71.250 ;
        RECT 674.550 65.400 676.350 71.250 ;
        RECT 677.550 65.400 679.350 71.250 ;
        RECT 710.550 65.400 712.350 71.250 ;
        RECT 713.550 65.400 715.350 71.250 ;
        RECT 716.550 65.400 718.350 71.250 ;
        RECT 752.550 65.400 754.350 71.250 ;
        RECT 755.550 65.400 757.350 71.250 ;
        RECT 615.450 57.600 617.250 57.900 ;
        RECT 625.050 54.150 625.950 58.800 ;
        RECT 631.950 57.600 636.150 58.800 ;
        RECT 635.250 55.800 637.050 57.600 ;
        RECT 616.950 53.100 619.050 54.150 ;
        RECT 608.100 51.150 609.900 52.950 ;
        RECT 611.100 52.050 619.050 53.100 ;
        RECT 622.950 52.050 625.950 54.150 ;
        RECT 611.100 51.300 612.900 52.050 ;
        RECT 609.000 50.400 609.900 51.150 ;
        RECT 614.100 50.400 615.900 51.000 ;
        RECT 609.000 49.200 615.900 50.400 ;
        RECT 614.850 48.000 615.900 49.200 ;
        RECT 625.050 48.000 625.950 52.050 ;
        RECT 634.950 51.750 637.050 52.050 ;
        RECT 633.150 49.950 637.050 51.750 ;
        RECT 638.250 49.950 639.450 59.400 ;
        RECT 674.550 57.150 675.750 65.400 ;
        RECT 713.550 57.150 714.750 65.400 ;
        RECT 670.950 53.850 673.050 55.950 ;
        RECT 673.950 55.050 676.050 57.150 ;
        RECT 671.100 52.050 672.900 53.850 ;
        RECT 614.850 47.100 625.950 48.000 ;
        RECT 634.950 47.850 639.450 49.950 ;
        RECT 614.850 46.200 615.900 47.100 ;
        RECT 625.050 46.800 625.950 47.100 ;
        RECT 606.150 39.750 607.950 45.600 ;
        RECT 610.950 43.500 613.050 45.600 ;
        RECT 614.550 44.400 616.350 46.200 ;
        RECT 617.850 45.450 619.650 46.200 ;
        RECT 617.850 44.400 622.800 45.450 ;
        RECT 625.050 45.000 626.850 46.800 ;
        RECT 638.250 45.600 639.450 47.850 ;
        RECT 674.550 47.700 675.750 55.050 ;
        RECT 676.950 53.850 679.050 55.950 ;
        RECT 709.950 53.850 712.050 55.950 ;
        RECT 712.950 55.050 715.050 57.150 ;
        RECT 677.100 52.050 678.900 53.850 ;
        RECT 710.100 52.050 711.900 53.850 ;
        RECT 713.550 47.700 714.750 55.050 ;
        RECT 715.950 53.850 718.050 55.950 ;
        RECT 716.100 52.050 717.900 53.850 ;
        RECT 755.400 52.950 756.600 65.400 ;
        RECT 752.100 51.150 753.900 52.950 ;
        RECT 751.950 49.050 754.050 51.150 ;
        RECT 754.950 50.850 757.050 52.950 ;
        RECT 674.550 46.800 678.150 47.700 ;
        RECT 713.550 46.800 717.150 47.700 ;
        RECT 631.950 44.700 634.050 45.600 ;
        RECT 612.000 42.600 613.050 43.500 ;
        RECT 621.750 42.600 622.800 44.400 ;
        RECT 630.300 43.500 634.050 44.700 ;
        RECT 630.300 42.600 631.350 43.500 ;
        RECT 609.150 39.750 610.950 42.600 ;
        RECT 612.000 41.700 615.750 42.600 ;
        RECT 613.950 39.750 615.750 41.700 ;
        RECT 618.450 39.750 620.250 42.600 ;
        RECT 621.750 39.750 623.550 42.600 ;
        RECT 625.650 39.750 627.450 42.600 ;
        RECT 629.850 39.750 631.650 42.600 ;
        RECT 634.350 39.750 636.150 42.600 ;
        RECT 637.650 39.750 639.450 45.600 ;
        RECT 671.850 39.750 673.650 45.600 ;
        RECT 676.350 39.750 678.150 46.800 ;
        RECT 710.850 39.750 712.650 45.600 ;
        RECT 715.350 39.750 717.150 46.800 ;
        RECT 755.400 42.600 756.600 50.850 ;
        RECT 752.550 39.750 754.350 42.600 ;
        RECT 755.550 39.750 757.350 42.600 ;
        RECT 31.650 32.400 33.450 35.250 ;
        RECT 34.650 32.400 36.450 35.250 ;
        RECT 32.400 24.150 33.600 32.400 ;
        RECT 39.150 29.400 40.950 35.250 ;
        RECT 42.150 32.400 43.950 35.250 ;
        RECT 46.950 33.300 48.750 35.250 ;
        RECT 45.000 32.400 48.750 33.300 ;
        RECT 51.450 32.400 53.250 35.250 ;
        RECT 54.750 32.400 56.550 35.250 ;
        RECT 58.650 32.400 60.450 35.250 ;
        RECT 62.850 32.400 64.650 35.250 ;
        RECT 67.350 32.400 69.150 35.250 ;
        RECT 45.000 31.500 46.050 32.400 ;
        RECT 43.950 29.400 46.050 31.500 ;
        RECT 54.750 30.600 55.800 32.400 ;
        RECT 31.950 22.050 34.050 24.150 ;
        RECT 34.950 23.850 37.050 25.950 ;
        RECT 35.100 22.050 36.900 23.850 ;
        RECT 32.400 9.600 33.600 22.050 ;
        RECT 39.150 16.800 40.050 29.400 ;
        RECT 47.550 28.800 49.350 30.600 ;
        RECT 50.850 29.550 55.800 30.600 ;
        RECT 63.300 31.500 64.350 32.400 ;
        RECT 63.300 30.300 67.050 31.500 ;
        RECT 50.850 28.800 52.650 29.550 ;
        RECT 47.850 27.900 48.900 28.800 ;
        RECT 58.050 28.200 59.850 30.000 ;
        RECT 64.950 29.400 67.050 30.300 ;
        RECT 70.650 29.400 72.450 35.250 ;
        RECT 104.550 32.400 106.350 35.250 ;
        RECT 107.550 32.400 109.350 35.250 ;
        RECT 110.550 32.400 112.350 35.250 ;
        RECT 148.650 32.400 150.450 35.250 ;
        RECT 151.650 32.400 153.450 35.250 ;
        RECT 58.050 27.900 58.950 28.200 ;
        RECT 47.850 27.000 58.950 27.900 ;
        RECT 71.250 27.150 72.450 29.400 ;
        RECT 47.850 25.800 48.900 27.000 ;
        RECT 42.000 24.600 48.900 25.800 ;
        RECT 42.000 23.850 42.900 24.600 ;
        RECT 47.100 24.000 48.900 24.600 ;
        RECT 41.100 22.050 42.900 23.850 ;
        RECT 44.100 22.950 45.900 23.700 ;
        RECT 58.050 22.950 58.950 27.000 ;
        RECT 67.950 25.050 72.450 27.150 ;
        RECT 108.000 25.950 109.050 32.400 ;
        RECT 66.150 23.250 70.050 25.050 ;
        RECT 67.950 22.950 70.050 23.250 ;
        RECT 44.100 21.900 52.050 22.950 ;
        RECT 49.950 20.850 52.050 21.900 ;
        RECT 55.950 20.850 58.950 22.950 ;
        RECT 48.450 17.100 50.250 17.400 ;
        RECT 48.450 16.800 56.850 17.100 ;
        RECT 39.150 16.200 56.850 16.800 ;
        RECT 39.150 15.600 50.250 16.200 ;
        RECT 31.650 3.750 33.450 9.600 ;
        RECT 34.650 3.750 36.450 9.600 ;
        RECT 39.150 3.750 40.950 15.600 ;
        RECT 53.250 14.700 55.050 15.300 ;
        RECT 47.550 13.500 55.050 14.700 ;
        RECT 55.950 14.100 56.850 16.200 ;
        RECT 58.050 16.200 58.950 20.850 ;
        RECT 68.250 17.400 70.050 19.200 ;
        RECT 64.950 16.200 69.150 17.400 ;
        RECT 58.050 15.300 64.050 16.200 ;
        RECT 64.950 15.300 67.050 16.200 ;
        RECT 71.250 15.600 72.450 25.050 ;
        RECT 106.950 23.850 109.050 25.950 ;
        RECT 149.400 24.150 150.600 32.400 ;
        RECT 156.150 29.400 157.950 35.250 ;
        RECT 159.150 32.400 160.950 35.250 ;
        RECT 163.950 33.300 165.750 35.250 ;
        RECT 162.000 32.400 165.750 33.300 ;
        RECT 168.450 32.400 170.250 35.250 ;
        RECT 171.750 32.400 173.550 35.250 ;
        RECT 175.650 32.400 177.450 35.250 ;
        RECT 179.850 32.400 181.650 35.250 ;
        RECT 184.350 32.400 186.150 35.250 ;
        RECT 162.000 31.500 163.050 32.400 ;
        RECT 160.950 29.400 163.050 31.500 ;
        RECT 171.750 30.600 172.800 32.400 ;
        RECT 103.950 20.850 106.050 22.950 ;
        RECT 104.100 19.050 105.900 20.850 ;
        RECT 108.000 16.650 109.050 23.850 ;
        RECT 109.950 20.850 112.050 22.950 ;
        RECT 148.950 22.050 151.050 24.150 ;
        RECT 151.950 23.850 154.050 25.950 ;
        RECT 152.100 22.050 153.900 23.850 ;
        RECT 110.100 19.050 111.900 20.850 ;
        RECT 108.000 15.600 110.550 16.650 ;
        RECT 63.150 14.400 64.050 15.300 ;
        RECT 60.450 14.100 62.250 14.400 ;
        RECT 47.550 12.600 48.750 13.500 ;
        RECT 55.950 13.200 62.250 14.100 ;
        RECT 60.450 12.600 62.250 13.200 ;
        RECT 63.150 12.600 65.850 14.400 ;
        RECT 43.950 10.500 48.750 12.600 ;
        RECT 51.150 10.500 58.050 12.300 ;
        RECT 47.550 9.600 48.750 10.500 ;
        RECT 42.150 3.750 43.950 9.600 ;
        RECT 47.250 3.750 49.050 9.600 ;
        RECT 52.050 3.750 53.850 9.600 ;
        RECT 55.050 3.750 56.850 10.500 ;
        RECT 63.150 9.600 67.050 11.700 ;
        RECT 58.950 3.750 60.750 9.600 ;
        RECT 63.150 3.750 64.950 9.600 ;
        RECT 67.650 3.750 69.450 6.600 ;
        RECT 70.650 3.750 72.450 15.600 ;
        RECT 104.550 3.750 106.350 15.600 ;
        RECT 108.750 3.750 110.550 15.600 ;
        RECT 149.400 9.600 150.600 22.050 ;
        RECT 156.150 16.800 157.050 29.400 ;
        RECT 164.550 28.800 166.350 30.600 ;
        RECT 167.850 29.550 172.800 30.600 ;
        RECT 180.300 31.500 181.350 32.400 ;
        RECT 180.300 30.300 184.050 31.500 ;
        RECT 167.850 28.800 169.650 29.550 ;
        RECT 164.850 27.900 165.900 28.800 ;
        RECT 175.050 28.200 176.850 30.000 ;
        RECT 181.950 29.400 184.050 30.300 ;
        RECT 187.650 29.400 189.450 35.250 ;
        RECT 175.050 27.900 175.950 28.200 ;
        RECT 164.850 27.000 175.950 27.900 ;
        RECT 188.250 27.150 189.450 29.400 ;
        RECT 164.850 25.800 165.900 27.000 ;
        RECT 159.000 24.600 165.900 25.800 ;
        RECT 159.000 23.850 159.900 24.600 ;
        RECT 164.100 24.000 165.900 24.600 ;
        RECT 158.100 22.050 159.900 23.850 ;
        RECT 161.100 22.950 162.900 23.700 ;
        RECT 175.050 22.950 175.950 27.000 ;
        RECT 184.950 25.050 189.450 27.150 ;
        RECT 183.150 23.250 187.050 25.050 ;
        RECT 184.950 22.950 187.050 23.250 ;
        RECT 161.100 21.900 169.050 22.950 ;
        RECT 166.950 20.850 169.050 21.900 ;
        RECT 172.950 20.850 175.950 22.950 ;
        RECT 165.450 17.100 167.250 17.400 ;
        RECT 165.450 16.800 173.850 17.100 ;
        RECT 156.150 16.200 173.850 16.800 ;
        RECT 156.150 15.600 167.250 16.200 ;
        RECT 148.650 3.750 150.450 9.600 ;
        RECT 151.650 3.750 153.450 9.600 ;
        RECT 156.150 3.750 157.950 15.600 ;
        RECT 170.250 14.700 172.050 15.300 ;
        RECT 164.550 13.500 172.050 14.700 ;
        RECT 172.950 14.100 173.850 16.200 ;
        RECT 175.050 16.200 175.950 20.850 ;
        RECT 185.250 17.400 187.050 19.200 ;
        RECT 181.950 16.200 186.150 17.400 ;
        RECT 175.050 15.300 181.050 16.200 ;
        RECT 181.950 15.300 184.050 16.200 ;
        RECT 188.250 15.600 189.450 25.050 ;
        RECT 180.150 14.400 181.050 15.300 ;
        RECT 177.450 14.100 179.250 14.400 ;
        RECT 164.550 12.600 165.750 13.500 ;
        RECT 172.950 13.200 179.250 14.100 ;
        RECT 177.450 12.600 179.250 13.200 ;
        RECT 180.150 12.600 182.850 14.400 ;
        RECT 160.950 10.500 165.750 12.600 ;
        RECT 168.150 10.500 175.050 12.300 ;
        RECT 164.550 9.600 165.750 10.500 ;
        RECT 159.150 3.750 160.950 9.600 ;
        RECT 164.250 3.750 166.050 9.600 ;
        RECT 169.050 3.750 170.850 9.600 ;
        RECT 172.050 3.750 173.850 10.500 ;
        RECT 180.150 9.600 184.050 11.700 ;
        RECT 175.950 3.750 177.750 9.600 ;
        RECT 180.150 3.750 181.950 9.600 ;
        RECT 184.650 3.750 186.450 6.600 ;
        RECT 187.650 3.750 189.450 15.600 ;
        RECT 191.550 29.400 193.350 35.250 ;
        RECT 194.850 32.400 196.650 35.250 ;
        RECT 199.350 32.400 201.150 35.250 ;
        RECT 203.550 32.400 205.350 35.250 ;
        RECT 207.450 32.400 209.250 35.250 ;
        RECT 210.750 32.400 212.550 35.250 ;
        RECT 215.250 33.300 217.050 35.250 ;
        RECT 215.250 32.400 219.000 33.300 ;
        RECT 220.050 32.400 221.850 35.250 ;
        RECT 199.650 31.500 200.700 32.400 ;
        RECT 196.950 30.300 200.700 31.500 ;
        RECT 208.200 30.600 209.250 32.400 ;
        RECT 217.950 31.500 219.000 32.400 ;
        RECT 196.950 29.400 199.050 30.300 ;
        RECT 191.550 27.150 192.750 29.400 ;
        RECT 204.150 28.200 205.950 30.000 ;
        RECT 208.200 29.550 213.150 30.600 ;
        RECT 211.350 28.800 213.150 29.550 ;
        RECT 214.650 28.800 216.450 30.600 ;
        RECT 217.950 29.400 220.050 31.500 ;
        RECT 223.050 29.400 224.850 35.250 ;
        RECT 205.050 27.900 205.950 28.200 ;
        RECT 215.100 27.900 216.150 28.800 ;
        RECT 191.550 25.050 196.050 27.150 ;
        RECT 205.050 27.000 216.150 27.900 ;
        RECT 191.550 15.600 192.750 25.050 ;
        RECT 193.950 23.250 197.850 25.050 ;
        RECT 193.950 22.950 196.050 23.250 ;
        RECT 205.050 22.950 205.950 27.000 ;
        RECT 215.100 25.800 216.150 27.000 ;
        RECT 215.100 24.600 222.000 25.800 ;
        RECT 215.100 24.000 216.900 24.600 ;
        RECT 221.100 23.850 222.000 24.600 ;
        RECT 218.100 22.950 219.900 23.700 ;
        RECT 205.050 20.850 208.050 22.950 ;
        RECT 211.950 21.900 219.900 22.950 ;
        RECT 221.100 22.050 222.900 23.850 ;
        RECT 211.950 20.850 214.050 21.900 ;
        RECT 193.950 17.400 195.750 19.200 ;
        RECT 194.850 16.200 199.050 17.400 ;
        RECT 205.050 16.200 205.950 20.850 ;
        RECT 213.750 17.100 215.550 17.400 ;
        RECT 191.550 3.750 193.350 15.600 ;
        RECT 196.950 15.300 199.050 16.200 ;
        RECT 199.950 15.300 205.950 16.200 ;
        RECT 207.150 16.800 215.550 17.100 ;
        RECT 223.950 16.800 224.850 29.400 ;
        RECT 260.850 28.200 262.650 35.250 ;
        RECT 265.350 29.400 267.150 35.250 ;
        RECT 298.650 29.400 300.450 35.250 ;
        RECT 260.850 27.300 264.450 28.200 ;
        RECT 260.100 21.150 261.900 22.950 ;
        RECT 259.950 19.050 262.050 21.150 ;
        RECT 263.250 19.950 264.450 27.300 ;
        RECT 299.250 27.300 300.450 29.400 ;
        RECT 301.650 30.300 303.450 35.250 ;
        RECT 304.650 31.200 306.450 35.250 ;
        RECT 307.650 30.300 309.450 35.250 ;
        RECT 301.650 28.950 309.450 30.300 ;
        RECT 312.150 29.400 313.950 35.250 ;
        RECT 315.150 32.400 316.950 35.250 ;
        RECT 319.950 33.300 321.750 35.250 ;
        RECT 318.000 32.400 321.750 33.300 ;
        RECT 324.450 32.400 326.250 35.250 ;
        RECT 327.750 32.400 329.550 35.250 ;
        RECT 331.650 32.400 333.450 35.250 ;
        RECT 335.850 32.400 337.650 35.250 ;
        RECT 340.350 32.400 342.150 35.250 ;
        RECT 318.000 31.500 319.050 32.400 ;
        RECT 316.950 29.400 319.050 31.500 ;
        RECT 327.750 30.600 328.800 32.400 ;
        RECT 299.250 26.250 303.000 27.300 ;
        RECT 301.950 22.950 303.150 26.250 ;
        RECT 305.100 24.150 306.900 25.950 ;
        RECT 266.100 21.150 267.900 22.950 ;
        RECT 262.950 17.850 265.050 19.950 ;
        RECT 265.950 19.050 268.050 21.150 ;
        RECT 301.950 20.850 304.050 22.950 ;
        RECT 304.950 22.050 307.050 24.150 ;
        RECT 307.950 20.850 310.050 22.950 ;
        RECT 298.950 17.850 301.050 19.950 ;
        RECT 207.150 16.200 224.850 16.800 ;
        RECT 199.950 14.400 200.850 15.300 ;
        RECT 198.150 12.600 200.850 14.400 ;
        RECT 201.750 14.100 203.550 14.400 ;
        RECT 207.150 14.100 208.050 16.200 ;
        RECT 213.750 15.600 224.850 16.200 ;
        RECT 201.750 13.200 208.050 14.100 ;
        RECT 208.950 14.700 210.750 15.300 ;
        RECT 208.950 13.500 216.450 14.700 ;
        RECT 201.750 12.600 203.550 13.200 ;
        RECT 215.250 12.600 216.450 13.500 ;
        RECT 196.950 9.600 200.850 11.700 ;
        RECT 205.950 10.500 212.850 12.300 ;
        RECT 215.250 10.500 220.050 12.600 ;
        RECT 194.550 3.750 196.350 6.600 ;
        RECT 199.050 3.750 200.850 9.600 ;
        RECT 203.250 3.750 205.050 9.600 ;
        RECT 207.150 3.750 208.950 10.500 ;
        RECT 215.250 9.600 216.450 10.500 ;
        RECT 210.150 3.750 211.950 9.600 ;
        RECT 214.950 3.750 216.750 9.600 ;
        RECT 220.050 3.750 221.850 9.600 ;
        RECT 223.050 3.750 224.850 15.600 ;
        RECT 263.250 9.600 264.450 17.850 ;
        RECT 299.250 16.050 301.050 17.850 ;
        RECT 302.850 15.600 304.050 20.850 ;
        RECT 308.100 19.050 309.900 20.850 ;
        RECT 312.150 16.800 313.050 29.400 ;
        RECT 320.550 28.800 322.350 30.600 ;
        RECT 323.850 29.550 328.800 30.600 ;
        RECT 336.300 31.500 337.350 32.400 ;
        RECT 336.300 30.300 340.050 31.500 ;
        RECT 323.850 28.800 325.650 29.550 ;
        RECT 320.850 27.900 321.900 28.800 ;
        RECT 331.050 28.200 332.850 30.000 ;
        RECT 337.950 29.400 340.050 30.300 ;
        RECT 343.650 29.400 345.450 35.250 ;
        RECT 331.050 27.900 331.950 28.200 ;
        RECT 320.850 27.000 331.950 27.900 ;
        RECT 344.250 27.150 345.450 29.400 ;
        RECT 380.850 28.200 382.650 35.250 ;
        RECT 385.350 29.400 387.150 35.250 ;
        RECT 418.650 29.400 420.450 35.250 ;
        RECT 380.850 27.300 384.450 28.200 ;
        RECT 320.850 25.800 321.900 27.000 ;
        RECT 315.000 24.600 321.900 25.800 ;
        RECT 315.000 23.850 315.900 24.600 ;
        RECT 320.100 24.000 321.900 24.600 ;
        RECT 314.100 22.050 315.900 23.850 ;
        RECT 317.100 22.950 318.900 23.700 ;
        RECT 331.050 22.950 331.950 27.000 ;
        RECT 340.950 25.050 345.450 27.150 ;
        RECT 339.150 23.250 343.050 25.050 ;
        RECT 340.950 22.950 343.050 23.250 ;
        RECT 317.100 21.900 325.050 22.950 ;
        RECT 322.950 20.850 325.050 21.900 ;
        RECT 328.950 20.850 331.950 22.950 ;
        RECT 321.450 17.100 323.250 17.400 ;
        RECT 321.450 16.800 329.850 17.100 ;
        RECT 312.150 16.200 329.850 16.800 ;
        RECT 312.150 15.600 323.250 16.200 ;
        RECT 259.650 3.750 261.450 9.600 ;
        RECT 262.650 3.750 264.450 9.600 ;
        RECT 265.650 3.750 267.450 9.600 ;
        RECT 299.400 3.750 301.200 9.600 ;
        RECT 302.700 3.750 304.500 15.600 ;
        RECT 306.900 3.750 308.700 15.600 ;
        RECT 312.150 3.750 313.950 15.600 ;
        RECT 326.250 14.700 328.050 15.300 ;
        RECT 320.550 13.500 328.050 14.700 ;
        RECT 328.950 14.100 329.850 16.200 ;
        RECT 331.050 16.200 331.950 20.850 ;
        RECT 341.250 17.400 343.050 19.200 ;
        RECT 337.950 16.200 342.150 17.400 ;
        RECT 331.050 15.300 337.050 16.200 ;
        RECT 337.950 15.300 340.050 16.200 ;
        RECT 344.250 15.600 345.450 25.050 ;
        RECT 380.100 21.150 381.900 22.950 ;
        RECT 379.950 19.050 382.050 21.150 ;
        RECT 383.250 19.950 384.450 27.300 ;
        RECT 419.250 27.300 420.450 29.400 ;
        RECT 421.650 30.300 423.450 35.250 ;
        RECT 424.650 31.200 426.450 35.250 ;
        RECT 427.650 30.300 429.450 35.250 ;
        RECT 421.650 28.950 429.450 30.300 ;
        RECT 464.850 28.200 466.650 35.250 ;
        RECT 469.350 29.400 471.150 35.250 ;
        RECT 505.650 29.400 507.450 35.250 ;
        RECT 464.850 27.300 468.450 28.200 ;
        RECT 419.250 26.250 423.000 27.300 ;
        RECT 421.950 22.950 423.150 26.250 ;
        RECT 425.100 24.150 426.900 25.950 ;
        RECT 386.100 21.150 387.900 22.950 ;
        RECT 382.950 17.850 385.050 19.950 ;
        RECT 385.950 19.050 388.050 21.150 ;
        RECT 421.950 20.850 424.050 22.950 ;
        RECT 424.950 22.050 427.050 24.150 ;
        RECT 427.950 20.850 430.050 22.950 ;
        RECT 464.100 21.150 465.900 22.950 ;
        RECT 418.950 17.850 421.050 19.950 ;
        RECT 336.150 14.400 337.050 15.300 ;
        RECT 333.450 14.100 335.250 14.400 ;
        RECT 320.550 12.600 321.750 13.500 ;
        RECT 328.950 13.200 335.250 14.100 ;
        RECT 333.450 12.600 335.250 13.200 ;
        RECT 336.150 12.600 338.850 14.400 ;
        RECT 316.950 10.500 321.750 12.600 ;
        RECT 324.150 10.500 331.050 12.300 ;
        RECT 320.550 9.600 321.750 10.500 ;
        RECT 315.150 3.750 316.950 9.600 ;
        RECT 320.250 3.750 322.050 9.600 ;
        RECT 325.050 3.750 326.850 9.600 ;
        RECT 328.050 3.750 329.850 10.500 ;
        RECT 336.150 9.600 340.050 11.700 ;
        RECT 331.950 3.750 333.750 9.600 ;
        RECT 336.150 3.750 337.950 9.600 ;
        RECT 340.650 3.750 342.450 6.600 ;
        RECT 343.650 3.750 345.450 15.600 ;
        RECT 383.250 9.600 384.450 17.850 ;
        RECT 419.250 16.050 421.050 17.850 ;
        RECT 422.850 15.600 424.050 20.850 ;
        RECT 428.100 19.050 429.900 20.850 ;
        RECT 463.950 19.050 466.050 21.150 ;
        RECT 467.250 19.950 468.450 27.300 ;
        RECT 506.250 27.300 507.450 29.400 ;
        RECT 508.650 30.300 510.450 35.250 ;
        RECT 511.650 31.200 513.450 35.250 ;
        RECT 514.650 30.300 516.450 35.250 ;
        RECT 508.650 28.950 516.450 30.300 ;
        RECT 551.850 28.200 553.650 35.250 ;
        RECT 556.350 29.400 558.150 35.250 ;
        RECT 592.650 29.400 594.450 35.250 ;
        RECT 551.850 27.300 555.450 28.200 ;
        RECT 506.250 26.250 510.000 27.300 ;
        RECT 508.950 22.950 510.150 26.250 ;
        RECT 512.100 24.150 513.900 25.950 ;
        RECT 470.100 21.150 471.900 22.950 ;
        RECT 466.950 17.850 469.050 19.950 ;
        RECT 469.950 19.050 472.050 21.150 ;
        RECT 508.950 20.850 511.050 22.950 ;
        RECT 511.950 22.050 514.050 24.150 ;
        RECT 514.950 20.850 517.050 22.950 ;
        RECT 551.100 21.150 552.900 22.950 ;
        RECT 505.950 17.850 508.050 19.950 ;
        RECT 379.650 3.750 381.450 9.600 ;
        RECT 382.650 3.750 384.450 9.600 ;
        RECT 385.650 3.750 387.450 9.600 ;
        RECT 419.400 3.750 421.200 9.600 ;
        RECT 422.700 3.750 424.500 15.600 ;
        RECT 426.900 3.750 428.700 15.600 ;
        RECT 467.250 9.600 468.450 17.850 ;
        RECT 506.250 16.050 508.050 17.850 ;
        RECT 509.850 15.600 511.050 20.850 ;
        RECT 515.100 19.050 516.900 20.850 ;
        RECT 550.950 19.050 553.050 21.150 ;
        RECT 554.250 19.950 555.450 27.300 ;
        RECT 593.250 27.300 594.450 29.400 ;
        RECT 595.650 30.300 597.450 35.250 ;
        RECT 598.650 31.200 600.450 35.250 ;
        RECT 601.650 30.300 603.450 35.250 ;
        RECT 595.650 28.950 603.450 30.300 ;
        RECT 606.150 29.400 607.950 35.250 ;
        RECT 609.150 32.400 610.950 35.250 ;
        RECT 613.950 33.300 615.750 35.250 ;
        RECT 612.000 32.400 615.750 33.300 ;
        RECT 618.450 32.400 620.250 35.250 ;
        RECT 621.750 32.400 623.550 35.250 ;
        RECT 625.650 32.400 627.450 35.250 ;
        RECT 629.850 32.400 631.650 35.250 ;
        RECT 634.350 32.400 636.150 35.250 ;
        RECT 612.000 31.500 613.050 32.400 ;
        RECT 610.950 29.400 613.050 31.500 ;
        RECT 621.750 30.600 622.800 32.400 ;
        RECT 593.250 26.250 597.000 27.300 ;
        RECT 595.950 22.950 597.150 26.250 ;
        RECT 599.100 24.150 600.900 25.950 ;
        RECT 557.100 21.150 558.900 22.950 ;
        RECT 553.950 17.850 556.050 19.950 ;
        RECT 556.950 19.050 559.050 21.150 ;
        RECT 595.950 20.850 598.050 22.950 ;
        RECT 598.950 22.050 601.050 24.150 ;
        RECT 601.950 20.850 604.050 22.950 ;
        RECT 592.950 17.850 595.050 19.950 ;
        RECT 463.650 3.750 465.450 9.600 ;
        RECT 466.650 3.750 468.450 9.600 ;
        RECT 469.650 3.750 471.450 9.600 ;
        RECT 506.400 3.750 508.200 9.600 ;
        RECT 509.700 3.750 511.500 15.600 ;
        RECT 513.900 3.750 515.700 15.600 ;
        RECT 554.250 9.600 555.450 17.850 ;
        RECT 593.250 16.050 595.050 17.850 ;
        RECT 596.850 15.600 598.050 20.850 ;
        RECT 602.100 19.050 603.900 20.850 ;
        RECT 606.150 16.800 607.050 29.400 ;
        RECT 614.550 28.800 616.350 30.600 ;
        RECT 617.850 29.550 622.800 30.600 ;
        RECT 630.300 31.500 631.350 32.400 ;
        RECT 630.300 30.300 634.050 31.500 ;
        RECT 617.850 28.800 619.650 29.550 ;
        RECT 614.850 27.900 615.900 28.800 ;
        RECT 625.050 28.200 626.850 30.000 ;
        RECT 631.950 29.400 634.050 30.300 ;
        RECT 637.650 29.400 639.450 35.250 ;
        RECT 671.550 32.400 673.350 35.250 ;
        RECT 674.550 32.400 676.350 35.250 ;
        RECT 625.050 27.900 625.950 28.200 ;
        RECT 614.850 27.000 625.950 27.900 ;
        RECT 638.250 27.150 639.450 29.400 ;
        RECT 614.850 25.800 615.900 27.000 ;
        RECT 609.000 24.600 615.900 25.800 ;
        RECT 609.000 23.850 609.900 24.600 ;
        RECT 614.100 24.000 615.900 24.600 ;
        RECT 608.100 22.050 609.900 23.850 ;
        RECT 611.100 22.950 612.900 23.700 ;
        RECT 625.050 22.950 625.950 27.000 ;
        RECT 634.950 25.050 639.450 27.150 ;
        RECT 633.150 23.250 637.050 25.050 ;
        RECT 634.950 22.950 637.050 23.250 ;
        RECT 611.100 21.900 619.050 22.950 ;
        RECT 616.950 20.850 619.050 21.900 ;
        RECT 622.950 20.850 625.950 22.950 ;
        RECT 615.450 17.100 617.250 17.400 ;
        RECT 615.450 16.800 623.850 17.100 ;
        RECT 606.150 16.200 623.850 16.800 ;
        RECT 606.150 15.600 617.250 16.200 ;
        RECT 550.650 3.750 552.450 9.600 ;
        RECT 553.650 3.750 555.450 9.600 ;
        RECT 556.650 3.750 558.450 9.600 ;
        RECT 593.400 3.750 595.200 9.600 ;
        RECT 596.700 3.750 598.500 15.600 ;
        RECT 600.900 3.750 602.700 15.600 ;
        RECT 606.150 3.750 607.950 15.600 ;
        RECT 620.250 14.700 622.050 15.300 ;
        RECT 614.550 13.500 622.050 14.700 ;
        RECT 622.950 14.100 623.850 16.200 ;
        RECT 625.050 16.200 625.950 20.850 ;
        RECT 635.250 17.400 637.050 19.200 ;
        RECT 631.950 16.200 636.150 17.400 ;
        RECT 625.050 15.300 631.050 16.200 ;
        RECT 631.950 15.300 634.050 16.200 ;
        RECT 638.250 15.600 639.450 25.050 ;
        RECT 670.950 23.850 673.050 25.950 ;
        RECT 674.400 24.150 675.600 32.400 ;
        RECT 713.850 28.200 715.650 35.250 ;
        RECT 718.350 29.400 720.150 35.250 ;
        RECT 749.850 29.400 751.650 35.250 ;
        RECT 754.350 28.200 756.150 35.250 ;
        RECT 713.850 27.300 717.450 28.200 ;
        RECT 671.100 22.050 672.900 23.850 ;
        RECT 673.950 22.050 676.050 24.150 ;
        RECT 630.150 14.400 631.050 15.300 ;
        RECT 627.450 14.100 629.250 14.400 ;
        RECT 614.550 12.600 615.750 13.500 ;
        RECT 622.950 13.200 629.250 14.100 ;
        RECT 627.450 12.600 629.250 13.200 ;
        RECT 630.150 12.600 632.850 14.400 ;
        RECT 610.950 10.500 615.750 12.600 ;
        RECT 618.150 10.500 625.050 12.300 ;
        RECT 614.550 9.600 615.750 10.500 ;
        RECT 609.150 3.750 610.950 9.600 ;
        RECT 614.250 3.750 616.050 9.600 ;
        RECT 619.050 3.750 620.850 9.600 ;
        RECT 622.050 3.750 623.850 10.500 ;
        RECT 630.150 9.600 634.050 11.700 ;
        RECT 625.950 3.750 627.750 9.600 ;
        RECT 630.150 3.750 631.950 9.600 ;
        RECT 634.650 3.750 636.450 6.600 ;
        RECT 637.650 3.750 639.450 15.600 ;
        RECT 674.400 9.600 675.600 22.050 ;
        RECT 713.100 21.150 714.900 22.950 ;
        RECT 712.950 19.050 715.050 21.150 ;
        RECT 716.250 19.950 717.450 27.300 ;
        RECT 752.550 27.300 756.150 28.200 ;
        RECT 719.100 21.150 720.900 22.950 ;
        RECT 749.100 21.150 750.900 22.950 ;
        RECT 715.950 17.850 718.050 19.950 ;
        RECT 718.950 19.050 721.050 21.150 ;
        RECT 748.950 19.050 751.050 21.150 ;
        RECT 752.550 19.950 753.750 27.300 ;
        RECT 755.100 21.150 756.900 22.950 ;
        RECT 751.950 17.850 754.050 19.950 ;
        RECT 754.950 19.050 757.050 21.150 ;
        RECT 716.250 9.600 717.450 17.850 ;
        RECT 752.550 9.600 753.750 17.850 ;
        RECT 671.550 3.750 673.350 9.600 ;
        RECT 674.550 3.750 676.350 9.600 ;
        RECT 712.650 3.750 714.450 9.600 ;
        RECT 715.650 3.750 717.450 9.600 ;
        RECT 718.650 3.750 720.450 9.600 ;
        RECT 749.550 3.750 751.350 9.600 ;
        RECT 752.550 3.750 754.350 9.600 ;
        RECT 755.550 3.750 757.350 9.600 ;
      LAYER metal2 ;
        RECT 91.950 749.400 94.050 751.500 ;
        RECT 112.950 749.400 115.050 751.500 ;
        RECT 169.950 749.400 172.050 751.500 ;
        RECT 190.950 749.400 193.050 751.500 ;
        RECT 457.950 749.400 460.050 751.500 ;
        RECT 478.950 749.400 481.050 751.500 ;
        RECT 535.950 749.400 538.050 751.500 ;
        RECT 556.950 749.400 559.050 751.500 ;
        RECT 76.950 742.950 79.050 745.050 ;
        RECT 82.950 744.450 85.050 745.050 ;
        RECT 80.250 743.250 81.750 744.150 ;
        RECT 82.950 743.400 87.450 744.450 ;
        RECT 82.950 742.950 85.050 743.400 ;
        RECT 28.950 740.250 30.750 741.150 ;
        RECT 31.950 739.950 34.050 742.050 ;
        RECT 35.250 740.250 37.050 741.150 ;
        RECT 73.950 739.950 76.050 742.050 ;
        RECT 77.250 740.850 78.750 741.750 ;
        RECT 79.950 739.950 82.050 742.050 ;
        RECT 83.250 740.850 85.050 741.750 ;
        RECT 32.250 737.850 33.750 738.750 ;
        RECT 34.950 736.950 37.050 739.050 ;
        RECT 73.950 737.850 76.050 738.750 ;
        RECT 80.400 736.050 81.450 739.950 ;
        RECT 86.400 739.050 87.450 743.400 ;
        RECT 85.950 736.950 88.050 739.050 ;
        RECT 34.950 733.950 37.050 736.050 ;
        RECT 79.950 733.950 82.050 736.050 ;
        RECT 86.400 735.450 87.450 736.950 ;
        RECT 86.400 734.400 90.450 735.450 ;
        RECT 35.400 703.050 36.450 733.950 ;
        RECT 76.950 706.950 79.050 709.050 ;
        RECT 82.950 707.250 85.050 708.150 ;
        RECT 77.400 706.050 78.450 706.950 ;
        RECT 76.950 703.950 79.050 706.050 ;
        RECT 80.250 704.250 81.750 705.150 ;
        RECT 82.950 703.950 85.050 706.050 ;
        RECT 86.250 704.250 88.050 705.150 ;
        RECT 34.950 700.950 37.050 703.050 ;
        RECT 40.950 702.450 43.050 703.050 ;
        RECT 40.950 701.400 45.450 702.450 ;
        RECT 76.950 701.850 78.750 702.750 ;
        RECT 40.950 700.950 43.050 701.400 ;
        RECT 34.950 698.850 37.050 699.750 ;
        RECT 40.950 698.850 43.050 699.750 ;
        RECT 37.950 673.950 40.050 676.050 ;
        RECT 34.950 671.250 37.050 672.150 ;
        RECT 37.950 671.850 40.050 672.750 ;
        RECT 34.950 667.950 37.050 670.050 ;
        RECT 35.400 667.050 36.450 667.950 ;
        RECT 34.950 664.950 37.050 667.050 ;
        RECT 44.400 637.050 45.450 701.400 ;
        RECT 79.950 700.950 82.050 703.050 ;
        RECT 80.400 693.450 81.450 700.950 ;
        RECT 83.400 697.050 84.450 703.950 ;
        RECT 85.950 700.950 88.050 703.050 ;
        RECT 86.400 700.050 87.450 700.950 ;
        RECT 89.400 700.050 90.450 734.400 ;
        RECT 92.400 732.600 93.600 749.400 ;
        RECT 103.950 745.950 106.050 748.050 ;
        RECT 104.400 745.050 105.450 745.950 ;
        RECT 97.950 742.950 100.050 745.050 ;
        RECT 103.950 744.450 106.050 745.050 ;
        RECT 101.400 743.400 106.050 744.450 ;
        RECT 97.950 740.850 100.050 741.750 ;
        RECT 91.950 730.500 94.050 732.600 ;
        RECT 85.950 697.950 88.050 700.050 ;
        RECT 88.950 697.950 91.050 700.050 ;
        RECT 82.950 694.950 85.050 697.050 ;
        RECT 80.400 692.400 84.450 693.450 ;
        RECT 46.950 673.950 49.050 676.050 ;
        RECT 47.400 670.050 48.450 673.950 ;
        RECT 64.950 670.950 67.050 673.050 ;
        RECT 73.950 670.950 76.050 673.050 ;
        RECT 76.950 670.950 79.050 673.050 ;
        RECT 46.950 667.950 49.050 670.050 ;
        RECT 37.950 634.950 40.050 637.050 ;
        RECT 43.950 634.950 46.050 637.050 ;
        RECT 38.400 634.050 39.450 634.950 ;
        RECT 31.950 631.950 34.050 634.050 ;
        RECT 35.250 632.250 36.750 633.150 ;
        RECT 37.950 631.950 40.050 634.050 ;
        RECT 40.950 631.950 43.050 634.050 ;
        RECT 31.950 629.850 33.750 630.750 ;
        RECT 34.950 628.950 37.050 631.050 ;
        RECT 38.250 629.850 40.050 630.750 ;
        RECT 41.400 607.050 42.450 631.950 ;
        RECT 40.950 604.950 43.050 607.050 ;
        RECT 37.950 601.950 40.050 604.050 ;
        RECT 41.400 601.050 42.450 604.950 ;
        RECT 47.400 601.050 48.450 667.950 ;
        RECT 65.400 631.050 66.450 670.950 ;
        RECT 70.950 669.450 73.050 670.050 ;
        RECT 68.400 668.400 73.050 669.450 ;
        RECT 68.400 667.050 69.450 668.400 ;
        RECT 70.950 667.950 73.050 668.400 ;
        RECT 74.400 667.050 75.450 670.950 ;
        RECT 77.400 670.050 78.450 670.950 ;
        RECT 76.950 667.950 79.050 670.050 ;
        RECT 80.250 668.250 82.050 669.150 ;
        RECT 67.950 664.950 70.050 667.050 ;
        RECT 70.950 665.850 72.750 666.750 ;
        RECT 73.950 664.950 76.050 667.050 ;
        RECT 77.250 665.850 78.750 666.750 ;
        RECT 79.950 666.450 82.050 667.050 ;
        RECT 83.400 666.450 84.450 692.400 ;
        RECT 85.950 670.950 88.050 673.050 ;
        RECT 86.400 667.050 87.450 670.950 ;
        RECT 79.950 665.400 84.450 666.450 ;
        RECT 79.950 664.950 82.050 665.400 ;
        RECT 85.950 664.950 88.050 667.050 ;
        RECT 73.950 662.850 76.050 663.750 ;
        RECT 79.950 634.950 82.050 637.050 ;
        RECT 80.400 634.050 81.450 634.950 ;
        RECT 73.950 631.950 76.050 634.050 ;
        RECT 77.250 632.250 78.750 633.150 ;
        RECT 79.950 631.950 82.050 634.050 ;
        RECT 86.400 631.050 87.450 664.950 ;
        RECT 64.950 628.950 67.050 631.050 ;
        RECT 73.950 629.850 75.750 630.750 ;
        RECT 76.950 628.950 79.050 631.050 ;
        RECT 80.250 629.850 82.050 630.750 ;
        RECT 85.950 628.950 88.050 631.050 ;
        RECT 76.950 604.950 79.050 607.050 ;
        RECT 79.950 604.950 82.050 607.050 ;
        RECT 85.950 605.400 88.050 607.500 ;
        RECT 77.400 604.050 78.450 604.950 ;
        RECT 76.950 601.950 79.050 604.050 ;
        RECT 34.950 598.950 37.050 601.050 ;
        RECT 38.250 599.850 39.750 600.750 ;
        RECT 40.950 598.950 43.050 601.050 ;
        RECT 46.950 598.950 49.050 601.050 ;
        RECT 73.950 599.250 76.050 600.150 ;
        RECT 76.950 599.850 79.050 600.750 ;
        RECT 34.950 596.850 37.050 597.750 ;
        RECT 40.950 596.850 43.050 597.750 ;
        RECT 34.950 560.250 37.050 561.150 ;
        RECT 40.950 559.950 43.050 562.050 ;
        RECT 41.400 559.050 42.450 559.950 ;
        RECT 34.950 556.950 37.050 559.050 ;
        RECT 38.250 557.250 39.750 558.150 ;
        RECT 40.950 556.950 43.050 559.050 ;
        RECT 44.250 557.250 46.050 558.150 ;
        RECT 37.950 553.950 40.050 556.050 ;
        RECT 41.250 554.850 42.750 555.750 ;
        RECT 43.950 553.950 46.050 556.050 ;
        RECT 38.400 541.050 39.450 553.950 ;
        RECT 13.950 538.950 16.050 541.050 ;
        RECT 37.950 538.950 40.050 541.050 ;
        RECT 7.950 533.400 10.050 535.500 ;
        RECT 8.400 516.600 9.600 533.400 ;
        RECT 14.400 529.050 15.450 538.950 ;
        RECT 28.950 533.400 31.050 535.500 ;
        RECT 22.950 529.950 25.050 532.050 ;
        RECT 13.950 526.950 16.050 529.050 ;
        RECT 19.950 528.450 22.050 529.050 ;
        RECT 23.400 528.450 24.450 529.950 ;
        RECT 19.950 527.400 24.450 528.450 ;
        RECT 19.950 526.950 22.050 527.400 ;
        RECT 13.950 524.850 16.050 525.750 ;
        RECT 19.950 524.850 22.050 525.750 ;
        RECT 7.950 514.500 10.050 516.600 ;
        RECT 7.950 494.400 10.050 496.500 ;
        RECT 8.400 477.600 9.600 494.400 ;
        RECT 13.950 485.250 16.050 486.150 ;
        RECT 19.950 485.250 22.050 486.150 ;
        RECT 13.950 481.950 16.050 484.050 ;
        RECT 19.950 481.950 22.050 484.050 ;
        RECT 14.400 481.050 15.450 481.950 ;
        RECT 13.950 478.950 16.050 481.050 ;
        RECT 7.950 475.500 10.050 477.600 ;
        RECT 20.400 475.050 21.450 481.950 ;
        RECT 23.400 475.050 24.450 527.400 ;
        RECT 29.250 521.400 30.450 533.400 ;
        RECT 31.950 530.250 34.050 531.150 ;
        RECT 31.950 526.950 34.050 529.050 ;
        RECT 28.950 519.300 31.050 521.400 ;
        RECT 47.400 520.050 48.450 598.950 ;
        RECT 73.950 595.950 76.050 598.050 ;
        RECT 80.400 564.450 81.450 604.950 ;
        RECT 86.400 588.600 87.600 605.400 ;
        RECT 91.950 600.450 94.050 601.050 ;
        RECT 97.950 600.450 100.050 601.050 ;
        RECT 101.400 600.450 102.450 743.400 ;
        RECT 103.950 742.950 106.050 743.400 ;
        RECT 103.950 740.850 106.050 741.750 ;
        RECT 113.250 737.400 114.450 749.400 ;
        RECT 115.950 746.250 118.050 747.150 ;
        RECT 115.950 742.950 118.050 745.050 ;
        RECT 154.950 742.950 157.050 745.050 ;
        RECT 160.950 744.450 163.050 745.050 ;
        RECT 158.250 743.250 159.750 744.150 ;
        RECT 160.950 743.400 165.450 744.450 ;
        RECT 160.950 742.950 163.050 743.400 ;
        RECT 112.950 735.300 115.050 737.400 ;
        RECT 113.250 731.700 114.450 735.300 ;
        RECT 112.950 729.600 115.050 731.700 ;
        RECT 116.400 706.050 117.450 742.950 ;
        RECT 164.400 742.050 165.450 743.400 ;
        RECT 127.950 739.950 130.050 742.050 ;
        RECT 151.950 739.950 154.050 742.050 ;
        RECT 155.250 740.850 156.750 741.750 ;
        RECT 157.950 739.950 160.050 742.050 ;
        RECT 161.250 740.850 163.050 741.750 ;
        RECT 163.950 739.950 166.050 742.050 ;
        RECT 121.950 707.250 124.050 708.150 ;
        RECT 128.400 706.050 129.450 739.950 ;
        RECT 151.950 737.850 154.050 738.750 ;
        RECT 115.950 703.950 118.050 706.050 ;
        RECT 118.950 704.250 120.750 705.150 ;
        RECT 121.950 703.950 124.050 706.050 ;
        RECT 125.250 704.250 126.750 705.150 ;
        RECT 127.950 703.950 130.050 706.050 ;
        RECT 122.400 703.050 123.450 703.950 ;
        RECT 115.950 700.950 118.050 703.050 ;
        RECT 118.950 700.950 121.050 703.050 ;
        RECT 121.950 700.950 124.050 703.050 ;
        RECT 124.950 700.950 127.050 703.050 ;
        RECT 128.250 701.850 130.050 702.750 ;
        RECT 109.950 673.950 112.050 676.050 ;
        RECT 110.400 637.050 111.450 673.950 ;
        RECT 116.400 664.050 117.450 700.950 ;
        RECT 119.400 700.050 120.450 700.950 ;
        RECT 118.950 697.950 121.050 700.050 ;
        RECT 125.400 696.450 126.450 700.950 ;
        RECT 158.400 700.050 159.450 739.950 ;
        RECT 170.400 732.600 171.600 749.400 ;
        RECT 181.950 745.950 184.050 748.050 ;
        RECT 182.400 745.050 183.450 745.950 ;
        RECT 175.950 742.950 178.050 745.050 ;
        RECT 181.950 742.950 184.050 745.050 ;
        RECT 175.950 740.850 178.050 741.750 ;
        RECT 181.950 740.850 184.050 741.750 ;
        RECT 191.250 737.400 192.450 749.400 ;
        RECT 193.950 746.250 196.050 747.150 ;
        RECT 196.950 745.950 199.050 748.050 ;
        RECT 229.950 745.950 232.050 748.050 ;
        RECT 268.950 745.950 271.050 748.050 ;
        RECT 283.950 745.950 286.050 748.050 ;
        RECT 193.950 744.450 196.050 745.050 ;
        RECT 197.400 744.450 198.450 745.950 ;
        RECT 193.950 743.400 198.450 744.450 ;
        RECT 229.950 743.850 232.050 744.750 ;
        RECT 193.950 742.950 196.050 743.400 ;
        RECT 232.950 743.250 235.050 744.150 ;
        RECT 268.950 743.850 270.750 744.750 ;
        RECT 271.950 742.950 274.050 745.050 ;
        RECT 277.950 743.250 280.050 744.150 ;
        RECT 232.950 739.950 235.050 742.050 ;
        RECT 235.950 739.950 238.050 742.050 ;
        RECT 271.950 740.850 274.050 741.750 ;
        RECT 277.950 739.950 280.050 742.050 ;
        RECT 190.950 735.300 193.050 737.400 ;
        RECT 169.950 730.500 172.050 732.600 ;
        RECT 191.250 731.700 192.450 735.300 ;
        RECT 190.950 729.600 193.050 731.700 ;
        RECT 220.950 703.950 223.050 706.050 ;
        RECT 166.950 701.250 169.050 702.150 ;
        RECT 172.950 701.250 175.050 702.150 ;
        RECT 208.950 700.950 211.050 703.050 ;
        RECT 157.950 697.950 160.050 700.050 ;
        RECT 166.950 697.950 169.050 700.050 ;
        RECT 172.950 697.950 175.050 700.050 ;
        RECT 208.950 698.850 211.050 699.750 ;
        RECT 211.950 698.250 214.050 699.150 ;
        RECT 122.400 695.400 126.450 696.450 ;
        RECT 122.400 670.050 123.450 695.400 ;
        RECT 169.950 694.950 172.050 697.050 ;
        RECT 157.950 673.950 160.050 676.050 ;
        RECT 154.950 670.950 157.050 673.050 ;
        RECT 118.950 668.250 120.750 669.150 ;
        RECT 121.950 667.950 124.050 670.050 ;
        RECT 125.250 668.250 127.050 669.150 ;
        RECT 118.950 664.950 121.050 667.050 ;
        RECT 122.250 665.850 123.750 666.750 ;
        RECT 124.950 664.950 127.050 667.050 ;
        RECT 115.950 661.950 118.050 664.050 ;
        RECT 121.950 661.950 124.050 664.050 ;
        RECT 109.950 634.950 112.050 637.050 ;
        RECT 115.950 635.250 118.050 636.150 ;
        RECT 110.400 630.450 111.450 634.950 ;
        RECT 122.400 634.050 123.450 661.950 ;
        RECT 112.950 632.250 114.750 633.150 ;
        RECT 115.950 631.950 118.050 634.050 ;
        RECT 119.250 632.250 120.750 633.150 ;
        RECT 121.950 631.950 124.050 634.050 ;
        RECT 112.950 630.450 115.050 631.050 ;
        RECT 110.400 629.400 115.050 630.450 ;
        RECT 112.950 628.950 115.050 629.400 ;
        RECT 106.950 605.400 109.050 607.500 ;
        RECT 116.400 607.050 117.450 631.950 ;
        RECT 118.950 628.950 121.050 631.050 ;
        RECT 122.250 629.850 124.050 630.750 ;
        RECT 91.950 599.400 96.450 600.450 ;
        RECT 91.950 598.950 94.050 599.400 ;
        RECT 91.950 596.850 94.050 597.750 ;
        RECT 85.950 586.500 88.050 588.600 ;
        RECT 77.400 563.400 81.450 564.450 ;
        RECT 77.400 562.050 78.450 563.400 ;
        RECT 64.950 559.950 67.050 562.050 ;
        RECT 76.950 561.450 79.050 562.050 ;
        RECT 74.400 560.400 79.050 561.450 ;
        RECT 29.250 515.700 30.450 519.300 ;
        RECT 31.950 517.950 34.050 520.050 ;
        RECT 46.950 517.950 49.050 520.050 ;
        RECT 28.950 513.600 31.050 515.700 ;
        RECT 28.950 495.300 31.050 497.400 ;
        RECT 29.250 491.700 30.450 495.300 ;
        RECT 28.950 489.600 31.050 491.700 ;
        RECT 29.250 477.600 30.450 489.600 ;
        RECT 32.400 484.050 33.450 517.950 ;
        RECT 65.400 517.050 66.450 559.950 ;
        RECT 74.400 529.050 75.450 560.400 ;
        RECT 76.950 559.950 79.050 560.400 ;
        RECT 80.250 560.250 81.750 561.150 ;
        RECT 82.950 559.950 85.050 562.050 ;
        RECT 76.950 557.850 78.750 558.750 ;
        RECT 79.950 556.950 82.050 559.050 ;
        RECT 83.250 557.850 85.050 558.750 ;
        RECT 95.400 553.050 96.450 599.400 ;
        RECT 97.950 599.400 102.450 600.450 ;
        RECT 97.950 598.950 100.050 599.400 ;
        RECT 97.950 596.850 100.050 597.750 ;
        RECT 94.950 550.950 97.050 553.050 ;
        RECT 85.950 533.400 88.050 535.500 ;
        RECT 73.950 526.950 76.050 529.050 ;
        RECT 67.950 524.250 69.750 525.150 ;
        RECT 70.950 523.950 73.050 526.050 ;
        RECT 74.250 524.250 76.050 525.150 ;
        RECT 76.950 523.950 79.050 526.050 ;
        RECT 67.950 520.950 70.050 523.050 ;
        RECT 71.250 521.850 72.750 522.750 ;
        RECT 73.950 520.950 76.050 523.050 ;
        RECT 68.400 520.050 69.450 520.950 ;
        RECT 67.950 517.950 70.050 520.050 ;
        RECT 74.400 517.050 75.450 520.950 ;
        RECT 64.950 514.950 67.050 517.050 ;
        RECT 67.950 514.950 70.050 517.050 ;
        RECT 73.950 514.950 76.050 517.050 ;
        RECT 68.400 487.050 69.450 514.950 ;
        RECT 73.950 488.250 76.050 489.150 ;
        RECT 61.950 484.950 64.050 487.050 ;
        RECT 64.950 485.250 66.750 486.150 ;
        RECT 67.950 484.950 70.050 487.050 ;
        RECT 73.950 486.450 76.050 487.050 ;
        RECT 77.400 486.450 78.450 523.950 ;
        RECT 86.400 516.600 87.600 533.400 ;
        RECT 101.400 532.050 102.450 599.400 ;
        RECT 107.250 593.400 108.450 605.400 ;
        RECT 115.950 604.950 118.050 607.050 ;
        RECT 109.950 602.250 112.050 603.150 ;
        RECT 109.950 598.950 112.050 601.050 ;
        RECT 106.950 591.300 109.050 593.400 ;
        RECT 107.250 587.700 108.450 591.300 ;
        RECT 106.950 585.600 109.050 587.700 ;
        RECT 110.400 568.050 111.450 598.950 ;
        RECT 125.400 598.050 126.450 664.950 ;
        RECT 155.400 663.450 156.450 670.950 ;
        RECT 158.400 670.050 159.450 673.950 ;
        RECT 163.950 670.950 166.050 673.050 ;
        RECT 164.400 670.050 165.450 670.950 ;
        RECT 157.950 667.950 160.050 670.050 ;
        RECT 160.950 667.950 163.050 670.050 ;
        RECT 163.950 667.950 166.050 670.050 ;
        RECT 167.250 668.250 169.050 669.150 ;
        RECT 161.400 667.050 162.450 667.950 ;
        RECT 157.950 665.850 159.750 666.750 ;
        RECT 160.950 664.950 163.050 667.050 ;
        RECT 164.250 665.850 165.750 666.750 ;
        RECT 166.950 666.450 169.050 667.050 ;
        RECT 170.400 666.450 171.450 694.950 ;
        RECT 173.400 691.050 174.450 697.950 ;
        RECT 211.950 694.950 214.050 697.050 ;
        RECT 172.950 688.950 175.050 691.050 ;
        RECT 212.400 682.050 213.450 694.950 ;
        RECT 211.950 679.950 214.050 682.050 ;
        RECT 205.950 676.950 208.050 679.050 ;
        RECT 206.400 676.050 207.450 676.950 ;
        RECT 221.400 676.050 222.450 703.950 ;
        RECT 232.950 679.950 235.050 682.050 ;
        RECT 205.950 673.950 208.050 676.050 ;
        RECT 220.950 673.950 223.050 676.050 ;
        RECT 206.400 673.050 207.450 673.950 ;
        RECT 221.400 673.050 222.450 673.950 ;
        RECT 205.950 670.950 208.050 673.050 ;
        RECT 211.950 670.950 214.050 673.050 ;
        RECT 220.950 670.950 223.050 673.050 ;
        RECT 205.950 668.850 208.050 669.750 ;
        RECT 211.950 668.850 214.050 669.750 ;
        RECT 166.950 665.400 171.450 666.450 ;
        RECT 166.950 664.950 169.050 665.400 ;
        RECT 155.400 662.400 159.450 663.450 ;
        RECT 160.950 662.850 163.050 663.750 ;
        RECT 151.950 631.950 154.050 634.050 ;
        RECT 148.950 598.950 151.050 601.050 ;
        RECT 124.950 595.950 127.050 598.050 ;
        RECT 145.950 595.950 148.050 598.050 ;
        RECT 149.400 595.050 150.450 598.950 ;
        RECT 152.400 598.050 153.450 631.950 ;
        RECT 151.950 595.950 154.050 598.050 ;
        RECT 155.250 596.250 157.050 597.150 ;
        RECT 145.950 593.850 147.750 594.750 ;
        RECT 148.950 592.950 151.050 595.050 ;
        RECT 152.250 593.850 153.750 594.750 ;
        RECT 154.950 594.450 157.050 595.050 ;
        RECT 158.400 594.450 159.450 662.400 ;
        RECT 169.950 634.950 172.050 637.050 ;
        RECT 208.950 634.950 211.050 637.050 ;
        RECT 160.950 631.950 163.050 634.050 ;
        RECT 166.950 633.450 169.050 634.050 ;
        RECT 170.400 633.450 171.450 634.950 ;
        RECT 209.400 634.050 210.450 634.950 ;
        RECT 164.250 632.250 165.750 633.150 ;
        RECT 166.950 632.400 171.450 633.450 ;
        RECT 166.950 631.950 169.050 632.400 ;
        RECT 160.950 629.850 162.750 630.750 ;
        RECT 163.950 628.950 166.050 631.050 ;
        RECT 167.250 629.850 169.050 630.750 ;
        RECT 170.400 601.050 171.450 632.400 ;
        RECT 190.950 631.950 193.050 634.050 ;
        RECT 202.950 631.950 205.050 634.050 ;
        RECT 206.250 632.250 207.750 633.150 ;
        RECT 208.950 631.950 211.050 634.050 ;
        RECT 191.400 604.050 192.450 631.950 ;
        RECT 202.950 629.850 204.750 630.750 ;
        RECT 205.950 628.950 208.050 631.050 ;
        RECT 209.250 629.850 211.050 630.750 ;
        RECT 190.950 601.950 193.050 604.050 ;
        RECT 169.950 598.950 172.050 601.050 ;
        RECT 184.950 600.450 187.050 601.050 ;
        RECT 187.950 600.450 190.050 601.050 ;
        RECT 184.950 599.400 190.050 600.450 ;
        RECT 184.950 598.950 187.050 599.400 ;
        RECT 187.950 598.950 190.050 599.400 ;
        RECT 154.950 593.400 159.450 594.450 ;
        RECT 154.950 592.950 157.050 593.400 ;
        RECT 148.950 590.850 151.050 591.750 ;
        RECT 109.950 565.950 112.050 568.050 ;
        RECT 160.950 565.950 163.050 568.050 ;
        RECT 121.950 562.950 124.050 565.050 ;
        RECT 122.400 559.050 123.450 562.950 ;
        RECT 161.400 562.050 162.450 565.950 ;
        RECT 166.950 562.950 169.050 565.050 ;
        RECT 167.400 562.050 168.450 562.950 ;
        RECT 127.950 560.250 130.050 561.150 ;
        RECT 160.950 559.950 163.050 562.050 ;
        RECT 164.250 560.250 165.750 561.150 ;
        RECT 166.950 559.950 169.050 562.050 ;
        RECT 112.950 556.950 115.050 559.050 ;
        RECT 118.950 557.250 120.750 558.150 ;
        RECT 121.950 556.950 124.050 559.050 ;
        RECT 125.250 557.250 126.750 558.150 ;
        RECT 127.950 556.950 130.050 559.050 ;
        RECT 160.950 557.850 162.750 558.750 ;
        RECT 163.950 556.950 166.050 559.050 ;
        RECT 167.250 557.850 169.050 558.750 ;
        RECT 106.950 533.400 109.050 535.500 ;
        RECT 97.950 529.950 100.050 532.050 ;
        RECT 100.950 529.950 103.050 532.050 ;
        RECT 98.400 529.050 99.450 529.950 ;
        RECT 91.950 528.450 94.050 529.050 ;
        RECT 91.950 527.400 96.450 528.450 ;
        RECT 91.950 526.950 94.050 527.400 ;
        RECT 91.950 524.850 94.050 525.750 ;
        RECT 85.950 514.500 88.050 516.600 ;
        RECT 71.250 485.250 72.750 486.150 ;
        RECT 73.950 485.400 78.450 486.450 ;
        RECT 73.950 484.950 76.050 485.400 ;
        RECT 31.950 481.950 34.050 484.050 ;
        RECT 31.950 479.850 34.050 480.750 ;
        RECT 28.950 475.500 31.050 477.600 ;
        RECT 19.950 472.950 22.050 475.050 ;
        RECT 22.950 472.950 25.050 475.050 ;
        RECT 52.950 472.950 55.050 475.050 ;
        RECT 34.950 455.250 37.050 456.150 ;
        RECT 53.400 453.450 54.450 472.950 ;
        RECT 55.950 455.250 58.050 456.150 ;
        RECT 55.950 453.450 58.050 454.050 ;
        RECT 53.400 452.400 58.050 453.450 ;
        RECT 55.950 451.950 58.050 452.400 ;
        RECT 7.950 422.400 10.050 424.500 ;
        RECT 28.950 423.300 31.050 425.400 ;
        RECT 8.400 405.600 9.600 422.400 ;
        RECT 29.250 419.700 30.450 423.300 ;
        RECT 43.950 422.400 46.050 424.500 ;
        RECT 28.950 417.600 31.050 419.700 ;
        RECT 13.950 413.250 16.050 414.150 ;
        RECT 19.950 413.250 22.050 414.150 ;
        RECT 13.950 409.950 16.050 412.050 ;
        RECT 19.950 409.950 22.050 412.050 ;
        RECT 22.950 409.950 25.050 412.050 ;
        RECT 7.950 403.500 10.050 405.600 ;
        RECT 14.400 400.050 15.450 409.950 ;
        RECT 20.400 408.450 21.450 409.950 ;
        RECT 23.400 408.450 24.450 409.950 ;
        RECT 20.400 407.400 24.450 408.450 ;
        RECT 13.950 397.950 16.050 400.050 ;
        RECT 7.950 350.400 10.050 352.500 ;
        RECT 8.400 333.600 9.600 350.400 ;
        RECT 13.950 341.250 16.050 342.150 ;
        RECT 19.950 341.250 22.050 342.150 ;
        RECT 19.950 337.950 22.050 340.050 ;
        RECT 7.950 331.500 10.050 333.600 ;
        RECT 7.950 317.400 10.050 319.500 ;
        RECT 8.400 300.600 9.600 317.400 ;
        RECT 20.400 313.050 21.450 337.950 ;
        RECT 13.950 312.450 16.050 313.050 ;
        RECT 19.950 312.450 22.050 313.050 ;
        RECT 23.400 312.450 24.450 407.400 ;
        RECT 29.250 405.600 30.450 417.600 ;
        RECT 31.950 411.450 34.050 412.050 ;
        RECT 31.950 410.400 36.450 411.450 ;
        RECT 31.950 409.950 34.050 410.400 ;
        RECT 31.950 407.850 34.050 408.750 ;
        RECT 28.950 403.500 31.050 405.600 ;
        RECT 35.400 403.050 36.450 410.400 ;
        RECT 44.400 405.600 45.600 422.400 ;
        RECT 49.950 413.250 52.050 414.150 ;
        RECT 55.950 413.250 58.050 414.150 ;
        RECT 49.950 409.950 52.050 412.050 ;
        RECT 55.950 409.950 58.050 412.050 ;
        RECT 43.950 403.500 46.050 405.600 ;
        RECT 34.950 400.950 37.050 403.050 ;
        RECT 50.400 400.050 51.450 409.950 ;
        RECT 56.400 409.050 57.450 409.950 ;
        RECT 55.950 406.950 58.050 409.050 ;
        RECT 37.950 397.950 40.050 400.050 ;
        RECT 49.950 397.950 52.050 400.050 ;
        RECT 38.400 385.050 39.450 397.950 ;
        RECT 43.950 385.950 46.050 388.050 ;
        RECT 44.400 385.050 45.450 385.950 ;
        RECT 34.950 382.950 37.050 385.050 ;
        RECT 37.950 382.950 40.050 385.050 ;
        RECT 41.250 383.250 42.750 384.150 ;
        RECT 43.950 382.950 46.050 385.050 ;
        RECT 46.950 382.950 49.050 385.050 ;
        RECT 35.400 382.050 36.450 382.950 ;
        RECT 34.950 379.950 37.050 382.050 ;
        RECT 38.250 380.850 39.750 381.750 ;
        RECT 40.950 379.950 43.050 382.050 ;
        RECT 44.250 380.850 46.050 381.750 ;
        RECT 34.950 377.850 37.050 378.750 ;
        RECT 28.950 351.300 31.050 353.400 ;
        RECT 29.250 347.700 30.450 351.300 ;
        RECT 28.950 345.600 31.050 347.700 ;
        RECT 29.250 333.600 30.450 345.600 ;
        RECT 31.950 339.450 34.050 340.050 ;
        RECT 31.950 338.400 36.450 339.450 ;
        RECT 31.950 337.950 34.050 338.400 ;
        RECT 35.400 337.050 36.450 338.400 ;
        RECT 31.950 335.850 34.050 336.750 ;
        RECT 34.950 334.950 37.050 337.050 ;
        RECT 28.950 331.500 31.050 333.600 ;
        RECT 28.950 317.400 31.050 319.500 ;
        RECT 13.950 311.400 18.450 312.450 ;
        RECT 13.950 310.950 16.050 311.400 ;
        RECT 13.950 308.850 16.050 309.750 ;
        RECT 7.950 298.500 10.050 300.600 ;
        RECT 17.400 265.050 18.450 311.400 ;
        RECT 19.950 311.400 24.450 312.450 ;
        RECT 19.950 310.950 22.050 311.400 ;
        RECT 19.950 308.850 22.050 309.750 ;
        RECT 16.950 262.950 19.050 265.050 ;
        RECT 23.400 199.050 24.450 311.400 ;
        RECT 29.250 305.400 30.450 317.400 ;
        RECT 31.950 314.250 34.050 315.150 ;
        RECT 31.950 310.950 34.050 313.050 ;
        RECT 28.950 303.300 31.050 305.400 ;
        RECT 29.250 299.700 30.450 303.300 ;
        RECT 32.400 301.050 33.450 310.950 ;
        RECT 41.400 310.050 42.450 379.950 ;
        RECT 47.400 340.050 48.450 382.950 ;
        RECT 46.950 337.950 49.050 340.050 ;
        RECT 40.950 307.950 43.050 310.050 ;
        RECT 52.950 307.950 55.050 310.050 ;
        RECT 28.950 297.600 31.050 299.700 ;
        RECT 31.950 298.950 34.050 301.050 ;
        RECT 32.400 276.450 33.450 298.950 ;
        RECT 29.400 275.400 33.450 276.450 ;
        RECT 29.400 270.450 30.450 275.400 ;
        RECT 31.950 272.250 34.050 273.150 ;
        RECT 31.950 270.450 34.050 271.050 ;
        RECT 29.400 269.400 34.050 270.450 ;
        RECT 31.950 268.950 34.050 269.400 ;
        RECT 35.250 269.250 36.750 270.150 ;
        RECT 37.950 268.950 40.050 271.050 ;
        RECT 41.250 269.250 43.050 270.150 ;
        RECT 49.950 268.950 52.050 271.050 ;
        RECT 34.950 265.950 37.050 268.050 ;
        RECT 38.250 266.850 39.750 267.750 ;
        RECT 40.950 265.950 43.050 268.050 ;
        RECT 46.950 265.950 49.050 268.050 ;
        RECT 35.400 238.050 36.450 265.950 ;
        RECT 37.950 262.950 40.050 265.050 ;
        RECT 38.400 241.050 39.450 262.950 ;
        RECT 37.950 238.950 40.050 241.050 ;
        RECT 41.250 239.250 42.750 240.150 ;
        RECT 43.950 238.950 46.050 241.050 ;
        RECT 34.950 235.950 37.050 238.050 ;
        RECT 38.250 236.850 39.750 237.750 ;
        RECT 40.950 235.950 43.050 238.050 ;
        RECT 44.250 236.850 46.050 237.750 ;
        RECT 34.950 233.850 37.050 234.750 ;
        RECT 22.950 196.950 25.050 199.050 ;
        RECT 34.950 196.950 37.050 199.050 ;
        RECT 34.950 194.850 37.050 195.750 ;
        RECT 34.950 190.950 37.050 193.050 ;
        RECT 35.400 169.050 36.450 190.950 ;
        RECT 31.950 167.250 33.750 168.150 ;
        RECT 34.950 166.950 37.050 169.050 ;
        RECT 31.950 163.950 34.050 166.050 ;
        RECT 35.250 164.850 37.050 165.750 ;
        RECT 32.400 162.450 33.450 163.950 ;
        RECT 32.400 161.400 36.450 162.450 ;
        RECT 7.950 135.300 10.050 137.400 ;
        RECT 8.550 131.700 9.750 135.300 ;
        RECT 28.950 134.400 31.050 136.500 ;
        RECT 4.950 127.950 7.050 130.050 ;
        RECT 7.950 129.600 10.050 131.700 ;
        RECT 5.400 124.050 6.450 127.950 ;
        RECT 4.950 121.950 7.050 124.050 ;
        RECT 4.950 119.850 7.050 120.750 ;
        RECT 8.550 117.600 9.750 129.600 ;
        RECT 10.950 127.950 13.050 130.050 ;
        RECT 7.950 115.500 10.050 117.600 ;
        RECT 7.950 62.400 10.050 64.500 ;
        RECT 8.400 45.600 9.600 62.400 ;
        RECT 11.400 51.450 12.450 127.950 ;
        RECT 16.950 125.250 19.050 126.150 ;
        RECT 19.950 124.950 22.050 127.050 ;
        RECT 22.950 125.250 25.050 126.150 ;
        RECT 16.950 123.450 19.050 124.050 ;
        RECT 20.400 123.450 21.450 124.950 ;
        RECT 16.950 122.400 21.450 123.450 ;
        RECT 16.950 121.950 19.050 122.400 ;
        RECT 22.950 121.950 25.050 124.050 ;
        RECT 13.950 53.250 16.050 54.150 ;
        RECT 13.950 51.450 16.050 52.050 ;
        RECT 11.400 50.400 16.050 51.450 ;
        RECT 17.400 51.450 18.450 121.950 ;
        RECT 29.400 117.600 30.600 134.400 ;
        RECT 35.400 130.050 36.450 161.400 ;
        RECT 34.950 127.950 37.050 130.050 ;
        RECT 28.950 115.500 31.050 117.600 ;
        RECT 35.400 97.050 36.450 127.950 ;
        RECT 47.400 124.050 48.450 265.950 ;
        RECT 50.400 193.050 51.450 268.950 ;
        RECT 53.400 238.050 54.450 307.950 ;
        RECT 52.950 235.950 55.050 238.050 ;
        RECT 62.400 202.050 63.450 484.950 ;
        RECT 64.950 481.950 67.050 484.050 ;
        RECT 68.250 482.850 69.750 483.750 ;
        RECT 70.950 481.950 73.050 484.050 ;
        RECT 71.400 481.050 72.450 481.950 ;
        RECT 95.400 481.050 96.450 527.400 ;
        RECT 97.950 526.950 100.050 529.050 ;
        RECT 97.950 524.850 100.050 525.750 ;
        RECT 107.250 521.400 108.450 533.400 ;
        RECT 109.950 530.250 112.050 531.150 ;
        RECT 109.950 526.950 112.050 529.050 ;
        RECT 106.950 519.300 109.050 521.400 ;
        RECT 107.250 515.700 108.450 519.300 ;
        RECT 106.950 513.600 109.050 515.700 ;
        RECT 110.400 496.050 111.450 526.950 ;
        RECT 109.950 493.950 112.050 496.050 ;
        RECT 113.400 490.050 114.450 556.950 ;
        RECT 118.950 553.950 121.050 556.050 ;
        RECT 122.250 554.850 123.750 555.750 ;
        RECT 124.950 553.950 127.050 556.050 ;
        RECT 109.950 487.950 112.050 490.050 ;
        RECT 112.950 487.950 115.050 490.050 ;
        RECT 115.950 488.250 118.050 489.150 ;
        RECT 110.400 487.050 111.450 487.950 ;
        RECT 106.950 485.250 108.750 486.150 ;
        RECT 109.950 484.950 112.050 487.050 ;
        RECT 113.250 485.250 114.750 486.150 ;
        RECT 115.950 484.950 118.050 487.050 ;
        RECT 106.950 481.950 109.050 484.050 ;
        RECT 110.250 482.850 111.750 483.750 ;
        RECT 112.950 481.950 115.050 484.050 ;
        RECT 70.950 478.950 73.050 481.050 ;
        RECT 94.950 478.950 97.050 481.050 ;
        RECT 94.950 455.250 97.050 456.150 ;
        RECT 97.950 455.850 100.050 456.750 ;
        RECT 94.950 451.950 97.050 454.050 ;
        RECT 64.950 423.300 67.050 425.400 ;
        RECT 65.250 419.700 66.450 423.300 ;
        RECT 79.950 422.400 82.050 424.500 ;
        RECT 64.950 417.600 67.050 419.700 ;
        RECT 65.250 405.600 66.450 417.600 ;
        RECT 67.950 412.950 70.050 415.050 ;
        RECT 68.400 412.050 69.450 412.950 ;
        RECT 67.950 409.950 70.050 412.050 ;
        RECT 67.950 407.850 70.050 408.750 ;
        RECT 80.400 405.600 81.600 422.400 ;
        RECT 85.950 413.250 88.050 414.150 ;
        RECT 91.950 413.250 94.050 414.150 ;
        RECT 85.950 409.950 88.050 412.050 ;
        RECT 91.950 409.950 94.050 412.050 ;
        RECT 92.400 409.050 93.450 409.950 ;
        RECT 91.950 406.950 94.050 409.050 ;
        RECT 64.950 403.500 67.050 405.600 ;
        RECT 79.950 403.500 82.050 405.600 ;
        RECT 67.950 400.950 70.050 403.050 ;
        RECT 64.950 340.950 67.050 343.050 ;
        RECT 68.400 342.450 69.450 400.950 ;
        RECT 79.950 397.950 82.050 400.050 ;
        RECT 80.400 385.050 81.450 397.950 ;
        RECT 95.400 388.050 96.450 451.950 ;
        RECT 100.950 423.300 103.050 425.400 ;
        RECT 101.250 419.700 102.450 423.300 ;
        RECT 100.950 417.600 103.050 419.700 ;
        RECT 101.250 405.600 102.450 417.600 ;
        RECT 103.950 415.950 106.050 418.050 ;
        RECT 104.400 412.050 105.450 415.950 ;
        RECT 103.950 409.950 106.050 412.050 ;
        RECT 103.950 407.850 106.050 408.750 ;
        RECT 100.950 403.500 103.050 405.600 ;
        RECT 94.950 385.950 97.050 388.050 ;
        RECT 73.950 382.950 76.050 385.050 ;
        RECT 77.250 383.250 78.750 384.150 ;
        RECT 79.950 382.950 82.050 385.050 ;
        RECT 107.400 382.050 108.450 481.950 ;
        RECT 113.400 481.050 114.450 481.950 ;
        RECT 112.950 478.950 115.050 481.050 ;
        RECT 119.400 454.050 120.450 553.950 ;
        RECT 125.400 553.050 126.450 553.950 ;
        RECT 185.400 553.050 186.450 598.950 ;
        RECT 187.950 596.850 190.050 597.750 ;
        RECT 191.400 594.450 192.450 601.950 ;
        RECT 196.950 598.950 199.050 601.050 ;
        RECT 193.950 596.250 196.050 597.150 ;
        RECT 196.950 596.850 199.050 597.750 ;
        RECT 193.950 594.450 196.050 595.050 ;
        RECT 191.400 593.400 196.050 594.450 ;
        RECT 193.950 592.950 196.050 593.400 ;
        RECT 202.950 557.250 205.050 558.150 ;
        RECT 208.950 557.250 211.050 558.150 ;
        RECT 193.950 553.950 196.050 556.050 ;
        RECT 202.950 553.950 205.050 556.050 ;
        RECT 206.250 554.250 207.750 555.150 ;
        RECT 208.950 553.950 211.050 556.050 ;
        RECT 124.950 550.950 127.050 553.050 ;
        RECT 184.950 550.950 187.050 553.050 ;
        RECT 157.950 532.950 160.050 535.050 ;
        RECT 166.950 533.400 169.050 535.500 ;
        RECT 187.950 533.400 190.050 535.500 ;
        RECT 158.400 529.050 159.450 532.950 ;
        RECT 151.950 526.950 154.050 529.050 ;
        RECT 155.250 527.250 156.750 528.150 ;
        RECT 157.950 526.950 160.050 529.050 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 148.950 523.950 151.050 526.050 ;
        RECT 152.250 524.850 153.750 525.750 ;
        RECT 154.950 523.950 157.050 526.050 ;
        RECT 158.250 524.850 160.050 525.750 ;
        RECT 134.400 454.050 135.450 523.950 ;
        RECT 148.950 521.850 151.050 522.750 ;
        RECT 155.400 510.450 156.450 523.950 ;
        RECT 167.400 516.600 168.600 533.400 ;
        RECT 175.950 529.950 178.050 532.050 ;
        RECT 178.950 529.950 181.050 532.050 ;
        RECT 172.950 526.950 175.050 529.050 ;
        RECT 172.950 524.850 175.050 525.750 ;
        RECT 166.950 514.500 169.050 516.600 ;
        RECT 152.400 509.400 156.450 510.450 ;
        RECT 118.950 451.950 121.050 454.050 ;
        RECT 130.950 452.250 132.750 453.150 ;
        RECT 133.950 451.950 136.050 454.050 ;
        RECT 137.250 452.250 139.050 453.150 ;
        RECT 139.950 451.950 142.050 454.050 ;
        RECT 130.950 448.950 133.050 451.050 ;
        RECT 134.250 449.850 135.750 450.750 ;
        RECT 131.400 448.050 132.450 448.950 ;
        RECT 130.950 445.950 133.050 448.050 ;
        RECT 127.950 412.950 130.050 415.050 ;
        RECT 140.400 414.450 141.450 451.950 ;
        RECT 152.400 448.050 153.450 509.400 ;
        RECT 160.950 493.950 163.050 496.050 ;
        RECT 169.950 494.400 172.050 496.500 ;
        RECT 161.400 490.050 162.450 493.950 ;
        RECT 166.950 490.950 169.050 493.050 ;
        RECT 154.950 487.950 157.050 490.050 ;
        RECT 158.250 488.250 159.750 489.150 ;
        RECT 160.950 487.950 163.050 490.050 ;
        RECT 163.950 487.950 166.050 490.050 ;
        RECT 154.950 485.850 156.750 486.750 ;
        RECT 157.950 484.950 160.050 487.050 ;
        RECT 161.250 485.850 163.050 486.750 ;
        RECT 151.950 445.950 154.050 448.050 ;
        RECT 142.950 416.250 145.050 417.150 ;
        RECT 142.950 414.450 145.050 415.050 ;
        RECT 140.400 413.400 145.050 414.450 ;
        RECT 142.950 412.950 145.050 413.400 ;
        RECT 146.250 413.250 147.750 414.150 ;
        RECT 148.950 412.950 151.050 415.050 ;
        RECT 152.250 413.250 154.050 414.150 ;
        RECT 154.950 412.950 157.050 415.050 ;
        RECT 128.400 406.050 129.450 412.950 ;
        RECT 145.950 409.950 148.050 412.050 ;
        RECT 149.250 410.850 150.750 411.750 ;
        RECT 151.950 409.950 154.050 412.050 ;
        RECT 155.400 408.450 156.450 412.950 ;
        RECT 164.400 409.050 165.450 487.950 ;
        RECT 167.400 450.450 168.450 490.950 ;
        RECT 170.400 477.600 171.600 494.400 ;
        RECT 176.400 489.450 177.450 529.950 ;
        RECT 179.400 529.050 180.450 529.950 ;
        RECT 178.950 526.950 181.050 529.050 ;
        RECT 178.950 524.850 181.050 525.750 ;
        RECT 188.250 521.400 189.450 533.400 ;
        RECT 190.950 530.250 193.050 531.150 ;
        RECT 190.950 526.950 193.050 529.050 ;
        RECT 187.950 519.300 190.050 521.400 ;
        RECT 188.250 515.700 189.450 519.300 ;
        RECT 187.950 513.600 190.050 515.700 ;
        RECT 190.950 495.300 193.050 497.400 ;
        RECT 191.250 491.700 192.450 495.300 ;
        RECT 190.950 489.600 193.050 491.700 ;
        RECT 176.400 488.400 180.450 489.450 ;
        RECT 175.950 485.250 178.050 486.150 ;
        RECT 175.950 481.950 178.050 484.050 ;
        RECT 179.400 483.450 180.450 488.400 ;
        RECT 181.950 485.250 184.050 486.150 ;
        RECT 181.950 483.450 184.050 484.050 ;
        RECT 179.400 482.400 184.050 483.450 ;
        RECT 181.950 481.950 184.050 482.400 ;
        RECT 176.400 481.050 177.450 481.950 ;
        RECT 175.950 478.950 178.050 481.050 ;
        RECT 191.250 477.600 192.450 489.600 ;
        RECT 194.400 484.050 195.450 553.950 ;
        RECT 203.400 550.050 204.450 553.950 ;
        RECT 205.950 550.950 208.050 553.050 ;
        RECT 202.950 547.950 205.050 550.050 ;
        RECT 203.400 529.050 204.450 547.950 ;
        RECT 202.950 526.950 205.050 529.050 ;
        RECT 193.950 481.950 196.050 484.050 ;
        RECT 193.950 479.850 196.050 480.750 ;
        RECT 169.950 475.500 172.050 477.600 ;
        RECT 190.950 475.500 193.050 477.600 ;
        RECT 217.950 460.950 220.050 463.050 ;
        RECT 218.400 460.050 219.450 460.950 ;
        RECT 217.950 457.950 220.050 460.050 ;
        RECT 214.950 455.250 217.050 456.150 ;
        RECT 217.950 455.850 220.050 456.750 ;
        RECT 169.950 452.250 171.750 453.150 ;
        RECT 172.950 451.950 175.050 454.050 ;
        RECT 176.250 452.250 178.050 453.150 ;
        RECT 214.950 451.950 217.050 454.050 ;
        RECT 169.950 450.450 172.050 451.050 ;
        RECT 167.400 449.400 172.050 450.450 ;
        RECT 173.250 449.850 174.750 450.750 ;
        RECT 167.400 418.050 168.450 449.400 ;
        RECT 169.950 448.950 172.050 449.400 ;
        RECT 175.950 448.950 178.050 451.050 ;
        RECT 176.400 421.050 177.450 448.950 ;
        RECT 175.950 418.950 178.050 421.050 ;
        RECT 196.950 418.950 199.050 421.050 ;
        RECT 166.950 415.950 169.050 418.050 ;
        RECT 176.400 412.050 177.450 418.950 ;
        RECT 190.950 415.950 193.050 418.050 ;
        RECT 191.400 415.050 192.450 415.950 ;
        RECT 197.400 415.050 198.450 418.950 ;
        RECT 208.950 415.950 211.050 418.050 ;
        RECT 187.950 413.250 189.750 414.150 ;
        RECT 190.950 412.950 193.050 415.050 ;
        RECT 194.250 413.250 195.750 414.150 ;
        RECT 196.950 412.950 199.050 415.050 ;
        RECT 200.250 413.250 202.050 414.150 ;
        RECT 175.950 409.950 178.050 412.050 ;
        RECT 187.950 409.950 190.050 412.050 ;
        RECT 191.250 410.850 192.750 411.750 ;
        RECT 193.950 409.950 196.050 412.050 ;
        RECT 197.250 410.850 198.750 411.750 ;
        RECT 199.950 409.950 202.050 412.050 ;
        RECT 152.400 407.400 156.450 408.450 ;
        RECT 127.950 403.950 130.050 406.050 ;
        RECT 121.950 383.250 124.050 384.150 ;
        RECT 124.950 383.850 127.050 384.750 ;
        RECT 73.950 380.850 75.750 381.750 ;
        RECT 76.950 379.950 79.050 382.050 ;
        RECT 80.250 380.850 81.750 381.750 ;
        RECT 82.950 381.450 85.050 382.050 ;
        RECT 82.950 380.400 87.450 381.450 ;
        RECT 82.950 379.950 85.050 380.400 ;
        RECT 82.950 377.850 85.050 378.750 ;
        RECT 70.950 344.250 73.050 345.150 ;
        RECT 70.950 342.450 73.050 343.050 ;
        RECT 68.400 341.400 73.050 342.450 ;
        RECT 70.950 340.950 73.050 341.400 ;
        RECT 74.250 341.250 75.750 342.150 ;
        RECT 76.950 340.950 79.050 343.050 ;
        RECT 80.250 341.250 82.050 342.150 ;
        RECT 65.400 316.050 66.450 340.950 ;
        RECT 73.950 337.950 76.050 340.050 ;
        RECT 77.250 338.850 78.750 339.750 ;
        RECT 79.950 337.950 82.050 340.050 ;
        RECT 80.400 337.050 81.450 337.950 ;
        RECT 86.400 337.050 87.450 380.400 ;
        RECT 106.950 379.950 109.050 382.050 ;
        RECT 121.950 379.950 124.050 382.050 ;
        RECT 121.950 344.250 124.050 345.150 ;
        RECT 128.400 343.050 129.450 403.950 ;
        RECT 152.400 343.050 153.450 407.400 ;
        RECT 160.950 406.950 163.050 409.050 ;
        RECT 163.950 406.950 166.050 409.050 ;
        RECT 157.950 383.250 160.050 384.150 ;
        RECT 157.950 381.450 160.050 382.050 ;
        RECT 161.400 381.450 162.450 406.950 ;
        RECT 163.950 385.950 166.050 388.050 ;
        RECT 166.950 387.450 169.050 388.050 ;
        RECT 166.950 386.400 171.450 387.450 ;
        RECT 166.950 385.950 169.050 386.400 ;
        RECT 164.400 385.050 165.450 385.950 ;
        RECT 163.950 382.950 166.050 385.050 ;
        RECT 167.250 383.850 169.050 384.750 ;
        RECT 157.950 380.400 162.450 381.450 ;
        RECT 163.950 380.850 166.050 381.750 ;
        RECT 157.950 379.950 160.050 380.400 ;
        RECT 170.400 379.050 171.450 386.400 ;
        RECT 176.400 382.050 177.450 409.950 ;
        RECT 188.400 409.050 189.450 409.950 ;
        RECT 178.950 406.950 181.050 409.050 ;
        RECT 187.950 406.950 190.050 409.050 ;
        RECT 175.950 379.950 178.050 382.050 ;
        RECT 169.950 376.950 172.050 379.050 ;
        RECT 157.950 345.450 160.050 346.050 ;
        RECT 155.400 344.400 160.050 345.450 ;
        RECT 112.950 341.250 114.750 342.150 ;
        RECT 115.950 340.950 118.050 343.050 ;
        RECT 119.250 341.250 120.750 342.150 ;
        RECT 121.950 340.950 124.050 343.050 ;
        RECT 127.950 340.950 130.050 343.050 ;
        RECT 151.950 340.950 154.050 343.050 ;
        RECT 112.950 337.950 115.050 340.050 ;
        RECT 116.250 338.850 117.750 339.750 ;
        RECT 118.950 337.950 121.050 340.050 ;
        RECT 155.400 339.450 156.450 344.400 ;
        RECT 157.950 343.950 160.050 344.400 ;
        RECT 161.250 344.250 162.750 345.150 ;
        RECT 163.950 343.950 166.050 346.050 ;
        RECT 157.950 341.850 159.750 342.750 ;
        RECT 160.950 340.950 163.050 343.050 ;
        RECT 164.250 341.850 166.050 342.750 ;
        RECT 155.400 338.400 159.450 339.450 ;
        RECT 70.950 334.950 73.050 337.050 ;
        RECT 79.950 334.950 82.050 337.050 ;
        RECT 85.950 334.950 88.050 337.050 ;
        RECT 64.950 313.950 67.050 316.050 ;
        RECT 64.950 311.850 66.750 312.750 ;
        RECT 67.950 312.450 70.050 313.050 ;
        RECT 71.400 312.450 72.450 334.950 ;
        RECT 113.400 322.050 114.450 337.950 ;
        RECT 119.400 337.050 120.450 337.950 ;
        RECT 118.950 334.950 121.050 337.050 ;
        RECT 112.950 319.950 115.050 322.050 ;
        RECT 76.950 313.950 79.050 316.050 ;
        RECT 136.950 313.950 139.050 316.050 ;
        RECT 67.950 311.400 72.450 312.450 ;
        RECT 67.950 310.950 70.050 311.400 ;
        RECT 67.950 308.850 70.050 309.750 ;
        RECT 71.400 268.050 72.450 311.400 ;
        RECT 73.950 311.250 76.050 312.150 ;
        RECT 73.950 307.950 76.050 310.050 ;
        RECT 77.400 271.050 78.450 313.950 ;
        RECT 112.950 310.950 115.050 313.050 ;
        RECT 118.950 312.450 121.050 313.050 ;
        RECT 118.950 311.400 123.450 312.450 ;
        RECT 118.950 310.950 121.050 311.400 ;
        RECT 112.950 308.850 115.050 309.750 ;
        RECT 118.950 308.850 121.050 309.750 ;
        RECT 94.950 278.400 97.050 280.500 ;
        RECT 115.950 279.300 118.050 281.400 ;
        RECT 82.950 272.250 85.050 273.150 ;
        RECT 73.950 269.250 75.750 270.150 ;
        RECT 76.950 268.950 79.050 271.050 ;
        RECT 80.250 269.250 81.750 270.150 ;
        RECT 82.950 268.950 85.050 271.050 ;
        RECT 83.400 268.050 84.450 268.950 ;
        RECT 70.950 265.950 73.050 268.050 ;
        RECT 73.950 265.950 76.050 268.050 ;
        RECT 77.250 266.850 78.750 267.750 ;
        RECT 79.950 265.950 82.050 268.050 ;
        RECT 82.950 265.950 85.050 268.050 ;
        RECT 67.950 238.950 70.050 241.050 ;
        RECT 61.950 199.950 64.050 202.050 ;
        RECT 55.950 194.850 58.050 195.750 ;
        RECT 49.950 190.950 52.050 193.050 ;
        RECT 68.400 172.050 69.450 238.950 ;
        RECT 80.400 238.050 81.450 265.950 ;
        RECT 82.950 259.950 85.050 262.050 ;
        RECT 95.400 261.600 96.600 278.400 ;
        RECT 116.250 275.700 117.450 279.300 ;
        RECT 115.950 273.600 118.050 275.700 ;
        RECT 100.950 269.250 103.050 270.150 ;
        RECT 106.950 269.250 109.050 270.150 ;
        RECT 100.950 265.950 103.050 268.050 ;
        RECT 106.950 265.950 109.050 268.050 ;
        RECT 101.400 262.050 102.450 265.950 ;
        RECT 83.400 241.050 84.450 259.950 ;
        RECT 94.950 259.500 97.050 261.600 ;
        RECT 100.950 259.950 103.050 262.050 ;
        RECT 82.950 238.950 85.050 241.050 ;
        RECT 86.250 239.250 87.750 240.150 ;
        RECT 88.950 238.950 91.050 241.050 ;
        RECT 103.950 238.950 106.050 241.050 ;
        RECT 79.950 235.950 82.050 238.050 ;
        RECT 83.250 236.850 84.750 237.750 ;
        RECT 85.950 235.950 88.050 238.050 ;
        RECT 89.250 236.850 91.050 237.750 ;
        RECT 79.950 233.850 82.050 234.750 ;
        RECT 85.950 199.950 88.050 202.050 ;
        RECT 94.950 199.950 97.050 202.050 ;
        RECT 98.250 200.250 99.750 201.150 ;
        RECT 100.950 199.950 103.050 202.050 ;
        RECT 76.950 172.950 79.050 175.050 ;
        RECT 67.950 169.950 70.050 172.050 ;
        RECT 68.400 169.050 69.450 169.950 ;
        RECT 67.950 166.950 70.050 169.050 ;
        RECT 71.250 167.250 72.750 168.150 ;
        RECT 73.950 166.950 76.050 169.050 ;
        RECT 77.400 166.050 78.450 172.950 ;
        RECT 86.400 166.050 87.450 199.950 ;
        RECT 94.950 197.850 96.750 198.750 ;
        RECT 97.950 196.950 100.050 199.050 ;
        RECT 101.250 197.850 103.050 198.750 ;
        RECT 88.950 173.400 91.050 175.500 ;
        RECT 98.400 175.050 99.450 196.950 ;
        RECT 100.950 193.950 103.050 196.050 ;
        RECT 67.950 164.850 69.750 165.750 ;
        RECT 70.950 163.950 73.050 166.050 ;
        RECT 74.250 164.850 75.750 165.750 ;
        RECT 76.950 163.950 79.050 166.050 ;
        RECT 85.950 163.950 88.050 166.050 ;
        RECT 71.400 144.450 72.450 163.950 ;
        RECT 76.950 161.850 79.050 162.750 ;
        RECT 89.400 156.600 90.600 173.400 ;
        RECT 97.950 172.950 100.050 175.050 ;
        RECT 101.400 169.050 102.450 193.950 ;
        RECT 94.950 166.950 97.050 169.050 ;
        RECT 100.950 166.950 103.050 169.050 ;
        RECT 94.950 164.850 97.050 165.750 ;
        RECT 100.950 164.850 103.050 165.750 ;
        RECT 104.400 162.450 105.450 238.950 ;
        RECT 107.400 196.050 108.450 265.950 ;
        RECT 116.250 261.600 117.450 273.600 ;
        RECT 118.950 265.950 121.050 268.050 ;
        RECT 118.950 263.850 121.050 264.750 ;
        RECT 115.950 259.500 118.050 261.600 ;
        RECT 122.400 247.050 123.450 311.400 ;
        RECT 133.950 310.950 136.050 313.050 ;
        RECT 127.950 271.950 130.050 274.050 ;
        RECT 121.950 244.950 124.050 247.050 ;
        RECT 128.400 238.050 129.450 271.950 ;
        RECT 134.400 241.050 135.450 310.950 ;
        RECT 133.950 238.950 136.050 241.050 ;
        RECT 124.950 236.250 126.750 237.150 ;
        RECT 127.950 235.950 130.050 238.050 ;
        RECT 131.250 236.250 133.050 237.150 ;
        RECT 124.950 232.950 127.050 235.050 ;
        RECT 128.250 233.850 129.750 234.750 ;
        RECT 130.950 234.450 133.050 235.050 ;
        RECT 134.400 234.450 135.450 238.950 ;
        RECT 130.950 233.400 135.450 234.450 ;
        RECT 130.950 232.950 133.050 233.400 ;
        RECT 109.950 206.400 112.050 208.500 ;
        RECT 106.950 193.950 109.050 196.050 ;
        RECT 110.400 189.600 111.600 206.400 ;
        RECT 125.400 202.050 126.450 232.950 ;
        RECT 130.950 207.300 133.050 209.400 ;
        RECT 131.250 203.700 132.450 207.300 ;
        RECT 124.950 199.950 127.050 202.050 ;
        RECT 127.950 199.950 130.050 202.050 ;
        RECT 130.950 201.600 133.050 203.700 ;
        RECT 115.950 197.250 118.050 198.150 ;
        RECT 118.950 196.950 121.050 199.050 ;
        RECT 121.950 197.250 124.050 198.150 ;
        RECT 115.950 195.450 118.050 196.050 ;
        RECT 119.400 195.450 120.450 196.950 ;
        RECT 115.950 194.400 120.450 195.450 ;
        RECT 115.950 193.950 118.050 194.400 ;
        RECT 121.950 193.950 124.050 196.050 ;
        RECT 109.950 187.500 112.050 189.600 ;
        RECT 109.950 173.400 112.050 175.500 ;
        RECT 104.400 161.400 108.450 162.450 ;
        RECT 110.250 161.400 111.450 173.400 ;
        RECT 112.950 170.250 115.050 171.150 ;
        RECT 125.400 169.050 126.450 199.950 ;
        RECT 112.950 166.950 115.050 169.050 ;
        RECT 124.950 166.950 127.050 169.050 ;
        RECT 88.950 154.500 91.050 156.600 ;
        RECT 71.400 143.400 75.450 144.450 ;
        RECT 70.950 124.950 73.050 127.050 ;
        RECT 40.950 121.950 43.050 124.050 ;
        RECT 46.950 121.950 49.050 124.050 ;
        RECT 70.950 122.850 73.050 123.750 ;
        RECT 37.950 97.950 40.050 100.050 ;
        RECT 41.400 97.050 42.450 121.950 ;
        RECT 67.950 97.950 70.050 100.050 ;
        RECT 34.950 94.950 37.050 97.050 ;
        RECT 38.250 95.850 39.750 96.750 ;
        RECT 40.950 94.950 43.050 97.050 ;
        RECT 34.950 92.850 37.050 93.750 ;
        RECT 40.950 92.850 43.050 93.750 ;
        RECT 28.950 63.300 31.050 65.400 ;
        RECT 29.250 59.700 30.450 63.300 ;
        RECT 28.950 57.600 31.050 59.700 ;
        RECT 19.950 53.250 22.050 54.150 ;
        RECT 19.950 51.450 22.050 52.050 ;
        RECT 17.400 50.400 22.050 51.450 ;
        RECT 13.950 49.950 16.050 50.400 ;
        RECT 19.950 49.950 22.050 50.400 ;
        RECT 7.950 43.500 10.050 45.600 ;
        RECT 20.400 25.050 21.450 49.950 ;
        RECT 29.250 45.600 30.450 57.600 ;
        RECT 68.400 55.050 69.450 97.950 ;
        RECT 74.400 91.050 75.450 143.400 ;
        RECT 103.950 134.400 106.050 136.500 ;
        RECT 85.950 121.950 88.050 124.050 ;
        RECT 91.950 122.850 94.050 123.750 ;
        RECT 76.950 92.250 78.750 93.150 ;
        RECT 79.950 91.950 82.050 94.050 ;
        RECT 83.250 92.250 85.050 93.150 ;
        RECT 70.950 88.950 73.050 91.050 ;
        RECT 73.950 88.950 76.050 91.050 ;
        RECT 76.950 88.950 79.050 91.050 ;
        RECT 80.250 89.850 81.750 90.750 ;
        RECT 82.950 90.450 85.050 91.050 ;
        RECT 86.400 90.450 87.450 121.950 ;
        RECT 104.400 117.600 105.600 134.400 ;
        RECT 103.950 115.500 106.050 117.600 ;
        RECT 107.400 112.050 108.450 161.400 ;
        RECT 109.950 159.300 112.050 161.400 ;
        RECT 110.250 155.700 111.450 159.300 ;
        RECT 109.950 153.600 112.050 155.700 ;
        RECT 124.950 135.300 127.050 137.400 ;
        RECT 125.250 131.700 126.450 135.300 ;
        RECT 124.950 129.600 127.050 131.700 ;
        RECT 109.950 125.250 112.050 126.150 ;
        RECT 112.950 124.950 115.050 127.050 ;
        RECT 115.950 125.250 118.050 126.150 ;
        RECT 109.950 121.950 112.050 124.050 ;
        RECT 113.400 123.450 114.450 124.950 ;
        RECT 115.950 123.450 118.050 124.050 ;
        RECT 113.400 122.400 118.050 123.450 ;
        RECT 115.950 121.950 118.050 122.400 ;
        RECT 110.400 121.050 111.450 121.950 ;
        RECT 109.950 118.950 112.050 121.050 ;
        RECT 121.950 118.950 124.050 121.050 ;
        RECT 106.950 109.950 109.050 112.050 ;
        RECT 115.950 109.950 118.050 112.050 ;
        RECT 116.400 97.050 117.450 109.950 ;
        RECT 122.400 97.050 123.450 118.950 ;
        RECT 125.250 117.600 126.450 129.600 ;
        RECT 128.400 124.050 129.450 199.950 ;
        RECT 131.250 189.600 132.450 201.600 ;
        RECT 133.950 195.450 136.050 196.050 ;
        RECT 137.400 195.450 138.450 313.950 ;
        RECT 158.400 310.050 159.450 338.400 ;
        RECT 154.950 308.250 156.750 309.150 ;
        RECT 157.950 307.950 160.050 310.050 ;
        RECT 161.250 308.250 163.050 309.150 ;
        RECT 154.950 304.950 157.050 307.050 ;
        RECT 158.250 305.850 159.750 306.750 ;
        RECT 160.950 304.950 163.050 307.050 ;
        RECT 155.400 298.050 156.450 304.950 ;
        RECT 154.950 295.950 157.050 298.050 ;
        RECT 157.950 268.950 160.050 271.050 ;
        RECT 154.950 266.250 157.050 267.150 ;
        RECT 157.950 266.850 160.050 267.750 ;
        RECT 154.950 262.950 157.050 265.050 ;
        RECT 155.400 250.050 156.450 262.950 ;
        RECT 154.950 247.950 157.050 250.050 ;
        RECT 155.400 202.050 156.450 247.950 ;
        RECT 161.400 244.050 162.450 304.950 ;
        RECT 160.950 241.950 163.050 244.050 ;
        RECT 166.950 243.450 169.050 244.050 ;
        RECT 166.950 242.400 171.450 243.450 ;
        RECT 166.950 241.950 169.050 242.400 ;
        RECT 161.400 237.450 162.450 241.950 ;
        RECT 163.950 239.250 166.050 240.150 ;
        RECT 166.950 239.850 169.050 240.750 ;
        RECT 163.950 237.450 166.050 238.050 ;
        RECT 161.400 236.400 166.050 237.450 ;
        RECT 163.950 235.950 166.050 236.400 ;
        RECT 170.400 235.050 171.450 242.400 ;
        RECT 169.950 232.950 172.050 235.050 ;
        RECT 179.400 202.050 180.450 406.950 ;
        RECT 196.950 385.950 199.050 388.050 ;
        RECT 202.950 385.950 205.050 388.050 ;
        RECT 197.400 375.450 198.450 385.950 ;
        RECT 209.400 385.050 210.450 415.950 ;
        RECT 215.400 412.050 216.450 451.950 ;
        RECT 214.950 409.950 217.050 412.050 ;
        RECT 199.950 383.250 202.050 384.150 ;
        RECT 202.950 383.850 205.050 384.750 ;
        RECT 205.950 383.250 207.750 384.150 ;
        RECT 208.950 382.950 211.050 385.050 ;
        RECT 199.950 381.450 202.050 382.050 ;
        RECT 199.950 380.400 204.450 381.450 ;
        RECT 199.950 379.950 202.050 380.400 ;
        RECT 200.400 379.050 201.450 379.950 ;
        RECT 199.950 376.950 202.050 379.050 ;
        RECT 197.400 374.400 201.450 375.450 ;
        RECT 200.400 343.050 201.450 374.400 ;
        RECT 199.950 340.950 202.050 343.050 ;
        RECT 203.400 340.050 204.450 380.400 ;
        RECT 205.950 379.950 208.050 382.050 ;
        RECT 209.250 380.850 211.050 381.750 ;
        RECT 196.950 338.250 199.050 339.150 ;
        RECT 199.950 338.850 202.050 339.750 ;
        RECT 202.950 337.950 205.050 340.050 ;
        RECT 196.950 334.950 199.050 337.050 ;
        RECT 197.400 316.050 198.450 334.950 ;
        RECT 193.950 313.950 196.050 316.050 ;
        RECT 196.950 313.950 199.050 316.050 ;
        RECT 193.950 311.850 196.050 312.750 ;
        RECT 196.950 311.250 199.050 312.150 ;
        RECT 196.950 307.950 199.050 310.050 ;
        RECT 197.400 307.050 198.450 307.950 ;
        RECT 196.950 304.950 199.050 307.050 ;
        RECT 202.950 295.950 205.050 298.050 ;
        RECT 193.950 275.250 196.050 276.150 ;
        RECT 190.950 272.250 192.750 273.150 ;
        RECT 193.950 271.950 196.050 274.050 ;
        RECT 197.250 272.250 198.750 273.150 ;
        RECT 199.950 271.950 202.050 274.050 ;
        RECT 203.400 271.050 204.450 295.950 ;
        RECT 211.950 274.950 214.050 277.050 ;
        RECT 190.950 268.950 193.050 271.050 ;
        RECT 196.950 268.950 199.050 271.050 ;
        RECT 200.250 269.850 202.050 270.750 ;
        RECT 202.950 268.950 205.050 271.050 ;
        RECT 199.950 262.950 202.050 265.050 ;
        RECT 200.400 234.450 201.450 262.950 ;
        RECT 208.950 247.950 211.050 250.050 ;
        RECT 202.950 236.250 204.750 237.150 ;
        RECT 205.950 235.950 208.050 238.050 ;
        RECT 209.400 235.050 210.450 247.950 ;
        RECT 212.400 241.050 213.450 274.950 ;
        RECT 221.400 247.050 222.450 670.950 ;
        RECT 233.400 601.050 234.450 679.950 ;
        RECT 236.400 640.050 237.450 739.950 ;
        RECT 278.400 739.050 279.450 739.950 ;
        RECT 277.950 736.950 280.050 739.050 ;
        RECT 259.950 733.950 262.050 736.050 ;
        RECT 247.950 702.450 250.050 703.050 ;
        RECT 247.950 701.400 252.450 702.450 ;
        RECT 247.950 700.950 250.050 701.400 ;
        RECT 244.950 698.250 247.050 699.150 ;
        RECT 247.950 698.850 250.050 699.750 ;
        RECT 251.400 697.050 252.450 701.400 ;
        RECT 244.950 694.950 247.050 697.050 ;
        RECT 250.950 694.950 253.050 697.050 ;
        RECT 241.950 679.950 244.050 682.050 ;
        RECT 238.950 673.950 241.050 676.050 ;
        RECT 239.400 670.050 240.450 673.950 ;
        RECT 242.400 672.450 243.450 679.950 ;
        RECT 245.400 676.050 246.450 694.950 ;
        RECT 260.400 694.050 261.450 733.950 ;
        RECT 284.400 733.050 285.450 745.950 ;
        RECT 292.950 742.950 295.050 745.050 ;
        RECT 391.950 742.950 394.050 745.050 ;
        RECT 397.950 742.950 400.050 745.050 ;
        RECT 401.250 743.250 402.750 744.150 ;
        RECT 403.950 742.950 406.050 745.050 ;
        RECT 283.950 730.950 286.050 733.050 ;
        RECT 284.400 702.450 285.450 730.950 ;
        RECT 286.950 704.250 289.050 705.150 ;
        RECT 293.400 703.050 294.450 742.950 ;
        RECT 313.950 740.250 315.750 741.150 ;
        RECT 316.950 739.950 319.050 742.050 ;
        RECT 320.250 740.250 322.050 741.150 ;
        RECT 352.950 739.950 355.050 742.050 ;
        RECT 355.950 740.250 357.750 741.150 ;
        RECT 358.950 739.950 361.050 742.050 ;
        RECT 362.250 740.250 364.050 741.150 ;
        RECT 313.950 736.950 316.050 739.050 ;
        RECT 317.250 737.850 318.750 738.750 ;
        RECT 319.950 736.950 322.050 739.050 ;
        RECT 353.400 738.450 354.450 739.950 ;
        RECT 355.950 738.450 358.050 739.050 ;
        RECT 353.400 737.400 358.050 738.450 ;
        RECT 359.250 737.850 360.750 738.750 ;
        RECT 355.950 736.950 358.050 737.400 ;
        RECT 361.950 736.950 364.050 739.050 ;
        RECT 314.400 703.050 315.450 736.950 ;
        RECT 320.400 733.050 321.450 736.950 ;
        RECT 319.950 730.950 322.050 733.050 ;
        RECT 392.400 706.050 393.450 742.950 ;
        RECT 397.950 740.850 399.750 741.750 ;
        RECT 400.950 739.950 403.050 742.050 ;
        RECT 404.250 740.850 405.750 741.750 ;
        RECT 406.950 739.950 409.050 742.050 ;
        RECT 439.950 740.250 441.750 741.150 ;
        RECT 442.950 739.950 445.050 742.050 ;
        RECT 446.250 740.250 448.050 741.150 ;
        RECT 406.950 737.850 409.050 738.750 ;
        RECT 439.950 736.950 442.050 739.050 ;
        RECT 443.250 737.850 444.750 738.750 ;
        RECT 445.950 736.950 448.050 739.050 ;
        RECT 439.950 710.400 442.050 712.500 ;
        RECT 376.950 703.950 379.050 706.050 ;
        RECT 391.950 703.950 394.050 706.050 ;
        RECT 427.950 703.950 430.050 706.050 ;
        RECT 377.400 703.050 378.450 703.950 ;
        RECT 286.950 702.450 289.050 703.050 ;
        RECT 284.400 701.400 289.050 702.450 ;
        RECT 259.950 691.950 262.050 694.050 ;
        RECT 253.950 676.950 256.050 679.050 ;
        RECT 244.950 673.950 247.050 676.050 ;
        RECT 244.950 672.450 247.050 673.050 ;
        RECT 242.400 671.400 247.050 672.450 ;
        RECT 244.950 670.950 247.050 671.400 ;
        RECT 248.250 671.250 249.750 672.150 ;
        RECT 250.950 670.950 253.050 673.050 ;
        RECT 254.400 670.050 255.450 676.950 ;
        RECT 238.950 667.950 241.050 670.050 ;
        RECT 244.950 668.850 246.750 669.750 ;
        RECT 247.950 667.950 250.050 670.050 ;
        RECT 251.250 668.850 252.750 669.750 ;
        RECT 253.950 667.950 256.050 670.050 ;
        RECT 235.950 637.950 238.050 640.050 ;
        RECT 235.950 601.950 238.050 604.050 ;
        RECT 239.400 601.050 240.450 667.950 ;
        RECT 253.950 665.850 256.050 666.750 ;
        RECT 241.950 632.250 244.050 633.150 ;
        RECT 241.950 628.950 244.050 631.050 ;
        RECT 245.250 629.250 246.750 630.150 ;
        RECT 247.950 628.950 250.050 631.050 ;
        RECT 251.250 629.250 253.050 630.150 ;
        RECT 242.400 622.050 243.450 628.950 ;
        RECT 244.950 625.950 247.050 628.050 ;
        RECT 248.250 626.850 249.750 627.750 ;
        RECT 250.950 625.950 253.050 628.050 ;
        RECT 241.950 619.950 244.050 622.050 ;
        RECT 232.950 600.450 235.050 601.050 ;
        RECT 230.400 599.400 235.050 600.450 ;
        RECT 236.250 599.850 237.750 600.750 ;
        RECT 238.950 600.450 241.050 601.050 ;
        RECT 230.400 568.050 231.450 599.400 ;
        RECT 232.950 598.950 235.050 599.400 ;
        RECT 238.950 599.400 243.450 600.450 ;
        RECT 238.950 598.950 241.050 599.400 ;
        RECT 232.950 596.850 235.050 597.750 ;
        RECT 238.950 596.850 241.050 597.750 ;
        RECT 229.950 565.950 232.050 568.050 ;
        RECT 232.950 553.950 235.050 556.050 ;
        RECT 233.400 532.050 234.450 553.950 ;
        RECT 232.950 529.950 235.050 532.050 ;
        RECT 229.950 527.250 232.050 528.150 ;
        RECT 232.950 527.850 235.050 528.750 ;
        RECT 229.950 523.950 232.050 526.050 ;
        RECT 230.400 520.050 231.450 523.950 ;
        RECT 229.950 517.950 232.050 520.050 ;
        RECT 230.400 490.050 231.450 517.950 ;
        RECT 242.400 496.050 243.450 599.400 ;
        RECT 251.400 589.050 252.450 625.950 ;
        RECT 250.950 586.950 253.050 589.050 ;
        RECT 247.950 558.450 250.050 559.050 ;
        RECT 247.950 557.400 252.450 558.450 ;
        RECT 247.950 556.950 250.050 557.400 ;
        RECT 244.950 554.250 247.050 555.150 ;
        RECT 247.950 554.850 250.050 555.750 ;
        RECT 251.400 553.050 252.450 557.400 ;
        RECT 260.400 556.050 261.450 691.950 ;
        RECT 284.400 679.050 285.450 701.400 ;
        RECT 286.950 700.950 289.050 701.400 ;
        RECT 290.250 701.250 291.750 702.150 ;
        RECT 292.950 700.950 295.050 703.050 ;
        RECT 296.250 701.250 298.050 702.150 ;
        RECT 313.950 700.950 316.050 703.050 ;
        RECT 328.950 701.250 331.050 702.150 ;
        RECT 334.950 700.950 337.050 703.050 ;
        RECT 370.950 702.450 373.050 703.050 ;
        RECT 368.400 701.400 373.050 702.450 ;
        RECT 368.400 700.050 369.450 701.400 ;
        RECT 370.950 700.950 373.050 701.400 ;
        RECT 376.950 700.950 379.050 703.050 ;
        RECT 380.250 701.250 382.050 702.150 ;
        RECT 289.950 697.950 292.050 700.050 ;
        RECT 293.250 698.850 294.750 699.750 ;
        RECT 295.950 697.950 298.050 700.050 ;
        RECT 322.950 697.950 325.050 700.050 ;
        RECT 325.950 698.250 327.750 699.150 ;
        RECT 328.950 697.950 331.050 700.050 ;
        RECT 334.950 698.850 337.050 699.750 ;
        RECT 367.950 697.950 370.050 700.050 ;
        RECT 370.950 698.850 373.050 699.750 ;
        RECT 373.950 698.250 376.050 699.150 ;
        RECT 376.950 698.850 378.750 699.750 ;
        RECT 379.950 697.950 382.050 700.050 ;
        RECT 296.400 694.050 297.450 697.950 ;
        RECT 323.400 696.450 324.450 697.950 ;
        RECT 329.400 697.050 330.450 697.950 ;
        RECT 325.950 696.450 328.050 697.050 ;
        RECT 323.400 695.400 328.050 696.450 ;
        RECT 325.950 694.950 328.050 695.400 ;
        RECT 328.950 694.950 331.050 697.050 ;
        RECT 373.950 694.950 376.050 697.050 ;
        RECT 295.950 691.950 298.050 694.050 ;
        RECT 283.950 676.950 286.050 679.050 ;
        RECT 382.950 676.950 385.050 679.050 ;
        RECT 284.400 628.050 285.450 676.950 ;
        RECT 289.950 673.950 292.050 676.050 ;
        RECT 290.400 673.050 291.450 673.950 ;
        RECT 289.950 670.950 292.050 673.050 ;
        RECT 295.950 672.450 298.050 673.050 ;
        RECT 293.400 671.400 298.050 672.450 ;
        RECT 293.400 670.050 294.450 671.400 ;
        RECT 295.950 670.950 298.050 671.400 ;
        RECT 310.950 670.950 313.050 673.050 ;
        RECT 334.950 670.950 337.050 673.050 ;
        RECT 376.950 670.950 379.050 673.050 ;
        RECT 289.950 668.850 292.050 669.750 ;
        RECT 292.950 667.950 295.050 670.050 ;
        RECT 295.950 668.850 298.050 669.750 ;
        RECT 286.950 634.950 289.050 637.050 ;
        RECT 287.400 634.050 288.450 634.950 ;
        RECT 293.400 634.050 294.450 667.950 ;
        RECT 311.400 637.050 312.450 670.950 ;
        RECT 331.950 667.950 334.050 670.050 ;
        RECT 335.400 669.450 336.450 670.950 ;
        RECT 377.400 670.050 378.450 670.950 ;
        RECT 383.400 670.050 384.450 676.950 ;
        RECT 337.950 669.450 340.050 670.050 ;
        RECT 335.400 668.400 340.050 669.450 ;
        RECT 337.950 667.950 340.050 668.400 ;
        RECT 341.250 668.250 343.050 669.150 ;
        RECT 376.950 667.950 379.050 670.050 ;
        RECT 382.950 667.950 385.050 670.050 ;
        RECT 386.250 668.250 388.050 669.150 ;
        RECT 328.950 664.950 331.050 667.050 ;
        RECT 331.950 665.850 333.750 666.750 ;
        RECT 334.950 664.950 337.050 667.050 ;
        RECT 338.250 665.850 339.750 666.750 ;
        RECT 340.950 664.950 343.050 667.050 ;
        RECT 376.950 665.850 378.750 666.750 ;
        RECT 379.950 664.950 382.050 667.050 ;
        RECT 383.250 665.850 384.750 666.750 ;
        RECT 385.950 664.950 388.050 667.050 ;
        RECT 295.950 634.950 298.050 637.050 ;
        RECT 310.950 634.950 313.050 637.050 ;
        RECT 286.950 631.950 289.050 634.050 ;
        RECT 290.250 632.250 291.750 633.150 ;
        RECT 292.950 631.950 295.050 634.050 ;
        RECT 286.950 629.850 288.750 630.750 ;
        RECT 289.950 628.950 292.050 631.050 ;
        RECT 293.250 629.850 295.050 630.750 ;
        RECT 290.400 628.050 291.450 628.950 ;
        RECT 283.950 625.950 286.050 628.050 ;
        RECT 289.950 625.950 292.050 628.050 ;
        RECT 274.950 601.950 277.050 604.050 ;
        RECT 275.400 598.050 276.450 601.950 ;
        RECT 280.950 598.950 283.050 601.050 ;
        RECT 281.400 598.050 282.450 598.950 ;
        RECT 274.950 595.950 277.050 598.050 ;
        RECT 277.950 595.950 280.050 598.050 ;
        RECT 280.950 595.950 283.050 598.050 ;
        RECT 284.250 596.250 286.050 597.150 ;
        RECT 278.400 595.050 279.450 595.950 ;
        RECT 296.400 595.050 297.450 634.950 ;
        RECT 329.400 634.050 330.450 664.950 ;
        RECT 334.950 662.850 337.050 663.750 ;
        RECT 346.950 661.950 349.050 664.050 ;
        RECT 379.950 662.850 382.050 663.750 ;
        RECT 316.950 631.950 319.050 634.050 ;
        RECT 322.950 631.950 325.050 634.050 ;
        RECT 328.950 633.450 331.050 634.050 ;
        RECT 326.250 632.250 327.750 633.150 ;
        RECT 328.950 632.400 333.450 633.450 ;
        RECT 328.950 631.950 331.050 632.400 ;
        RECT 317.400 622.050 318.450 631.950 ;
        RECT 322.950 629.850 324.750 630.750 ;
        RECT 325.950 628.950 328.050 631.050 ;
        RECT 329.250 629.850 331.050 630.750 ;
        RECT 316.950 619.950 319.050 622.050 ;
        RECT 313.950 601.950 316.050 604.050 ;
        RECT 274.950 593.850 276.750 594.750 ;
        RECT 277.950 592.950 280.050 595.050 ;
        RECT 281.250 593.850 282.750 594.750 ;
        RECT 283.950 592.950 286.050 595.050 ;
        RECT 295.950 592.950 298.050 595.050 ;
        RECT 307.950 592.950 310.050 595.050 ;
        RECT 277.950 590.850 280.050 591.750 ;
        RECT 280.950 589.950 283.050 592.050 ;
        RECT 271.950 586.950 274.050 589.050 ;
        RECT 259.950 553.950 262.050 556.050 ;
        RECT 244.950 550.950 247.050 553.050 ;
        RECT 250.950 550.950 253.050 553.050 ;
        RECT 245.400 550.050 246.450 550.950 ;
        RECT 244.950 547.950 247.050 550.050 ;
        RECT 251.400 535.050 252.450 550.950 ;
        RECT 250.950 532.950 253.050 535.050 ;
        RECT 272.400 526.050 273.450 586.950 ;
        RECT 281.400 559.050 282.450 589.950 ;
        RECT 292.950 560.250 295.050 561.150 ;
        RECT 280.950 556.950 283.050 559.050 ;
        RECT 283.950 557.250 285.750 558.150 ;
        RECT 286.950 556.950 289.050 559.050 ;
        RECT 290.250 557.250 291.750 558.150 ;
        RECT 292.950 556.950 295.050 559.050 ;
        RECT 268.950 524.250 270.750 525.150 ;
        RECT 271.950 523.950 274.050 526.050 ;
        RECT 275.250 524.250 277.050 525.150 ;
        RECT 268.950 520.950 271.050 523.050 ;
        RECT 272.250 521.850 273.750 522.750 ;
        RECT 274.950 520.950 277.050 523.050 ;
        RECT 241.950 493.950 244.050 496.050 ;
        RECT 269.400 490.050 270.450 520.950 ;
        RECT 275.400 519.450 276.450 520.950 ;
        RECT 272.400 518.400 276.450 519.450 ;
        RECT 229.950 487.950 232.050 490.050 ;
        RECT 235.950 488.250 238.050 489.150 ;
        RECT 262.950 487.950 265.050 490.050 ;
        RECT 268.950 487.950 271.050 490.050 ;
        RECT 226.950 485.250 228.750 486.150 ;
        RECT 229.950 484.950 232.050 487.050 ;
        RECT 233.250 485.250 234.750 486.150 ;
        RECT 235.950 484.950 238.050 487.050 ;
        RECT 259.950 484.950 262.050 487.050 ;
        RECT 236.400 484.050 237.450 484.950 ;
        RECT 226.950 481.950 229.050 484.050 ;
        RECT 230.250 482.850 231.750 483.750 ;
        RECT 232.950 481.950 235.050 484.050 ;
        RECT 235.950 481.950 238.050 484.050 ;
        RECT 253.950 481.950 256.050 484.050 ;
        RECT 233.400 481.050 234.450 481.950 ;
        RECT 232.950 478.950 235.050 481.050 ;
        RECT 254.400 454.050 255.450 481.950 ;
        RECT 250.950 452.250 252.750 453.150 ;
        RECT 253.950 451.950 256.050 454.050 ;
        RECT 257.250 452.250 259.050 453.150 ;
        RECT 254.250 449.850 255.750 450.750 ;
        RECT 256.950 450.450 259.050 451.050 ;
        RECT 260.400 450.450 261.450 484.950 ;
        RECT 256.950 449.400 261.450 450.450 ;
        RECT 256.950 448.950 259.050 449.400 ;
        RECT 257.400 448.050 258.450 448.950 ;
        RECT 256.950 445.950 259.050 448.050 ;
        RECT 229.950 413.250 232.050 414.150 ;
        RECT 235.950 413.250 238.050 414.150 ;
        RECT 229.950 409.950 232.050 412.050 ;
        RECT 233.250 410.250 234.750 411.150 ;
        RECT 235.950 409.950 238.050 412.050 ;
        RECT 230.400 403.050 231.450 409.950 ;
        RECT 232.950 406.950 235.050 409.050 ;
        RECT 236.400 406.050 237.450 409.950 ;
        RECT 235.950 403.950 238.050 406.050 ;
        RECT 229.950 400.950 232.050 403.050 ;
        RECT 244.950 400.950 247.050 403.050 ;
        RECT 245.400 388.050 246.450 400.950 ;
        RECT 244.950 385.950 247.050 388.050 ;
        RECT 244.950 383.850 247.050 384.750 ;
        RECT 247.950 383.250 250.050 384.150 ;
        RECT 250.950 382.950 253.050 385.050 ;
        RECT 247.950 379.950 250.050 382.050 ;
        RECT 223.950 343.950 226.050 346.050 ;
        RECT 235.950 343.950 238.050 346.050 ;
        RECT 238.950 344.250 241.050 345.150 ;
        RECT 220.950 244.950 223.050 247.050 ;
        RECT 211.950 238.950 214.050 241.050 ;
        RECT 212.400 238.050 213.450 238.950 ;
        RECT 211.950 235.950 214.050 238.050 ;
        RECT 202.950 234.450 205.050 235.050 ;
        RECT 200.400 233.400 205.050 234.450 ;
        RECT 206.250 233.850 207.750 234.750 ;
        RECT 202.950 232.950 205.050 233.400 ;
        RECT 208.950 232.950 211.050 235.050 ;
        RECT 212.250 233.850 214.050 234.750 ;
        RECT 208.950 230.850 211.050 231.750 ;
        RECT 217.950 203.250 220.050 204.150 ;
        RECT 224.400 202.050 225.450 343.950 ;
        RECT 226.950 313.950 229.050 316.050 ;
        RECT 154.950 199.950 157.050 202.050 ;
        RECT 166.950 199.950 169.050 202.050 ;
        RECT 172.950 200.250 175.050 201.150 ;
        RECT 178.950 199.950 181.050 202.050 ;
        RECT 214.950 200.250 216.750 201.150 ;
        RECT 217.950 199.950 220.050 202.050 ;
        RECT 221.250 200.250 222.750 201.150 ;
        RECT 223.950 199.950 226.050 202.050 ;
        RECT 154.950 196.950 157.050 199.050 ;
        RECT 133.950 194.400 138.450 195.450 ;
        RECT 133.950 193.950 136.050 194.400 ;
        RECT 133.950 191.850 136.050 192.750 ;
        RECT 130.950 187.500 133.050 189.600 ;
        RECT 137.400 163.050 138.450 194.400 ;
        RECT 155.400 166.050 156.450 196.950 ;
        RECT 151.950 164.250 153.750 165.150 ;
        RECT 154.950 163.950 157.050 166.050 ;
        RECT 158.250 164.250 160.050 165.150 ;
        RECT 136.950 160.950 139.050 163.050 ;
        RECT 151.950 160.950 154.050 163.050 ;
        RECT 155.250 161.850 156.750 162.750 ;
        RECT 157.950 160.950 160.050 163.050 ;
        RECT 152.400 130.050 153.450 160.950 ;
        RECT 167.400 130.050 168.450 199.950 ;
        RECT 179.400 199.050 180.450 199.950 ;
        RECT 172.950 196.950 175.050 199.050 ;
        RECT 176.250 197.250 177.750 198.150 ;
        RECT 178.950 196.950 181.050 199.050 ;
        RECT 182.250 197.250 184.050 198.150 ;
        RECT 214.950 196.950 217.050 199.050 ;
        RECT 215.400 196.050 216.450 196.950 ;
        RECT 175.950 193.950 178.050 196.050 ;
        RECT 179.250 194.850 180.750 195.750 ;
        RECT 181.950 193.950 184.050 196.050 ;
        RECT 214.950 193.950 217.050 196.050 ;
        RECT 182.400 172.050 183.450 193.950 ;
        RECT 181.950 169.950 184.050 172.050 ;
        RECT 182.400 166.050 183.450 169.950 ;
        RECT 218.400 169.050 219.450 199.950 ;
        RECT 220.950 196.950 223.050 199.050 ;
        RECT 224.250 197.850 226.050 198.750 ;
        RECT 190.950 167.250 193.050 168.150 ;
        RECT 193.950 167.850 196.050 168.750 ;
        RECT 217.950 166.950 220.050 169.050 ;
        RECT 181.950 163.950 184.050 166.050 ;
        RECT 190.950 163.950 193.050 166.050 ;
        RECT 208.950 163.950 211.050 166.050 ;
        RECT 184.950 130.950 187.050 133.050 ;
        RECT 151.950 127.950 154.050 130.050 ;
        RECT 166.950 127.950 169.050 130.050 ;
        RECT 172.950 128.250 175.050 129.150 ;
        RECT 178.950 127.950 181.050 130.050 ;
        RECT 167.400 127.050 168.450 127.950 ;
        RECT 148.950 124.950 151.050 127.050 ;
        RECT 163.950 125.250 165.750 126.150 ;
        RECT 166.950 124.950 169.050 127.050 ;
        RECT 170.250 125.250 171.750 126.150 ;
        RECT 172.950 124.950 175.050 127.050 ;
        RECT 127.950 121.950 130.050 124.050 ;
        RECT 127.950 119.850 130.050 120.750 ;
        RECT 124.950 115.500 127.050 117.600 ;
        RECT 136.950 101.400 139.050 103.500 ;
        RECT 115.950 94.950 118.050 97.050 ;
        RECT 119.250 95.250 120.750 96.150 ;
        RECT 121.950 94.950 124.050 97.050 ;
        RECT 115.950 92.850 117.750 93.750 ;
        RECT 118.950 91.950 121.050 94.050 ;
        RECT 122.250 92.850 123.750 93.750 ;
        RECT 124.950 91.950 127.050 94.050 ;
        RECT 119.400 91.050 120.450 91.950 ;
        RECT 82.950 89.400 87.450 90.450 ;
        RECT 82.950 88.950 85.050 89.400 ;
        RECT 118.950 88.950 121.050 91.050 ;
        RECT 124.950 89.850 127.050 90.750 ;
        RECT 71.400 58.050 72.450 88.950 ;
        RECT 137.400 84.600 138.600 101.400 ;
        RECT 142.950 100.950 145.050 103.050 ;
        RECT 143.400 97.050 144.450 100.950 ;
        RECT 149.400 100.050 150.450 124.950 ;
        RECT 163.950 121.950 166.050 124.050 ;
        RECT 167.250 122.850 168.750 123.750 ;
        RECT 169.950 121.950 172.050 124.050 ;
        RECT 164.400 112.050 165.450 121.950 ;
        RECT 163.950 109.950 166.050 112.050 ;
        RECT 157.950 101.400 160.050 103.500 ;
        RECT 170.400 103.050 171.450 121.950 ;
        RECT 148.950 97.950 151.050 100.050 ;
        RECT 149.400 97.050 150.450 97.950 ;
        RECT 142.950 94.950 145.050 97.050 ;
        RECT 148.950 94.950 151.050 97.050 ;
        RECT 142.950 92.850 145.050 93.750 ;
        RECT 148.950 92.850 151.050 93.750 ;
        RECT 158.250 89.400 159.450 101.400 ;
        RECT 169.950 100.950 172.050 103.050 ;
        RECT 172.950 101.400 175.050 103.500 ;
        RECT 160.950 98.250 163.050 99.150 ;
        RECT 169.950 98.250 172.050 99.150 ;
        RECT 160.950 94.950 163.050 97.050 ;
        RECT 169.950 94.950 172.050 97.050 ;
        RECT 170.400 94.050 171.450 94.950 ;
        RECT 169.950 91.950 172.050 94.050 ;
        RECT 173.550 89.400 174.750 101.400 ;
        RECT 175.950 97.950 178.050 100.050 ;
        RECT 157.950 87.300 160.050 89.400 ;
        RECT 172.950 87.300 175.050 89.400 ;
        RECT 136.950 82.500 139.050 84.600 ;
        RECT 158.250 83.700 159.450 87.300 ;
        RECT 173.550 83.700 174.750 87.300 ;
        RECT 157.950 81.600 160.050 83.700 ;
        RECT 172.950 81.600 175.050 83.700 ;
        RECT 76.950 59.250 79.050 60.150 ;
        RECT 70.950 55.950 73.050 58.050 ;
        RECT 74.250 56.250 75.750 57.150 ;
        RECT 76.950 55.950 79.050 58.050 ;
        RECT 157.950 57.450 160.050 58.050 ;
        RECT 80.250 56.250 82.050 57.150 ;
        RECT 155.400 56.400 160.050 57.450 ;
        RECT 67.950 52.950 70.050 55.050 ;
        RECT 70.950 53.850 72.750 54.750 ;
        RECT 73.950 52.950 76.050 55.050 ;
        RECT 74.400 52.050 75.450 52.950 ;
        RECT 31.950 51.450 34.050 52.050 ;
        RECT 31.950 50.400 36.450 51.450 ;
        RECT 31.950 49.950 34.050 50.400 ;
        RECT 31.950 47.850 34.050 48.750 ;
        RECT 28.950 43.500 31.050 45.600 ;
        RECT 35.400 28.050 36.450 50.400 ;
        RECT 73.950 49.950 76.050 52.050 ;
        RECT 77.400 46.050 78.450 55.950 ;
        RECT 79.950 52.950 82.050 55.050 ;
        RECT 112.950 53.250 115.050 54.150 ;
        RECT 118.950 53.250 121.050 54.150 ;
        RECT 151.950 53.250 154.050 54.150 ;
        RECT 76.950 43.950 79.050 46.050 ;
        RECT 43.950 29.400 46.050 31.500 ;
        RECT 64.950 29.400 67.050 31.500 ;
        RECT 34.950 25.950 37.050 28.050 ;
        RECT 19.950 22.950 22.050 25.050 ;
        RECT 31.950 23.250 34.050 24.150 ;
        RECT 34.950 23.850 37.050 24.750 ;
        RECT 31.950 19.950 34.050 22.050 ;
        RECT 44.400 12.600 45.600 29.400 ;
        RECT 49.950 25.950 52.050 28.050 ;
        RECT 50.400 25.050 51.450 25.950 ;
        RECT 49.950 22.950 52.050 25.050 ;
        RECT 55.950 22.950 58.050 25.050 ;
        RECT 49.950 20.850 52.050 21.750 ;
        RECT 55.950 20.850 58.050 21.750 ;
        RECT 65.250 17.400 66.450 29.400 ;
        RECT 67.950 26.250 70.050 27.150 ;
        RECT 77.400 25.050 78.450 43.950 ;
        RECT 80.400 25.050 81.450 52.950 ;
        RECT 112.950 49.950 115.050 52.050 ;
        RECT 116.250 50.250 117.750 51.150 ;
        RECT 118.950 49.950 121.050 52.050 ;
        RECT 151.950 49.950 154.050 52.050 ;
        RECT 106.950 28.950 109.050 31.050 ;
        RECT 107.400 28.050 108.450 28.950 ;
        RECT 113.400 28.050 114.450 49.950 ;
        RECT 115.950 46.950 118.050 49.050 ;
        RECT 119.400 46.050 120.450 49.950 ;
        RECT 118.950 43.950 121.050 46.050 ;
        RECT 152.400 28.050 153.450 49.950 ;
        RECT 155.400 49.050 156.450 56.400 ;
        RECT 157.950 55.950 160.050 56.400 ;
        RECT 157.950 53.850 160.050 54.750 ;
        RECT 160.950 53.250 163.050 54.150 ;
        RECT 160.950 49.950 163.050 52.050 ;
        RECT 154.950 46.950 157.050 49.050 ;
        RECT 166.950 43.950 169.050 46.050 ;
        RECT 160.950 29.400 163.050 31.500 ;
        RECT 106.950 25.950 109.050 28.050 ;
        RECT 112.950 25.950 115.050 28.050 ;
        RECT 151.950 25.950 154.050 28.050 ;
        RECT 67.950 22.950 70.050 25.050 ;
        RECT 76.950 22.950 79.050 25.050 ;
        RECT 79.950 22.950 82.050 25.050 ;
        RECT 103.950 22.950 106.050 25.050 ;
        RECT 107.250 23.850 108.750 24.750 ;
        RECT 109.950 24.450 112.050 25.050 ;
        RECT 109.950 23.400 114.450 24.450 ;
        RECT 109.950 22.950 112.050 23.400 ;
        RECT 80.400 22.050 81.450 22.950 ;
        RECT 113.400 22.050 114.450 23.400 ;
        RECT 148.950 23.250 151.050 24.150 ;
        RECT 151.950 23.850 154.050 24.750 ;
        RECT 79.950 19.950 82.050 22.050 ;
        RECT 103.950 20.850 106.050 21.750 ;
        RECT 109.950 20.850 112.050 21.750 ;
        RECT 112.950 19.950 115.050 22.050 ;
        RECT 148.950 19.950 151.050 22.050 ;
        RECT 64.950 15.300 67.050 17.400 ;
        RECT 43.950 10.500 46.050 12.600 ;
        RECT 65.250 11.700 66.450 15.300 ;
        RECT 161.400 12.600 162.600 29.400 ;
        RECT 167.400 25.050 168.450 43.950 ;
        RECT 176.400 25.050 177.450 97.950 ;
        RECT 179.400 55.050 180.450 127.950 ;
        RECT 181.950 97.950 184.050 100.050 ;
        RECT 182.400 97.050 183.450 97.950 ;
        RECT 181.950 94.950 184.050 97.050 ;
        RECT 185.400 94.050 186.450 130.950 ;
        RECT 209.400 130.050 210.450 163.950 ;
        RECT 208.950 127.950 211.050 130.050 ;
        RECT 212.250 128.250 213.750 129.150 ;
        RECT 214.950 127.950 217.050 130.050 ;
        RECT 208.950 125.850 210.750 126.750 ;
        RECT 211.950 124.950 214.050 127.050 ;
        RECT 215.250 125.850 217.050 126.750 ;
        RECT 187.950 100.950 190.050 103.050 ;
        RECT 190.950 100.950 193.050 103.050 ;
        RECT 193.950 101.400 196.050 103.500 ;
        RECT 188.400 97.050 189.450 100.950 ;
        RECT 187.950 94.950 190.050 97.050 ;
        RECT 181.950 92.850 184.050 93.750 ;
        RECT 184.950 91.950 187.050 94.050 ;
        RECT 187.950 92.850 190.050 93.750 ;
        RECT 178.950 52.950 181.050 55.050 ;
        RECT 181.950 29.400 184.050 31.500 ;
        RECT 166.950 22.950 169.050 25.050 ;
        RECT 172.950 24.450 175.050 25.050 ;
        RECT 175.950 24.450 178.050 25.050 ;
        RECT 172.950 23.400 178.050 24.450 ;
        RECT 172.950 22.950 175.050 23.400 ;
        RECT 175.950 22.950 178.050 23.400 ;
        RECT 166.950 20.850 169.050 21.750 ;
        RECT 172.950 20.850 175.050 21.750 ;
        RECT 182.250 17.400 183.450 29.400 ;
        RECT 184.950 26.250 187.050 27.150 ;
        RECT 184.950 22.950 187.050 25.050 ;
        RECT 191.400 24.450 192.450 100.950 ;
        RECT 194.400 84.600 195.600 101.400 ;
        RECT 218.400 100.050 219.450 166.950 ;
        RECT 227.400 166.050 228.450 313.950 ;
        RECT 236.400 310.050 237.450 343.950 ;
        RECT 238.950 340.950 241.050 343.050 ;
        RECT 242.250 341.250 243.750 342.150 ;
        RECT 244.950 340.950 247.050 343.050 ;
        RECT 248.250 341.250 250.050 342.150 ;
        RECT 239.400 337.050 240.450 340.950 ;
        RECT 241.950 337.950 244.050 340.050 ;
        RECT 245.250 338.850 246.750 339.750 ;
        RECT 247.950 339.450 250.050 340.050 ;
        RECT 251.400 339.450 252.450 382.950 ;
        RECT 253.950 340.950 256.050 343.050 ;
        RECT 247.950 338.400 252.450 339.450 ;
        RECT 247.950 337.950 250.050 338.400 ;
        RECT 238.950 334.950 241.050 337.050 ;
        RECT 244.950 310.950 247.050 313.050 ;
        RECT 232.950 308.250 234.750 309.150 ;
        RECT 235.950 307.950 238.050 310.050 ;
        RECT 239.250 308.250 241.050 309.150 ;
        RECT 245.400 307.050 246.450 310.950 ;
        RECT 251.400 307.050 252.450 338.400 ;
        RECT 254.400 313.050 255.450 340.950 ;
        RECT 253.950 310.950 256.050 313.050 ;
        RECT 232.950 304.950 235.050 307.050 ;
        RECT 236.250 305.850 237.750 306.750 ;
        RECT 238.950 304.950 241.050 307.050 ;
        RECT 244.950 304.950 247.050 307.050 ;
        RECT 250.950 304.950 253.050 307.050 ;
        RECT 239.400 283.050 240.450 304.950 ;
        RECT 238.950 280.950 241.050 283.050 ;
        RECT 235.950 274.950 238.050 277.050 ;
        RECT 236.400 274.050 237.450 274.950 ;
        RECT 235.950 271.950 238.050 274.050 ;
        RECT 241.950 273.450 244.050 274.050 ;
        RECT 239.250 272.250 240.750 273.150 ;
        RECT 241.950 272.400 246.450 273.450 ;
        RECT 241.950 271.950 244.050 272.400 ;
        RECT 235.950 269.850 237.750 270.750 ;
        RECT 238.950 268.950 241.050 271.050 ;
        RECT 242.250 269.850 244.050 270.750 ;
        RECT 245.400 255.450 246.450 272.400 ;
        RECT 242.400 254.400 246.450 255.450 ;
        RECT 229.950 238.950 232.050 241.050 ;
        RECT 230.400 196.050 231.450 238.950 ;
        RECT 242.400 199.050 243.450 254.400 ;
        RECT 253.950 241.950 256.050 244.050 ;
        RECT 254.400 238.050 255.450 241.950 ;
        RECT 244.950 236.250 246.750 237.150 ;
        RECT 247.950 235.950 250.050 238.050 ;
        RECT 253.950 235.950 256.050 238.050 ;
        RECT 244.950 232.950 247.050 235.050 ;
        RECT 248.250 233.850 249.750 234.750 ;
        RECT 250.950 232.950 253.050 235.050 ;
        RECT 254.250 233.850 256.050 234.750 ;
        RECT 250.950 230.850 253.050 231.750 ;
        RECT 241.950 196.950 244.050 199.050 ;
        RECT 229.950 193.950 232.050 196.050 ;
        RECT 257.400 195.450 258.450 445.950 ;
        RECT 263.400 409.050 264.450 487.950 ;
        RECT 268.950 485.250 271.050 486.150 ;
        RECT 268.950 481.950 271.050 484.050 ;
        RECT 269.400 478.050 270.450 481.950 ;
        RECT 272.400 478.050 273.450 518.400 ;
        RECT 274.950 487.950 277.050 490.050 ;
        RECT 274.950 485.850 277.050 486.750 ;
        RECT 277.950 485.250 280.050 486.150 ;
        RECT 277.950 483.450 280.050 484.050 ;
        RECT 281.400 483.450 282.450 556.950 ;
        RECT 283.950 553.950 286.050 556.050 ;
        RECT 287.250 554.850 288.750 555.750 ;
        RECT 289.950 553.950 292.050 556.050 ;
        RECT 290.400 523.050 291.450 553.950 ;
        RECT 293.400 553.050 294.450 556.950 ;
        RECT 304.950 553.950 307.050 556.050 ;
        RECT 292.950 550.950 295.050 553.050 ;
        RECT 289.950 520.950 292.050 523.050 ;
        RECT 289.950 494.400 292.050 496.500 ;
        RECT 277.950 482.400 282.450 483.450 ;
        RECT 277.950 481.950 280.050 482.400 ;
        RECT 268.950 475.950 271.050 478.050 ;
        RECT 271.950 475.950 274.050 478.050 ;
        RECT 290.400 477.600 291.600 494.400 ;
        RECT 295.950 485.250 298.050 486.150 ;
        RECT 301.950 485.250 304.050 486.150 ;
        RECT 295.950 481.950 298.050 484.050 ;
        RECT 301.950 481.950 304.050 484.050 ;
        RECT 302.400 481.050 303.450 481.950 ;
        RECT 301.950 478.950 304.050 481.050 ;
        RECT 289.950 475.500 292.050 477.600 ;
        RECT 305.400 460.050 306.450 553.950 ;
        RECT 292.950 457.950 295.050 460.050 ;
        RECT 304.950 457.950 307.050 460.050 ;
        RECT 277.950 451.950 280.050 454.050 ;
        RECT 271.950 448.950 274.050 451.050 ;
        RECT 272.400 415.050 273.450 448.950 ;
        RECT 271.950 412.950 274.050 415.050 ;
        RECT 274.950 412.950 277.050 415.050 ;
        RECT 274.950 410.850 277.050 411.750 ;
        RECT 278.400 411.450 279.450 451.950 ;
        RECT 280.950 413.250 283.050 414.150 ;
        RECT 280.950 411.450 283.050 412.050 ;
        RECT 278.400 410.400 283.050 411.450 ;
        RECT 280.950 409.950 283.050 410.400 ;
        RECT 284.250 410.250 286.050 411.150 ;
        RECT 262.950 406.950 265.050 409.050 ;
        RECT 281.400 382.050 282.450 409.950 ;
        RECT 283.950 406.950 286.050 409.050 ;
        RECT 284.400 388.050 285.450 406.950 ;
        RECT 289.950 388.950 292.050 391.050 ;
        RECT 283.950 385.950 286.050 388.050 ;
        RECT 286.950 385.950 289.050 388.050 ;
        RECT 287.400 382.050 288.450 385.950 ;
        RECT 290.400 385.050 291.450 388.950 ;
        RECT 293.400 387.450 294.450 457.950 ;
        RECT 305.400 457.050 306.450 457.950 ;
        RECT 298.950 454.950 301.050 457.050 ;
        RECT 302.250 455.250 303.750 456.150 ;
        RECT 304.950 454.950 307.050 457.050 ;
        RECT 295.950 451.950 298.050 454.050 ;
        RECT 299.250 452.850 300.750 453.750 ;
        RECT 301.950 451.950 304.050 454.050 ;
        RECT 305.250 452.850 307.050 453.750 ;
        RECT 295.950 449.850 298.050 450.750 ;
        RECT 293.400 386.400 297.450 387.450 ;
        RECT 296.400 385.050 297.450 386.400 ;
        RECT 289.950 382.950 292.050 385.050 ;
        RECT 293.250 383.250 294.750 384.150 ;
        RECT 295.950 382.950 298.050 385.050 ;
        RECT 280.950 379.950 283.050 382.050 ;
        RECT 286.950 379.950 289.050 382.050 ;
        RECT 290.250 380.850 291.750 381.750 ;
        RECT 292.950 379.950 295.050 382.050 ;
        RECT 296.250 380.850 298.050 381.750 ;
        RECT 286.950 377.850 289.050 378.750 ;
        RECT 298.950 350.400 301.050 352.500 ;
        RECT 277.950 346.950 280.050 349.050 ;
        RECT 286.950 346.950 289.050 349.050 ;
        RECT 268.950 334.950 271.050 337.050 ;
        RECT 269.400 315.450 270.450 334.950 ;
        RECT 271.950 315.450 274.050 316.050 ;
        RECT 269.400 314.400 274.050 315.450 ;
        RECT 269.400 283.050 270.450 314.400 ;
        RECT 271.950 313.950 274.050 314.400 ;
        RECT 271.950 311.850 273.750 312.750 ;
        RECT 274.950 310.950 277.050 313.050 ;
        RECT 274.950 308.850 277.050 309.750 ;
        RECT 278.400 309.450 279.450 346.950 ;
        RECT 287.400 346.050 288.450 346.950 ;
        RECT 280.950 343.950 283.050 346.050 ;
        RECT 284.250 344.250 285.750 345.150 ;
        RECT 286.950 343.950 289.050 346.050 ;
        RECT 280.950 341.850 282.750 342.750 ;
        RECT 283.950 340.950 286.050 343.050 ;
        RECT 287.250 341.850 289.050 342.750 ;
        RECT 299.400 333.600 300.600 350.400 ;
        RECT 308.400 343.050 309.450 592.950 ;
        RECT 310.950 527.250 313.050 528.150 ;
        RECT 310.950 523.950 313.050 526.050 ;
        RECT 310.950 495.300 313.050 497.400 ;
        RECT 311.250 491.700 312.450 495.300 ;
        RECT 310.950 489.600 313.050 491.700 ;
        RECT 311.250 477.600 312.450 489.600 ;
        RECT 314.400 484.050 315.450 601.950 ;
        RECT 317.400 594.450 318.450 619.950 ;
        RECT 332.400 604.050 333.450 632.400 ;
        RECT 347.400 631.050 348.450 661.950 ;
        RECT 386.400 637.050 387.450 664.950 ;
        RECT 364.950 634.950 367.050 637.050 ;
        RECT 373.950 634.950 376.050 637.050 ;
        RECT 385.950 634.950 388.050 637.050 ;
        RECT 361.950 631.950 364.050 634.050 ;
        RECT 346.950 628.950 349.050 631.050 ;
        RECT 362.400 628.050 363.450 631.950 ;
        RECT 361.950 625.950 364.050 628.050 ;
        RECT 365.400 627.450 366.450 634.950 ;
        RECT 374.400 634.050 375.450 634.950 ;
        RECT 367.950 631.950 370.050 634.050 ;
        RECT 371.250 632.250 372.750 633.150 ;
        RECT 373.950 631.950 376.050 634.050 ;
        RECT 367.950 629.850 369.750 630.750 ;
        RECT 370.950 628.950 373.050 631.050 ;
        RECT 374.250 629.850 376.050 630.750 ;
        RECT 365.400 626.400 369.450 627.450 ;
        RECT 331.950 601.950 334.050 604.050 ;
        RECT 364.950 601.950 367.050 604.050 ;
        RECT 361.950 599.250 364.050 600.150 ;
        RECT 364.950 599.850 367.050 600.750 ;
        RECT 368.400 598.050 369.450 626.400 ;
        RECT 392.400 600.450 393.450 703.950 ;
        RECT 428.400 703.050 429.450 703.950 ;
        RECT 415.950 700.950 418.050 703.050 ;
        RECT 418.950 701.250 420.750 702.150 ;
        RECT 421.950 700.950 424.050 703.050 ;
        RECT 425.250 701.250 426.750 702.150 ;
        RECT 427.950 700.950 430.050 703.050 ;
        RECT 431.250 701.250 433.050 702.150 ;
        RECT 433.950 700.950 436.050 703.050 ;
        RECT 416.400 699.450 417.450 700.950 ;
        RECT 418.950 699.450 421.050 700.050 ;
        RECT 416.400 698.400 421.050 699.450 ;
        RECT 422.250 698.850 423.750 699.750 ;
        RECT 418.950 697.950 421.050 698.400 ;
        RECT 424.950 697.950 427.050 700.050 ;
        RECT 428.250 698.850 429.750 699.750 ;
        RECT 430.950 699.450 433.050 700.050 ;
        RECT 434.400 699.450 435.450 700.950 ;
        RECT 430.950 698.400 435.450 699.450 ;
        RECT 430.950 697.950 433.050 698.400 ;
        RECT 440.400 693.600 441.600 710.400 ;
        RECT 446.400 706.050 447.450 736.950 ;
        RECT 458.400 732.600 459.600 749.400 ;
        RECT 463.950 742.950 466.050 745.050 ;
        RECT 469.950 744.450 472.050 745.050 ;
        RECT 469.950 743.400 474.450 744.450 ;
        RECT 469.950 742.950 472.050 743.400 ;
        RECT 463.950 740.850 466.050 741.750 ;
        RECT 469.950 740.850 472.050 741.750 ;
        RECT 457.950 730.500 460.050 732.600 ;
        RECT 460.950 711.300 463.050 713.400 ;
        RECT 461.250 707.700 462.450 711.300 ;
        RECT 445.950 703.950 448.050 706.050 ;
        RECT 460.950 705.600 463.050 707.700 ;
        RECT 445.950 701.250 448.050 702.150 ;
        RECT 451.950 701.250 454.050 702.150 ;
        RECT 445.950 697.950 448.050 700.050 ;
        RECT 451.950 697.950 454.050 700.050 ;
        RECT 452.400 694.050 453.450 697.950 ;
        RECT 439.950 691.500 442.050 693.600 ;
        RECT 451.950 691.950 454.050 694.050 ;
        RECT 461.250 693.600 462.450 705.600 ;
        RECT 463.950 699.450 466.050 700.050 ;
        RECT 463.950 698.400 468.450 699.450 ;
        RECT 463.950 697.950 466.050 698.400 ;
        RECT 467.400 697.050 468.450 698.400 ;
        RECT 463.950 695.850 466.050 696.750 ;
        RECT 466.950 694.950 469.050 697.050 ;
        RECT 473.400 694.050 474.450 743.400 ;
        RECT 479.250 737.400 480.450 749.400 ;
        RECT 481.950 746.250 484.050 747.150 ;
        RECT 481.950 742.950 484.050 745.050 ;
        RECT 517.950 744.450 520.050 745.050 ;
        RECT 517.950 743.400 522.450 744.450 ;
        RECT 517.950 742.950 520.050 743.400 ;
        RECT 482.400 739.050 483.450 742.950 ;
        RECT 517.950 740.850 520.050 741.750 ;
        RECT 478.950 735.300 481.050 737.400 ;
        RECT 481.950 736.950 484.050 739.050 ;
        RECT 479.250 731.700 480.450 735.300 ;
        RECT 478.950 729.600 481.050 731.700 ;
        RECT 521.400 706.050 522.450 743.400 ;
        RECT 523.950 740.850 526.050 741.750 ;
        RECT 536.400 732.600 537.600 749.400 ;
        RECT 541.950 744.450 544.050 745.050 ;
        RECT 539.400 743.400 544.050 744.450 ;
        RECT 535.950 730.500 538.050 732.600 ;
        RECT 539.400 712.050 540.450 743.400 ;
        RECT 541.950 742.950 544.050 743.400 ;
        RECT 547.950 744.450 550.050 745.050 ;
        RECT 547.950 743.400 552.450 744.450 ;
        RECT 547.950 742.950 550.050 743.400 ;
        RECT 541.950 740.850 544.050 741.750 ;
        RECT 547.950 740.850 550.050 741.750 ;
        RECT 538.950 709.950 541.050 712.050 ;
        RECT 535.950 706.950 538.050 709.050 ;
        RECT 484.950 703.950 487.050 706.050 ;
        RECT 520.950 703.950 523.050 706.050 ;
        RECT 460.950 691.500 463.050 693.600 ;
        RECT 472.950 691.950 475.050 694.050 ;
        RECT 451.950 688.950 454.050 691.050 ;
        RECT 433.950 673.950 436.050 676.050 ;
        RECT 400.950 670.950 403.050 673.050 ;
        RECT 427.950 670.950 430.050 673.050 ;
        RECT 401.400 631.050 402.450 670.950 ;
        RECT 428.400 670.050 429.450 670.950 ;
        RECT 434.400 670.050 435.450 673.950 ;
        RECT 452.400 673.050 453.450 688.950 ;
        RECT 485.400 676.050 486.450 703.950 ;
        RECT 502.950 700.950 505.050 703.050 ;
        RECT 536.400 702.450 537.450 706.950 ;
        RECT 538.950 704.250 541.050 705.150 ;
        RECT 544.950 703.950 547.050 706.050 ;
        RECT 545.400 703.050 546.450 703.950 ;
        RECT 538.950 702.450 541.050 703.050 ;
        RECT 536.400 701.400 541.050 702.450 ;
        RECT 538.950 700.950 541.050 701.400 ;
        RECT 542.250 701.250 543.750 702.150 ;
        RECT 544.950 700.950 547.050 703.050 ;
        RECT 548.250 701.250 550.050 702.150 ;
        RECT 499.950 698.250 502.050 699.150 ;
        RECT 502.950 698.850 505.050 699.750 ;
        RECT 538.950 699.450 541.050 700.050 ;
        RECT 541.950 699.450 544.050 700.050 ;
        RECT 538.950 698.400 544.050 699.450 ;
        RECT 545.250 698.850 546.750 699.750 ;
        RECT 538.950 697.950 541.050 698.400 ;
        RECT 541.950 697.950 544.050 698.400 ;
        RECT 547.950 697.950 550.050 700.050 ;
        RECT 548.400 697.050 549.450 697.950 ;
        RECT 499.950 694.950 502.050 697.050 ;
        RECT 547.950 694.950 550.050 697.050 ;
        RECT 551.400 694.050 552.450 743.400 ;
        RECT 557.250 737.400 558.450 749.400 ;
        RECT 559.950 746.250 562.050 747.150 ;
        RECT 562.950 745.950 565.050 748.050 ;
        RECT 595.950 745.950 598.050 748.050 ;
        RECT 634.950 745.950 637.050 748.050 ;
        RECT 640.950 745.950 643.050 748.050 ;
        RECT 682.950 745.950 685.050 748.050 ;
        RECT 559.950 744.450 562.050 745.050 ;
        RECT 563.400 744.450 564.450 745.950 ;
        RECT 559.950 743.400 564.450 744.450 ;
        RECT 595.950 743.850 598.050 744.750 ;
        RECT 559.950 742.950 562.050 743.400 ;
        RECT 598.950 743.250 601.050 744.150 ;
        RECT 622.950 742.950 625.050 745.050 ;
        RECT 634.950 743.850 637.050 744.750 ;
        RECT 637.950 743.250 640.050 744.150 ;
        RECT 598.950 739.950 601.050 742.050 ;
        RECT 556.950 735.300 559.050 737.400 ;
        RECT 557.250 731.700 558.450 735.300 ;
        RECT 556.950 729.600 559.050 731.700 ;
        RECT 583.950 704.250 586.050 705.150 ;
        RECT 583.950 700.950 586.050 703.050 ;
        RECT 587.250 701.250 588.750 702.150 ;
        RECT 589.950 700.950 592.050 703.050 ;
        RECT 593.250 701.250 595.050 702.150 ;
        RECT 584.400 696.450 585.450 700.950 ;
        RECT 586.950 697.950 589.050 700.050 ;
        RECT 590.250 698.850 591.750 699.750 ;
        RECT 592.950 697.950 595.050 700.050 ;
        RECT 584.400 695.400 588.450 696.450 ;
        RECT 541.950 691.950 544.050 694.050 ;
        RECT 550.950 691.950 553.050 694.050 ;
        RECT 523.950 677.400 526.050 679.500 ;
        RECT 469.950 673.950 472.050 676.050 ;
        RECT 484.950 673.950 487.050 676.050 ;
        RECT 470.400 673.050 471.450 673.950 ;
        RECT 451.950 670.950 454.050 673.050 ;
        RECT 463.950 670.950 466.050 673.050 ;
        RECT 469.950 670.950 472.050 673.050 ;
        RECT 421.950 667.950 424.050 670.050 ;
        RECT 424.950 668.250 426.750 669.150 ;
        RECT 427.950 667.950 430.050 670.050 ;
        RECT 433.950 667.950 436.050 670.050 ;
        RECT 422.400 664.050 423.450 667.950 ;
        RECT 424.950 664.950 427.050 667.050 ;
        RECT 428.250 665.850 429.750 666.750 ;
        RECT 430.950 664.950 433.050 667.050 ;
        RECT 434.250 665.850 436.050 666.750 ;
        RECT 403.950 661.950 406.050 664.050 ;
        RECT 421.950 661.950 424.050 664.050 ;
        RECT 430.950 662.850 433.050 663.750 ;
        RECT 404.400 634.050 405.450 661.950 ;
        RECT 415.950 635.250 418.050 636.150 ;
        RECT 403.950 631.950 406.050 634.050 ;
        RECT 409.950 633.450 412.050 634.050 ;
        RECT 407.400 632.400 412.050 633.450 ;
        RECT 407.400 631.050 408.450 632.400 ;
        RECT 409.950 631.950 412.050 632.400 ;
        RECT 413.250 632.250 414.750 633.150 ;
        RECT 415.950 631.950 418.050 634.050 ;
        RECT 419.250 632.250 421.050 633.150 ;
        RECT 400.950 628.950 403.050 631.050 ;
        RECT 406.950 628.950 409.050 631.050 ;
        RECT 409.950 629.850 411.750 630.750 ;
        RECT 412.950 628.950 415.050 631.050 ;
        RECT 418.950 628.950 421.050 631.050 ;
        RECT 413.400 628.050 414.450 628.950 ;
        RECT 412.950 625.950 415.050 628.050 ;
        RECT 394.950 600.450 397.050 601.050 ;
        RECT 392.400 599.400 397.050 600.450 ;
        RECT 319.950 596.250 321.750 597.150 ;
        RECT 322.950 595.950 325.050 598.050 ;
        RECT 326.250 596.250 328.050 597.150 ;
        RECT 328.950 595.950 331.050 598.050 ;
        RECT 361.950 595.950 364.050 598.050 ;
        RECT 367.950 595.950 370.050 598.050 ;
        RECT 319.950 594.450 322.050 595.050 ;
        RECT 317.400 593.400 322.050 594.450 ;
        RECT 323.250 593.850 324.750 594.750 ;
        RECT 319.950 592.950 322.050 593.400 ;
        RECT 325.950 592.950 328.050 595.050 ;
        RECT 326.400 589.050 327.450 592.950 ;
        RECT 325.950 586.950 328.050 589.050 ;
        RECT 329.400 564.450 330.450 595.950 ;
        RECT 326.400 563.400 330.450 564.450 ;
        RECT 316.950 556.950 319.050 559.050 ;
        RECT 326.400 558.450 327.450 563.400 ;
        RECT 328.950 560.250 331.050 561.150 ;
        RECT 328.950 558.450 331.050 559.050 ;
        RECT 326.400 557.400 331.050 558.450 ;
        RECT 317.400 553.050 318.450 556.950 ;
        RECT 316.950 550.950 319.050 553.050 ;
        RECT 317.400 529.050 318.450 550.950 ;
        RECT 326.400 532.050 327.450 557.400 ;
        RECT 328.950 556.950 331.050 557.400 ;
        RECT 332.250 557.250 333.750 558.150 ;
        RECT 334.950 556.950 337.050 559.050 ;
        RECT 338.250 557.250 340.050 558.150 ;
        RECT 331.950 553.950 334.050 556.050 ;
        RECT 335.250 554.850 336.750 555.750 ;
        RECT 337.950 553.950 340.050 556.050 ;
        RECT 332.400 553.050 333.450 553.950 ;
        RECT 331.950 550.950 334.050 553.050 ;
        RECT 319.950 529.950 322.050 532.050 ;
        RECT 325.950 529.950 328.050 532.050 ;
        RECT 316.950 526.950 319.050 529.050 ;
        RECT 320.250 527.850 322.050 528.750 ;
        RECT 352.950 526.950 355.050 529.050 ;
        RECT 353.400 526.050 354.450 526.950 ;
        RECT 316.950 524.850 319.050 525.750 ;
        RECT 352.950 523.950 355.050 526.050 ;
        RECT 358.950 523.950 361.050 526.050 ;
        RECT 362.250 524.250 364.050 525.150 ;
        RECT 352.950 521.850 354.750 522.750 ;
        RECT 355.950 520.950 358.050 523.050 ;
        RECT 359.250 521.850 360.750 522.750 ;
        RECT 361.950 520.950 364.050 523.050 ;
        RECT 355.950 518.850 358.050 519.750 ;
        RECT 352.950 488.250 355.050 489.150 ;
        RECT 358.950 487.950 361.050 490.050 ;
        RECT 359.400 487.050 360.450 487.950 ;
        RECT 352.950 484.950 355.050 487.050 ;
        RECT 356.250 485.250 357.750 486.150 ;
        RECT 358.950 484.950 361.050 487.050 ;
        RECT 362.250 485.250 364.050 486.150 ;
        RECT 313.950 481.950 316.050 484.050 ;
        RECT 313.950 479.850 316.050 480.750 ;
        RECT 353.400 478.050 354.450 484.950 ;
        RECT 368.400 484.050 369.450 595.950 ;
        RECT 373.950 557.250 376.050 558.150 ;
        RECT 379.950 556.950 382.050 559.050 ;
        RECT 370.950 554.250 372.750 555.150 ;
        RECT 373.950 553.950 376.050 556.050 ;
        RECT 379.950 554.850 382.050 555.750 ;
        RECT 370.950 550.950 373.050 553.050 ;
        RECT 374.400 550.050 375.450 553.950 ;
        RECT 373.950 547.950 376.050 550.050 ;
        RECT 374.400 520.050 375.450 547.950 ;
        RECT 392.400 541.050 393.450 599.400 ;
        RECT 394.950 598.950 397.050 599.400 ;
        RECT 398.250 599.250 399.750 600.150 ;
        RECT 400.950 598.950 403.050 601.050 ;
        RECT 394.950 596.850 396.750 597.750 ;
        RECT 397.950 595.950 400.050 598.050 ;
        RECT 401.250 596.850 402.750 597.750 ;
        RECT 403.950 595.950 406.050 598.050 ;
        RECT 442.950 596.250 444.750 597.150 ;
        RECT 445.950 595.950 448.050 598.050 ;
        RECT 449.250 596.250 451.050 597.150 ;
        RECT 398.400 595.050 399.450 595.950 ;
        RECT 397.950 592.950 400.050 595.050 ;
        RECT 403.950 593.850 406.050 594.750 ;
        RECT 442.950 592.950 445.050 595.050 ;
        RECT 446.250 593.850 447.750 594.750 ;
        RECT 448.950 592.950 451.050 595.050 ;
        RECT 443.400 562.050 444.450 592.950 ;
        RECT 421.950 559.950 424.050 562.050 ;
        RECT 442.950 559.950 445.050 562.050 ;
        RECT 422.400 559.050 423.450 559.950 ;
        RECT 415.950 558.450 418.050 559.050 ;
        RECT 413.400 557.400 418.050 558.450 ;
        RECT 413.400 553.050 414.450 557.400 ;
        RECT 415.950 556.950 418.050 557.400 ;
        RECT 421.950 556.950 424.050 559.050 ;
        RECT 425.250 557.250 427.050 558.150 ;
        RECT 415.950 554.850 418.050 555.750 ;
        RECT 418.950 554.250 421.050 555.150 ;
        RECT 421.950 554.850 423.750 555.750 ;
        RECT 424.950 553.950 427.050 556.050 ;
        RECT 412.950 550.950 415.050 553.050 ;
        RECT 418.950 550.950 421.050 553.050 ;
        RECT 419.400 550.050 420.450 550.950 ;
        RECT 418.950 547.950 421.050 550.050 ;
        RECT 391.950 538.950 394.050 541.050 ;
        RECT 448.950 538.950 451.050 541.050 ;
        RECT 449.400 529.050 450.450 538.950 ;
        RECT 403.950 526.950 406.050 529.050 ;
        RECT 409.950 528.450 412.050 529.050 ;
        RECT 442.950 528.450 445.050 529.050 ;
        RECT 407.250 527.250 408.750 528.150 ;
        RECT 409.950 527.400 414.450 528.450 ;
        RECT 409.950 526.950 412.050 527.400 ;
        RECT 413.400 526.050 414.450 527.400 ;
        RECT 442.950 527.400 447.450 528.450 ;
        RECT 442.950 526.950 445.050 527.400 ;
        RECT 400.950 525.450 403.050 526.050 ;
        RECT 398.400 524.400 403.050 525.450 ;
        RECT 404.250 524.850 405.750 525.750 ;
        RECT 398.400 523.050 399.450 524.400 ;
        RECT 400.950 523.950 403.050 524.400 ;
        RECT 406.950 523.950 409.050 526.050 ;
        RECT 410.250 524.850 412.050 525.750 ;
        RECT 412.950 523.950 415.050 526.050 ;
        RECT 442.950 524.850 445.050 525.750 ;
        RECT 397.950 520.950 400.050 523.050 ;
        RECT 400.950 521.850 403.050 522.750 ;
        RECT 373.950 517.950 376.050 520.050 ;
        RECT 382.950 493.950 385.050 496.050 ;
        RECT 370.950 484.950 373.050 487.050 ;
        RECT 355.950 481.950 358.050 484.050 ;
        RECT 359.250 482.850 360.750 483.750 ;
        RECT 361.950 481.950 364.050 484.050 ;
        RECT 367.950 481.950 370.050 484.050 ;
        RECT 371.400 481.050 372.450 484.950 ;
        RECT 370.950 478.950 373.050 481.050 ;
        RECT 310.950 475.500 313.050 477.600 ;
        RECT 313.950 475.950 316.050 478.050 ;
        RECT 352.950 475.950 355.050 478.050 ;
        RECT 314.400 460.050 315.450 475.950 ;
        RECT 355.950 461.400 358.050 463.500 ;
        RECT 313.950 457.950 316.050 460.050 ;
        RECT 343.950 457.950 346.050 460.050 ;
        RECT 310.950 454.950 313.050 457.050 ;
        RECT 311.400 418.050 312.450 454.950 ;
        RECT 314.400 454.050 315.450 457.950 ;
        RECT 340.950 454.950 343.050 457.050 ;
        RECT 344.250 455.850 345.750 456.750 ;
        RECT 346.950 456.450 349.050 457.050 ;
        RECT 346.950 455.400 351.450 456.450 ;
        RECT 346.950 454.950 349.050 455.400 ;
        RECT 313.950 451.950 316.050 454.050 ;
        RECT 340.950 452.850 343.050 453.750 ;
        RECT 343.950 451.950 346.050 454.050 ;
        RECT 346.950 452.850 349.050 453.750 ;
        RECT 340.950 445.950 343.050 448.050 ;
        RECT 322.950 421.950 325.050 424.050 ;
        RECT 316.950 419.250 319.050 420.150 ;
        RECT 323.400 418.050 324.450 421.950 ;
        RECT 310.950 415.950 313.050 418.050 ;
        RECT 313.950 416.250 315.750 417.150 ;
        RECT 316.950 415.950 319.050 418.050 ;
        RECT 320.250 416.250 321.750 417.150 ;
        RECT 322.950 415.950 325.050 418.050 ;
        RECT 313.950 412.950 316.050 415.050 ;
        RECT 319.950 412.950 322.050 415.050 ;
        RECT 323.250 413.850 325.050 414.750 ;
        RECT 314.400 412.050 315.450 412.950 ;
        RECT 313.950 409.950 316.050 412.050 ;
        RECT 313.950 394.950 316.050 397.050 ;
        RECT 304.950 341.250 307.050 342.150 ;
        RECT 307.950 340.950 310.050 343.050 ;
        RECT 310.950 341.250 313.050 342.150 ;
        RECT 304.950 337.950 307.050 340.050 ;
        RECT 310.950 339.450 313.050 340.050 ;
        RECT 314.400 339.450 315.450 394.950 ;
        RECT 331.950 385.950 334.050 388.050 ;
        RECT 332.400 385.050 333.450 385.950 ;
        RECT 331.950 382.950 334.050 385.050 ;
        RECT 337.950 384.450 340.050 385.050 ;
        RECT 341.400 384.450 342.450 445.950 ;
        RECT 335.250 383.250 336.750 384.150 ;
        RECT 337.950 383.400 342.450 384.450 ;
        RECT 337.950 382.950 340.050 383.400 ;
        RECT 328.950 381.450 331.050 382.050 ;
        RECT 326.400 380.400 331.050 381.450 ;
        RECT 332.250 380.850 333.750 381.750 ;
        RECT 319.950 351.300 322.050 353.400 ;
        RECT 320.250 347.700 321.450 351.300 ;
        RECT 319.950 345.600 322.050 347.700 ;
        RECT 310.950 338.400 315.450 339.450 ;
        RECT 310.950 337.950 313.050 338.400 ;
        RECT 305.400 334.050 306.450 337.950 ;
        RECT 298.950 331.500 301.050 333.600 ;
        RECT 304.950 331.950 307.050 334.050 ;
        RECT 320.250 333.600 321.450 345.600 ;
        RECT 322.950 340.950 325.050 343.050 ;
        RECT 323.400 340.050 324.450 340.950 ;
        RECT 322.950 337.950 325.050 340.050 ;
        RECT 322.950 335.850 325.050 336.750 ;
        RECT 319.950 331.500 322.050 333.600 ;
        RECT 322.950 331.950 325.050 334.050 ;
        RECT 313.950 319.950 316.050 322.050 ;
        RECT 304.950 313.950 307.050 316.050 ;
        RECT 280.950 311.250 283.050 312.150 ;
        RECT 280.950 309.450 283.050 310.050 ;
        RECT 278.400 308.400 283.050 309.450 ;
        RECT 280.950 307.950 283.050 308.400 ;
        RECT 268.950 280.950 271.050 283.050 ;
        RECT 274.950 280.950 277.050 283.050 ;
        RECT 265.950 235.950 268.050 238.050 ;
        RECT 259.950 232.950 262.050 235.050 ;
        RECT 260.400 202.050 261.450 232.950 ;
        RECT 266.400 202.050 267.450 235.950 ;
        RECT 259.950 199.950 262.050 202.050 ;
        RECT 263.250 200.250 264.750 201.150 ;
        RECT 265.950 199.950 268.050 202.050 ;
        RECT 259.950 197.850 261.750 198.750 ;
        RECT 262.950 196.950 265.050 199.050 ;
        RECT 266.250 197.850 268.050 198.750 ;
        RECT 257.400 194.400 261.450 195.450 ;
        RECT 230.400 166.050 231.450 193.950 ;
        RECT 232.950 166.950 235.050 169.050 ;
        RECT 238.950 168.450 241.050 169.050 ;
        RECT 236.250 167.250 237.750 168.150 ;
        RECT 238.950 167.400 243.450 168.450 ;
        RECT 238.950 166.950 241.050 167.400 ;
        RECT 226.950 163.950 229.050 166.050 ;
        RECT 229.950 163.950 232.050 166.050 ;
        RECT 233.250 164.850 234.750 165.750 ;
        RECT 235.950 163.950 238.050 166.050 ;
        RECT 239.250 164.850 241.050 165.750 ;
        RECT 227.400 118.050 228.450 163.950 ;
        RECT 242.400 163.050 243.450 167.400 ;
        RECT 229.950 161.850 232.050 162.750 ;
        RECT 241.950 160.950 244.050 163.050 ;
        RECT 242.400 124.050 243.450 160.950 ;
        RECT 250.950 125.250 253.050 126.150 ;
        RECT 256.950 125.250 259.050 126.150 ;
        RECT 235.950 121.950 238.050 124.050 ;
        RECT 241.950 121.950 244.050 124.050 ;
        RECT 250.950 121.950 253.050 124.050 ;
        RECT 254.250 122.250 255.750 123.150 ;
        RECT 256.950 121.950 259.050 124.050 ;
        RECT 226.950 115.950 229.050 118.050 ;
        RECT 217.950 97.950 220.050 100.050 ;
        RECT 227.400 97.050 228.450 115.950 ;
        RECT 229.950 97.950 232.050 100.050 ;
        RECT 232.950 97.950 235.050 100.050 ;
        RECT 230.400 97.050 231.450 97.950 ;
        RECT 236.400 97.050 237.450 121.950 ;
        RECT 253.950 118.950 256.050 121.050 ;
        RECT 257.400 118.050 258.450 121.950 ;
        RECT 256.950 115.950 259.050 118.050 ;
        RECT 238.950 100.950 241.050 103.050 ;
        RECT 226.950 94.950 229.050 97.050 ;
        RECT 229.950 94.950 232.050 97.050 ;
        RECT 233.250 95.850 234.750 96.750 ;
        RECT 235.950 94.950 238.050 97.050 ;
        RECT 229.950 92.850 232.050 93.750 ;
        RECT 235.950 92.850 238.050 93.750 ;
        RECT 193.950 82.500 196.050 84.600 ;
        RECT 239.400 58.050 240.450 100.950 ;
        RECT 196.950 55.950 199.050 58.050 ;
        RECT 202.950 57.450 205.050 58.050 ;
        RECT 200.250 56.250 201.750 57.150 ;
        RECT 202.950 56.400 207.450 57.450 ;
        RECT 202.950 55.950 205.050 56.400 ;
        RECT 196.950 53.850 198.750 54.750 ;
        RECT 199.950 52.950 202.050 55.050 ;
        RECT 203.250 53.850 205.050 54.750 ;
        RECT 206.400 52.050 207.450 56.400 ;
        RECT 211.950 55.950 214.050 58.050 ;
        RECT 238.950 55.950 241.050 58.050 ;
        RECT 244.950 57.450 247.050 58.050 ;
        RECT 242.250 56.250 243.750 57.150 ;
        RECT 244.950 56.400 249.450 57.450 ;
        RECT 244.950 55.950 247.050 56.400 ;
        RECT 205.950 49.950 208.050 52.050 ;
        RECT 196.950 29.400 199.050 31.500 ;
        RECT 193.950 26.250 196.050 27.150 ;
        RECT 193.950 24.450 196.050 25.050 ;
        RECT 191.400 23.400 196.050 24.450 ;
        RECT 193.950 22.950 196.050 23.400 ;
        RECT 185.400 22.050 186.450 22.950 ;
        RECT 184.950 19.950 187.050 22.050 ;
        RECT 197.550 17.400 198.750 29.400 ;
        RECT 212.400 25.050 213.450 55.950 ;
        RECT 238.950 53.850 240.750 54.750 ;
        RECT 241.950 52.950 244.050 55.050 ;
        RECT 245.250 53.850 247.050 54.750 ;
        RECT 242.400 49.050 243.450 52.950 ;
        RECT 248.400 52.050 249.450 56.400 ;
        RECT 247.950 49.950 250.050 52.050 ;
        RECT 241.950 46.950 244.050 49.050 ;
        RECT 217.950 29.400 220.050 31.500 ;
        RECT 260.400 31.050 261.450 194.400 ;
        RECT 275.400 169.050 276.450 280.950 ;
        RECT 280.950 275.250 283.050 276.150 ;
        RECT 277.950 272.250 279.750 273.150 ;
        RECT 280.950 271.950 283.050 274.050 ;
        RECT 286.950 273.450 289.050 274.050 ;
        RECT 284.250 272.250 285.750 273.150 ;
        RECT 286.950 272.400 291.450 273.450 ;
        RECT 286.950 271.950 289.050 272.400 ;
        RECT 277.950 268.950 280.050 271.050 ;
        RECT 278.400 196.050 279.450 268.950 ;
        RECT 281.400 265.050 282.450 271.950 ;
        RECT 283.950 268.950 286.050 271.050 ;
        RECT 287.250 269.850 289.050 270.750 ;
        RECT 290.400 265.050 291.450 272.400 ;
        RECT 280.950 262.950 283.050 265.050 ;
        RECT 289.950 262.950 292.050 265.050 ;
        RECT 286.950 244.950 289.050 247.050 ;
        RECT 287.400 241.050 288.450 244.950 ;
        RECT 286.950 238.950 289.050 241.050 ;
        RECT 292.950 238.950 295.050 241.050 ;
        RECT 286.950 236.850 289.050 237.750 ;
        RECT 289.950 235.950 292.050 238.050 ;
        RECT 292.950 236.850 295.050 237.750 ;
        RECT 280.950 199.950 283.050 202.050 ;
        RECT 277.950 193.950 280.050 196.050 ;
        RECT 268.950 166.950 271.050 169.050 ;
        RECT 274.950 166.950 277.050 169.050 ;
        RECT 269.400 166.050 270.450 166.950 ;
        RECT 275.400 166.050 276.450 166.950 ;
        RECT 268.950 163.950 271.050 166.050 ;
        RECT 274.950 163.950 277.050 166.050 ;
        RECT 278.250 164.250 280.050 165.150 ;
        RECT 268.950 161.850 270.750 162.750 ;
        RECT 271.950 160.950 274.050 163.050 ;
        RECT 275.250 161.850 276.750 162.750 ;
        RECT 277.950 160.950 280.050 163.050 ;
        RECT 271.950 158.850 274.050 159.750 ;
        RECT 274.950 157.950 277.050 160.050 ;
        RECT 275.400 127.050 276.450 157.950 ;
        RECT 274.950 124.950 277.050 127.050 ;
        RECT 271.950 112.950 274.050 115.050 ;
        RECT 272.400 97.050 273.450 112.950 ;
        RECT 277.950 97.950 280.050 100.050 ;
        RECT 271.950 94.950 274.050 97.050 ;
        RECT 271.950 92.850 274.050 93.750 ;
        RECT 274.950 92.250 277.050 93.150 ;
        RECT 274.950 90.450 277.050 91.050 ;
        RECT 278.400 90.450 279.450 97.950 ;
        RECT 281.400 97.050 282.450 199.950 ;
        RECT 290.400 151.050 291.450 235.950 ;
        RECT 301.950 197.250 304.050 198.150 ;
        RECT 301.950 195.450 304.050 196.050 ;
        RECT 305.400 195.450 306.450 313.950 ;
        RECT 314.400 274.050 315.450 319.950 ;
        RECT 323.400 313.050 324.450 331.950 ;
        RECT 326.400 319.050 327.450 380.400 ;
        RECT 328.950 379.950 331.050 380.400 ;
        RECT 334.950 379.950 337.050 382.050 ;
        RECT 338.250 380.850 340.050 381.750 ;
        RECT 328.950 377.850 331.050 378.750 ;
        RECT 335.400 343.050 336.450 379.950 ;
        RECT 334.950 340.950 337.050 343.050 ;
        RECT 341.400 337.050 342.450 383.400 ;
        RECT 344.400 382.050 345.450 451.950 ;
        RECT 350.400 448.050 351.450 455.400 ;
        RECT 349.950 445.950 352.050 448.050 ;
        RECT 356.400 444.600 357.600 461.400 ;
        RECT 361.950 456.450 364.050 457.050 ;
        RECT 359.400 455.400 364.050 456.450 ;
        RECT 359.400 451.050 360.450 455.400 ;
        RECT 361.950 454.950 364.050 455.400 ;
        RECT 367.950 456.450 370.050 457.050 ;
        RECT 371.400 456.450 372.450 478.950 ;
        RECT 376.950 461.400 379.050 463.500 ;
        RECT 383.400 463.050 384.450 493.950 ;
        RECT 394.950 482.850 397.050 483.750 ;
        RECT 407.400 475.050 408.450 523.950 ;
        RECT 427.950 487.950 430.050 490.050 ;
        RECT 415.950 484.950 418.050 487.050 ;
        RECT 415.950 482.850 418.050 483.750 ;
        RECT 415.950 475.950 418.050 478.050 ;
        RECT 406.950 472.950 409.050 475.050 ;
        RECT 367.950 455.400 372.450 456.450 ;
        RECT 367.950 454.950 370.050 455.400 ;
        RECT 361.950 452.850 364.050 453.750 ;
        RECT 367.950 452.850 370.050 453.750 ;
        RECT 358.950 448.950 361.050 451.050 ;
        RECT 355.950 442.500 358.050 444.600 ;
        RECT 355.950 417.450 358.050 418.050 ;
        RECT 353.400 416.400 358.050 417.450 ;
        RECT 361.950 417.450 364.050 418.050 ;
        RECT 353.400 406.050 354.450 416.400 ;
        RECT 355.950 415.950 358.050 416.400 ;
        RECT 359.250 416.250 360.750 417.150 ;
        RECT 361.950 416.400 366.450 417.450 ;
        RECT 361.950 415.950 364.050 416.400 ;
        RECT 355.950 413.850 357.750 414.750 ;
        RECT 358.950 412.950 361.050 415.050 ;
        RECT 362.250 413.850 364.050 414.750 ;
        RECT 352.950 403.950 355.050 406.050 ;
        RECT 365.400 391.050 366.450 416.400 ;
        RECT 371.400 397.050 372.450 455.400 ;
        RECT 377.250 449.400 378.450 461.400 ;
        RECT 382.950 460.950 385.050 463.050 ;
        RECT 379.950 458.250 382.050 459.150 ;
        RECT 379.950 456.450 382.050 457.050 ;
        RECT 383.400 456.450 384.450 460.950 ;
        RECT 379.950 455.400 384.450 456.450 ;
        RECT 379.950 454.950 382.050 455.400 ;
        RECT 416.400 454.050 417.450 475.950 ;
        RECT 412.950 452.250 414.750 453.150 ;
        RECT 415.950 451.950 418.050 454.050 ;
        RECT 419.250 452.250 421.050 453.150 ;
        RECT 428.400 451.050 429.450 487.950 ;
        RECT 446.400 484.050 447.450 527.400 ;
        RECT 448.950 526.950 451.050 529.050 ;
        RECT 448.950 524.850 451.050 525.750 ;
        RECT 445.950 481.950 448.050 484.050 ;
        RECT 452.400 457.050 453.450 670.950 ;
        RECT 485.400 670.050 486.450 673.950 ;
        RECT 505.950 670.950 508.050 673.050 ;
        RECT 508.950 670.950 511.050 673.050 ;
        RECT 514.950 672.450 517.050 673.050 ;
        RECT 512.250 671.250 513.750 672.150 ;
        RECT 514.950 671.400 519.450 672.450 ;
        RECT 514.950 670.950 517.050 671.400 ;
        RECT 506.400 670.050 507.450 670.950 ;
        RECT 518.400 670.050 519.450 671.400 ;
        RECT 463.950 668.850 466.050 669.750 ;
        RECT 469.950 668.850 472.050 669.750 ;
        RECT 484.950 667.950 487.050 670.050 ;
        RECT 505.950 667.950 508.050 670.050 ;
        RECT 509.250 668.850 510.750 669.750 ;
        RECT 511.950 667.950 514.050 670.050 ;
        RECT 515.250 668.850 517.050 669.750 ;
        RECT 517.950 667.950 520.050 670.050 ;
        RECT 505.950 665.850 508.050 666.750 ;
        RECT 484.950 646.950 487.050 649.050 ;
        RECT 454.950 628.950 457.050 631.050 ;
        RECT 454.950 626.850 457.050 627.750 ;
        RECT 457.950 626.250 460.050 627.150 ;
        RECT 457.950 622.950 460.050 625.050 ;
        RECT 457.950 605.400 460.050 607.500 ;
        RECT 478.950 605.400 481.050 607.500 ;
        RECT 458.400 588.600 459.600 605.400 ;
        RECT 463.950 598.950 466.050 601.050 ;
        RECT 469.950 598.950 472.050 601.050 ;
        RECT 463.950 596.850 466.050 597.750 ;
        RECT 469.950 596.850 472.050 597.750 ;
        RECT 479.250 593.400 480.450 605.400 ;
        RECT 481.950 602.250 484.050 603.150 ;
        RECT 481.950 600.450 484.050 601.050 ;
        RECT 485.400 600.450 486.450 646.950 ;
        RECT 490.950 634.950 493.050 637.050 ;
        RECT 491.400 634.050 492.450 634.950 ;
        RECT 490.950 631.950 493.050 634.050 ;
        RECT 496.950 633.450 499.050 634.050 ;
        RECT 494.250 632.250 495.750 633.150 ;
        RECT 496.950 632.400 501.450 633.450 ;
        RECT 496.950 631.950 499.050 632.400 ;
        RECT 490.950 629.850 492.750 630.750 ;
        RECT 493.950 628.950 496.050 631.050 ;
        RECT 497.250 629.850 499.050 630.750 ;
        RECT 500.400 625.050 501.450 632.400 ;
        RECT 512.400 631.050 513.450 667.950 ;
        RECT 524.400 660.600 525.600 677.400 ;
        RECT 542.400 673.050 543.450 691.950 ;
        RECT 544.950 677.400 547.050 679.500 ;
        RECT 529.950 670.950 532.050 673.050 ;
        RECT 535.950 670.950 538.050 673.050 ;
        RECT 541.950 670.950 544.050 673.050 ;
        RECT 529.950 668.850 532.050 669.750 ;
        RECT 535.950 668.850 538.050 669.750 ;
        RECT 523.950 658.500 526.050 660.600 ;
        RECT 532.950 635.250 535.050 636.150 ;
        RECT 538.950 634.950 541.050 637.050 ;
        RECT 539.400 634.050 540.450 634.950 ;
        RECT 523.950 631.950 526.050 634.050 ;
        RECT 529.950 632.250 531.750 633.150 ;
        RECT 532.950 631.950 535.050 634.050 ;
        RECT 536.250 632.250 537.750 633.150 ;
        RECT 538.950 631.950 541.050 634.050 ;
        RECT 508.950 628.950 511.050 631.050 ;
        RECT 511.950 628.950 514.050 631.050 ;
        RECT 509.400 628.050 510.450 628.950 ;
        RECT 508.950 625.950 511.050 628.050 ;
        RECT 499.950 622.950 502.050 625.050 ;
        RECT 481.950 599.400 486.450 600.450 ;
        RECT 481.950 598.950 484.050 599.400 ;
        RECT 482.400 595.050 483.450 598.950 ;
        RECT 478.950 591.300 481.050 593.400 ;
        RECT 481.950 592.950 484.050 595.050 ;
        RECT 457.950 586.500 460.050 588.600 ;
        RECT 479.250 587.700 480.450 591.300 ;
        RECT 478.950 585.600 481.050 587.700 ;
        RECT 481.950 566.400 484.050 568.500 ;
        RECT 469.950 559.950 472.050 562.050 ;
        RECT 478.950 559.950 481.050 562.050 ;
        RECT 470.400 559.050 471.450 559.950 ;
        RECT 457.950 556.950 460.050 559.050 ;
        RECT 460.950 557.250 462.750 558.150 ;
        RECT 463.950 556.950 466.050 559.050 ;
        RECT 467.250 557.250 468.750 558.150 ;
        RECT 469.950 556.950 472.050 559.050 ;
        RECT 473.250 557.250 475.050 558.150 ;
        RECT 475.950 556.950 478.050 559.050 ;
        RECT 458.400 555.450 459.450 556.950 ;
        RECT 460.950 555.450 463.050 556.050 ;
        RECT 458.400 554.400 463.050 555.450 ;
        RECT 464.250 554.850 465.750 555.750 ;
        RECT 460.950 553.950 463.050 554.400 ;
        RECT 466.950 553.950 469.050 556.050 ;
        RECT 470.250 554.850 471.750 555.750 ;
        RECT 472.950 555.450 475.050 556.050 ;
        RECT 476.400 555.450 477.450 556.950 ;
        RECT 472.950 554.400 477.450 555.450 ;
        RECT 472.950 553.950 475.050 554.400 ;
        RECT 460.950 533.400 463.050 535.500 ;
        RECT 461.400 516.600 462.600 533.400 ;
        RECT 472.950 529.950 475.050 532.050 ;
        RECT 473.400 529.050 474.450 529.950 ;
        RECT 466.950 526.950 469.050 529.050 ;
        RECT 472.950 526.950 475.050 529.050 ;
        RECT 466.950 524.850 469.050 525.750 ;
        RECT 472.950 524.850 475.050 525.750 ;
        RECT 460.950 514.500 463.050 516.600 ;
        RECT 479.400 490.050 480.450 559.950 ;
        RECT 482.400 549.600 483.600 566.400 ;
        RECT 487.950 557.250 490.050 558.150 ;
        RECT 493.950 557.250 496.050 558.150 ;
        RECT 487.950 553.950 490.050 556.050 ;
        RECT 493.950 553.950 496.050 556.050 ;
        RECT 481.950 547.500 484.050 549.600 ;
        RECT 481.950 533.400 484.050 535.500 ;
        RECT 482.250 521.400 483.450 533.400 ;
        RECT 494.400 532.050 495.450 553.950 ;
        RECT 484.950 530.250 487.050 531.150 ;
        RECT 493.950 529.950 496.050 532.050 ;
        RECT 484.950 526.950 487.050 529.050 ;
        RECT 494.400 523.050 495.450 529.950 ;
        RECT 481.950 519.300 484.050 521.400 ;
        RECT 493.950 520.950 496.050 523.050 ;
        RECT 482.250 515.700 483.450 519.300 ;
        RECT 500.400 517.050 501.450 622.950 ;
        RECT 524.400 598.050 525.450 631.950 ;
        RECT 529.950 628.950 532.050 631.050 ;
        RECT 533.400 628.050 534.450 631.950 ;
        RECT 535.950 628.950 538.050 631.050 ;
        RECT 539.250 629.850 541.050 630.750 ;
        RECT 536.400 628.050 537.450 628.950 ;
        RECT 532.950 625.950 535.050 628.050 ;
        RECT 535.950 625.950 538.050 628.050 ;
        RECT 535.950 605.400 538.050 607.500 ;
        RECT 529.950 601.950 532.050 604.050 ;
        RECT 532.950 602.250 535.050 603.150 ;
        RECT 530.400 600.450 531.450 601.950 ;
        RECT 532.950 600.450 535.050 601.050 ;
        RECT 530.400 599.400 535.050 600.450 ;
        RECT 520.950 596.250 522.750 597.150 ;
        RECT 523.950 595.950 526.050 598.050 ;
        RECT 527.250 596.250 529.050 597.150 ;
        RECT 520.950 592.950 523.050 595.050 ;
        RECT 524.250 593.850 525.750 594.750 ;
        RECT 526.950 594.450 529.050 595.050 ;
        RECT 530.400 594.450 531.450 599.400 ;
        RECT 532.950 598.950 535.050 599.400 ;
        RECT 526.950 593.400 531.450 594.450 ;
        RECT 536.550 593.400 537.750 605.400 ;
        RECT 542.400 601.050 543.450 670.950 ;
        RECT 545.250 665.400 546.450 677.400 ;
        RECT 547.950 674.250 550.050 675.150 ;
        RECT 550.950 673.950 553.050 676.050 ;
        RECT 580.950 673.950 583.050 676.050 ;
        RECT 547.950 672.450 550.050 673.050 ;
        RECT 551.400 672.450 552.450 673.950 ;
        RECT 547.950 671.400 552.450 672.450 ;
        RECT 580.950 671.850 583.050 672.750 ;
        RECT 547.950 670.950 550.050 671.400 ;
        RECT 583.950 671.250 586.050 672.150 ;
        RECT 583.950 667.950 586.050 670.050 ;
        RECT 544.950 663.300 547.050 665.400 ;
        RECT 545.250 659.700 546.450 663.300 ;
        RECT 544.950 657.600 547.050 659.700 ;
        RECT 577.950 634.950 580.050 637.050 ;
        RECT 578.400 634.050 579.450 634.950 ;
        RECT 577.950 631.950 580.050 634.050 ;
        RECT 581.250 632.250 582.750 633.150 ;
        RECT 583.950 631.950 586.050 634.050 ;
        RECT 577.950 629.850 579.750 630.750 ;
        RECT 580.950 628.950 583.050 631.050 ;
        RECT 584.250 629.850 586.050 630.750 ;
        RECT 581.400 616.050 582.450 628.950 ;
        RECT 550.950 613.950 553.050 616.050 ;
        RECT 580.950 613.950 583.050 616.050 ;
        RECT 551.400 601.050 552.450 613.950 ;
        RECT 556.950 605.400 559.050 607.500 ;
        RECT 541.950 598.950 544.050 601.050 ;
        RECT 544.950 600.450 547.050 601.050 ;
        RECT 544.950 599.400 549.450 600.450 ;
        RECT 544.950 598.950 547.050 599.400 ;
        RECT 544.950 596.850 547.050 597.750 ;
        RECT 526.950 592.950 529.050 593.400 ;
        RECT 502.950 567.300 505.050 569.400 ;
        RECT 503.250 563.700 504.450 567.300 ;
        RECT 502.950 561.600 505.050 563.700 ;
        RECT 521.400 562.050 522.450 592.950 ;
        RECT 535.950 591.300 538.050 593.400 ;
        RECT 536.550 587.700 537.750 591.300 ;
        RECT 535.950 585.600 538.050 587.700 ;
        RECT 503.250 549.600 504.450 561.600 ;
        RECT 520.950 559.950 523.050 562.050 ;
        RECT 541.950 556.950 544.050 559.050 ;
        RECT 505.950 555.450 508.050 556.050 ;
        RECT 505.950 554.400 510.450 555.450 ;
        RECT 505.950 553.950 508.050 554.400 ;
        RECT 509.400 553.050 510.450 554.400 ;
        RECT 538.950 554.250 541.050 555.150 ;
        RECT 541.950 554.850 544.050 555.750 ;
        RECT 505.950 551.850 508.050 552.750 ;
        RECT 508.950 550.950 511.050 553.050 ;
        RECT 538.950 550.950 541.050 553.050 ;
        RECT 502.950 547.500 505.050 549.600 ;
        RECT 520.950 529.950 523.050 532.050 ;
        RECT 520.950 527.850 523.050 528.750 ;
        RECT 523.950 527.250 526.050 528.150 ;
        RECT 523.950 523.950 526.050 526.050 ;
        RECT 548.400 523.050 549.450 599.400 ;
        RECT 550.950 598.950 553.050 601.050 ;
        RECT 550.950 596.850 553.050 597.750 ;
        RECT 557.400 588.600 558.600 605.400 ;
        RECT 556.950 586.500 559.050 588.600 ;
        RECT 587.400 565.050 588.450 695.400 ;
        RECT 593.400 694.050 594.450 697.950 ;
        RECT 599.400 697.050 600.450 739.950 ;
        RECT 623.400 700.050 624.450 742.950 ;
        RECT 637.950 739.950 640.050 742.050 ;
        RECT 625.950 704.250 628.050 705.150 ;
        RECT 638.400 703.050 639.450 739.950 ;
        RECT 625.950 700.950 628.050 703.050 ;
        RECT 629.250 701.250 630.750 702.150 ;
        RECT 631.950 700.950 634.050 703.050 ;
        RECT 635.250 701.250 637.050 702.150 ;
        RECT 637.950 700.950 640.050 703.050 ;
        RECT 622.950 697.950 625.050 700.050 ;
        RECT 598.950 694.950 601.050 697.050 ;
        RECT 592.950 691.950 595.050 694.050 ;
        RECT 599.400 676.050 600.450 694.950 ;
        RECT 598.950 673.950 601.050 676.050 ;
        RECT 626.400 670.050 627.450 700.950 ;
        RECT 628.950 697.950 631.050 700.050 ;
        RECT 632.250 698.850 633.750 699.750 ;
        RECT 634.950 697.950 637.050 700.050 ;
        RECT 635.400 697.050 636.450 697.950 ;
        RECT 634.950 694.950 637.050 697.050 ;
        RECT 635.400 694.050 636.450 694.950 ;
        RECT 634.950 691.950 637.050 694.050 ;
        RECT 622.950 668.250 624.750 669.150 ;
        RECT 625.950 667.950 628.050 670.050 ;
        RECT 629.250 668.250 631.050 669.150 ;
        RECT 635.400 667.050 636.450 691.950 ;
        RECT 622.950 664.950 625.050 667.050 ;
        RECT 626.250 665.850 627.750 666.750 ;
        RECT 628.950 664.950 631.050 667.050 ;
        RECT 634.950 664.950 637.050 667.050 ;
        RECT 623.400 649.050 624.450 664.950 ;
        RECT 622.950 646.950 625.050 649.050 ;
        RECT 629.400 634.050 630.450 664.950 ;
        RECT 616.950 633.450 619.050 634.050 ;
        RECT 614.400 632.400 619.050 633.450 ;
        RECT 595.950 601.950 598.050 604.050 ;
        RECT 595.950 599.850 598.050 600.750 ;
        RECT 598.950 599.250 601.050 600.150 ;
        RECT 598.950 595.950 601.050 598.050 ;
        RECT 586.950 562.950 589.050 565.050 ;
        RECT 580.950 561.450 583.050 562.050 ;
        RECT 578.400 560.400 583.050 561.450 ;
        RECT 586.950 561.450 589.050 562.050 ;
        RECT 562.950 527.250 565.050 528.150 ;
        RECT 562.950 523.950 565.050 526.050 ;
        RECT 563.400 523.050 564.450 523.950 ;
        RECT 547.950 520.950 550.050 523.050 ;
        RECT 562.950 520.950 565.050 523.050 ;
        RECT 481.950 513.600 484.050 515.700 ;
        RECT 499.950 514.950 502.050 517.050 ;
        RECT 553.950 494.400 556.050 496.500 ;
        RECT 574.950 495.300 577.050 497.400 ;
        RECT 578.400 496.050 579.450 560.400 ;
        RECT 580.950 559.950 583.050 560.400 ;
        RECT 584.250 560.250 585.750 561.150 ;
        RECT 586.950 560.400 591.450 561.450 ;
        RECT 586.950 559.950 589.050 560.400 ;
        RECT 580.950 557.850 582.750 558.750 ;
        RECT 583.950 556.950 586.050 559.050 ;
        RECT 587.250 557.850 589.050 558.750 ;
        RECT 583.950 527.250 586.050 528.150 ;
        RECT 457.950 487.950 460.050 490.050 ;
        RECT 478.950 487.950 481.050 490.050 ;
        RECT 496.950 487.950 499.050 490.050 ;
        RECT 500.250 488.250 501.750 489.150 ;
        RECT 502.950 487.950 505.050 490.050 ;
        RECT 529.950 487.950 532.050 490.050 ;
        RECT 538.950 487.950 541.050 490.050 ;
        RECT 544.950 489.450 547.050 490.050 ;
        RECT 542.250 488.250 543.750 489.150 ;
        RECT 544.950 488.400 549.450 489.450 ;
        RECT 544.950 487.950 547.050 488.400 ;
        RECT 454.950 485.250 457.050 486.150 ;
        RECT 454.950 483.450 457.050 484.050 ;
        RECT 458.400 483.450 459.450 487.950 ;
        RECT 460.950 485.250 463.050 486.150 ;
        RECT 496.950 485.850 498.750 486.750 ;
        RECT 499.950 484.950 502.050 487.050 ;
        RECT 503.250 485.850 505.050 486.750 ;
        RECT 454.950 482.400 459.450 483.450 ;
        RECT 454.950 481.950 457.050 482.400 ;
        RECT 460.950 481.950 463.050 484.050 ;
        RECT 460.950 472.950 463.050 475.050 ;
        RECT 461.400 457.050 462.450 472.950 ;
        RECT 445.950 454.950 448.050 457.050 ;
        RECT 451.950 454.950 454.050 457.050 ;
        RECT 454.950 454.950 457.050 457.050 ;
        RECT 460.950 456.450 463.050 457.050 ;
        RECT 496.950 456.450 499.050 457.050 ;
        RECT 460.950 455.400 465.450 456.450 ;
        RECT 460.950 454.950 463.050 455.400 ;
        RECT 416.250 449.850 417.750 450.750 ;
        RECT 376.950 447.300 379.050 449.400 ;
        RECT 418.950 448.950 421.050 451.050 ;
        RECT 427.950 448.950 430.050 451.050 ;
        RECT 377.250 443.700 378.450 447.300 ;
        RECT 376.950 441.600 379.050 443.700 ;
        RECT 400.950 419.250 403.050 420.150 ;
        RECT 397.950 416.250 399.750 417.150 ;
        RECT 400.950 415.950 403.050 418.050 ;
        RECT 406.950 417.450 409.050 418.050 ;
        RECT 404.250 416.250 405.750 417.150 ;
        RECT 406.950 416.400 411.450 417.450 ;
        RECT 406.950 415.950 409.050 416.400 ;
        RECT 401.400 415.050 402.450 415.950 ;
        RECT 397.950 412.950 400.050 415.050 ;
        RECT 400.950 412.950 403.050 415.050 ;
        RECT 403.950 412.950 406.050 415.050 ;
        RECT 407.250 413.850 409.050 414.750 ;
        RECT 398.400 412.050 399.450 412.950 ;
        RECT 397.950 409.950 400.050 412.050 ;
        RECT 404.400 411.450 405.450 412.950 ;
        RECT 401.400 410.400 405.450 411.450 ;
        RECT 373.950 403.950 376.050 406.050 ;
        RECT 370.950 394.950 373.050 397.050 ;
        RECT 364.950 388.950 367.050 391.050 ;
        RECT 370.950 388.950 373.050 391.050 ;
        RECT 371.400 388.050 372.450 388.950 ;
        RECT 370.950 385.950 373.050 388.050 ;
        RECT 374.400 385.050 375.450 403.950 ;
        RECT 391.950 389.400 394.050 391.500 ;
        RECT 370.950 383.850 372.750 384.750 ;
        RECT 373.950 382.950 376.050 385.050 ;
        RECT 379.950 383.250 382.050 384.150 ;
        RECT 343.950 379.950 346.050 382.050 ;
        RECT 373.950 380.850 376.050 381.750 ;
        RECT 379.950 379.950 382.050 382.050 ;
        RECT 392.400 372.600 393.600 389.400 ;
        RECT 397.950 382.950 400.050 385.050 ;
        RECT 401.400 382.050 402.450 410.400 ;
        RECT 410.400 409.050 411.450 416.400 ;
        RECT 409.950 406.950 412.050 409.050 ;
        RECT 403.950 394.950 406.050 397.050 ;
        RECT 404.400 385.050 405.450 394.950 ;
        RECT 418.950 391.950 421.050 394.050 ;
        RECT 412.950 389.400 415.050 391.500 ;
        RECT 403.950 382.950 406.050 385.050 ;
        RECT 397.950 380.850 400.050 381.750 ;
        RECT 400.950 379.950 403.050 382.050 ;
        RECT 403.950 380.850 406.050 381.750 ;
        RECT 413.250 377.400 414.450 389.400 ;
        RECT 415.950 386.250 418.050 387.150 ;
        RECT 415.950 384.450 418.050 385.050 ;
        RECT 419.400 384.450 420.450 391.950 ;
        RECT 415.950 383.400 420.450 384.450 ;
        RECT 415.950 382.950 418.050 383.400 ;
        RECT 412.950 375.300 415.050 377.400 ;
        RECT 391.950 370.500 394.050 372.600 ;
        RECT 413.250 371.700 414.450 375.300 ;
        RECT 412.950 369.600 415.050 371.700 ;
        RECT 424.950 351.300 427.050 353.400 ;
        RECT 367.950 347.250 370.050 348.150 ;
        RECT 406.950 347.250 409.050 348.150 ;
        RECT 425.550 347.700 426.750 351.300 ;
        RECT 361.950 343.950 364.050 346.050 ;
        RECT 365.250 344.250 366.750 345.150 ;
        RECT 367.950 343.950 370.050 346.050 ;
        RECT 371.250 344.250 373.050 345.150 ;
        RECT 400.950 343.950 403.050 346.050 ;
        RECT 403.950 344.250 405.750 345.150 ;
        RECT 406.950 343.950 409.050 346.050 ;
        RECT 410.250 344.250 411.750 345.150 ;
        RECT 412.950 343.950 415.050 346.050 ;
        RECT 424.950 345.600 427.050 347.700 ;
        RECT 368.400 343.050 369.450 343.950 ;
        RECT 358.950 340.950 361.050 343.050 ;
        RECT 361.950 341.850 363.750 342.750 ;
        RECT 364.950 340.950 367.050 343.050 ;
        RECT 367.950 340.950 370.050 343.050 ;
        RECT 370.950 340.950 373.050 343.050 ;
        RECT 340.950 334.950 343.050 337.050 ;
        RECT 328.950 319.950 331.050 322.050 ;
        RECT 325.950 316.950 328.050 319.050 ;
        RECT 329.400 313.050 330.450 319.950 ;
        RECT 334.950 316.950 337.050 319.050 ;
        RECT 322.950 310.950 325.050 313.050 ;
        RECT 326.250 311.250 327.750 312.150 ;
        RECT 328.950 310.950 331.050 313.050 ;
        RECT 319.950 309.450 322.050 310.050 ;
        RECT 317.400 308.400 322.050 309.450 ;
        RECT 323.250 308.850 324.750 309.750 ;
        RECT 313.950 271.950 316.050 274.050 ;
        RECT 317.400 271.050 318.450 308.400 ;
        RECT 319.950 307.950 322.050 308.400 ;
        RECT 325.950 307.950 328.050 310.050 ;
        RECT 329.250 308.850 331.050 309.750 ;
        RECT 319.950 305.850 322.050 306.750 ;
        RECT 322.950 271.950 325.050 274.050 ;
        RECT 326.250 272.250 327.750 273.150 ;
        RECT 316.950 268.950 319.050 271.050 ;
        RECT 322.950 269.850 324.750 270.750 ;
        RECT 325.950 268.950 328.050 271.050 ;
        RECT 329.250 269.850 331.050 270.750 ;
        RECT 335.400 241.050 336.450 316.950 ;
        RECT 359.400 316.050 360.450 340.950 ;
        RECT 365.400 319.050 366.450 340.950 ;
        RECT 371.400 337.050 372.450 340.950 ;
        RECT 370.950 334.950 373.050 337.050 ;
        RECT 364.950 316.950 367.050 319.050 ;
        RECT 358.950 313.950 361.050 316.050 ;
        RECT 401.400 313.050 402.450 343.950 ;
        RECT 407.400 343.050 408.450 343.950 ;
        RECT 403.950 340.950 406.050 343.050 ;
        RECT 406.950 340.950 409.050 343.050 ;
        RECT 409.950 340.950 412.050 343.050 ;
        RECT 413.250 341.850 415.050 342.750 ;
        RECT 404.400 340.050 405.450 340.950 ;
        RECT 403.950 337.950 406.050 340.050 ;
        RECT 409.950 337.950 412.050 340.050 ;
        RECT 421.950 337.950 424.050 340.050 ;
        RECT 358.950 311.850 361.050 312.750 ;
        RECT 361.950 311.250 364.050 312.150 ;
        RECT 400.950 310.950 403.050 313.050 ;
        RECT 404.250 311.250 405.750 312.150 ;
        RECT 406.950 310.950 409.050 313.050 ;
        RECT 361.950 307.950 364.050 310.050 ;
        RECT 397.950 307.950 400.050 310.050 ;
        RECT 401.250 308.850 402.750 309.750 ;
        RECT 403.950 307.950 406.050 310.050 ;
        RECT 407.250 308.850 409.050 309.750 ;
        RECT 404.400 307.050 405.450 307.950 ;
        RECT 370.950 304.950 373.050 307.050 ;
        RECT 397.950 305.850 400.050 306.750 ;
        RECT 403.950 304.950 406.050 307.050 ;
        RECT 358.950 298.950 361.050 301.050 ;
        RECT 359.400 271.050 360.450 298.950 ;
        RECT 358.950 268.950 361.050 271.050 ;
        RECT 361.950 269.250 364.050 270.150 ;
        RECT 367.950 269.250 370.050 270.150 ;
        RECT 359.400 267.450 360.450 268.950 ;
        RECT 361.950 267.450 364.050 268.050 ;
        RECT 359.400 266.400 364.050 267.450 ;
        RECT 361.950 265.950 364.050 266.400 ;
        RECT 365.250 266.250 366.750 267.150 ;
        RECT 367.950 265.950 370.050 268.050 ;
        RECT 364.950 262.950 367.050 265.050 ;
        RECT 322.950 238.950 325.050 241.050 ;
        RECT 328.950 240.450 331.050 241.050 ;
        RECT 326.400 239.400 331.050 240.450 ;
        RECT 307.950 197.250 310.050 198.150 ;
        RECT 301.950 194.400 306.450 195.450 ;
        RECT 301.950 193.950 304.050 194.400 ;
        RECT 307.950 193.950 310.050 196.050 ;
        RECT 289.950 148.950 292.050 151.050 ;
        RECT 290.400 130.050 291.450 148.950 ;
        RECT 302.400 133.050 303.450 193.950 ;
        RECT 308.400 175.050 309.450 193.950 ;
        RECT 307.950 172.950 310.050 175.050 ;
        RECT 313.950 169.950 316.050 172.050 ;
        RECT 314.400 169.050 315.450 169.950 ;
        RECT 313.950 166.950 316.050 169.050 ;
        RECT 317.250 167.250 318.750 168.150 ;
        RECT 319.950 166.950 322.050 169.050 ;
        RECT 323.400 166.050 324.450 238.950 ;
        RECT 326.400 238.050 327.450 239.400 ;
        RECT 328.950 238.950 331.050 239.400 ;
        RECT 334.950 238.950 337.050 241.050 ;
        RECT 337.950 238.950 340.050 241.050 ;
        RECT 343.950 238.950 346.050 241.050 ;
        RECT 325.950 235.950 328.050 238.050 ;
        RECT 328.950 236.850 331.050 237.750 ;
        RECT 331.950 236.250 334.050 237.150 ;
        RECT 337.950 236.850 340.050 237.750 ;
        RECT 331.950 232.950 334.050 235.050 ;
        RECT 344.400 202.050 345.450 238.950 ;
        RECT 365.400 235.050 366.450 262.950 ;
        RECT 367.950 244.950 370.050 247.050 ;
        RECT 349.950 232.950 352.050 235.050 ;
        RECT 364.950 232.950 367.050 235.050 ;
        RECT 350.400 202.050 351.450 232.950 ;
        RECT 343.950 199.950 346.050 202.050 ;
        RECT 347.250 200.250 348.750 201.150 ;
        RECT 349.950 199.950 352.050 202.050 ;
        RECT 343.950 197.850 345.750 198.750 ;
        RECT 346.950 196.950 349.050 199.050 ;
        RECT 350.250 197.850 352.050 198.750 ;
        RECT 347.400 172.050 348.450 196.950 ;
        RECT 368.400 196.050 369.450 244.950 ;
        RECT 371.400 244.050 372.450 304.950 ;
        RECT 410.400 280.050 411.450 337.950 ;
        RECT 421.950 335.850 424.050 336.750 ;
        RECT 425.550 333.600 426.750 345.600 ;
        RECT 424.950 331.500 427.050 333.600 ;
        RECT 428.400 307.050 429.450 448.950 ;
        RECT 442.950 413.250 445.050 414.150 ;
        RECT 442.950 411.450 445.050 412.050 ;
        RECT 446.400 411.450 447.450 454.950 ;
        RECT 454.950 452.850 457.050 453.750 ;
        RECT 460.950 452.850 463.050 453.750 ;
        RECT 464.400 451.050 465.450 455.400 ;
        RECT 494.400 455.400 499.050 456.450 ;
        RECT 463.950 448.950 466.050 451.050 ;
        RECT 448.950 413.250 451.050 414.150 ;
        RECT 451.950 412.950 454.050 415.050 ;
        RECT 442.950 410.400 447.450 411.450 ;
        RECT 448.950 411.450 451.050 412.050 ;
        RECT 452.400 411.450 453.450 412.950 ;
        RECT 464.400 412.050 465.450 448.950 ;
        RECT 484.950 424.950 487.050 427.050 ;
        RECT 485.400 414.450 486.450 424.950 ;
        RECT 494.400 421.050 495.450 455.400 ;
        RECT 496.950 454.950 499.050 455.400 ;
        RECT 496.950 452.850 499.050 453.750 ;
        RECT 500.400 427.050 501.450 484.950 ;
        RECT 502.950 481.950 505.050 484.050 ;
        RECT 503.400 457.050 504.450 481.950 ;
        RECT 502.950 454.950 505.050 457.050 ;
        RECT 502.950 452.850 505.050 453.750 ;
        RECT 499.950 424.950 502.050 427.050 ;
        RECT 505.950 422.400 508.050 424.500 ;
        RECT 526.950 423.300 529.050 425.400 ;
        RECT 493.950 418.950 496.050 421.050 ;
        RECT 499.950 418.950 502.050 421.050 ;
        RECT 487.950 416.250 490.050 417.150 ;
        RECT 493.950 415.950 496.050 418.050 ;
        RECT 494.400 415.050 495.450 415.950 ;
        RECT 487.950 414.450 490.050 415.050 ;
        RECT 485.400 413.400 490.050 414.450 ;
        RECT 487.950 412.950 490.050 413.400 ;
        RECT 491.250 413.250 492.750 414.150 ;
        RECT 493.950 412.950 496.050 415.050 ;
        RECT 497.250 413.250 499.050 414.150 ;
        RECT 448.950 410.400 453.450 411.450 ;
        RECT 442.950 409.950 445.050 410.400 ;
        RECT 448.950 409.950 451.050 410.400 ;
        RECT 463.950 409.950 466.050 412.050 ;
        RECT 490.950 409.950 493.050 412.050 ;
        RECT 494.250 410.850 495.750 411.750 ;
        RECT 496.950 411.450 499.050 412.050 ;
        RECT 500.400 411.450 501.450 418.950 ;
        RECT 496.950 410.400 501.450 411.450 ;
        RECT 496.950 409.950 499.050 410.400 ;
        RECT 436.950 394.950 439.050 397.050 ;
        RECT 433.950 341.250 436.050 342.150 ;
        RECT 433.950 339.450 436.050 340.050 ;
        RECT 437.400 339.450 438.450 394.950 ;
        RECT 439.950 341.250 442.050 342.150 ;
        RECT 433.950 338.400 438.450 339.450 ;
        RECT 433.950 337.950 436.050 338.400 ;
        RECT 439.950 337.950 442.050 340.050 ;
        RECT 439.950 334.950 442.050 337.050 ;
        RECT 440.400 316.050 441.450 334.950 ;
        RECT 443.400 316.050 444.450 409.950 ;
        RECT 449.400 382.050 450.450 409.950 ;
        RECT 506.400 405.600 507.600 422.400 ;
        RECT 527.250 419.700 528.450 423.300 ;
        RECT 520.950 415.950 523.050 418.050 ;
        RECT 526.950 417.600 529.050 419.700 ;
        RECT 511.950 413.250 514.050 414.150 ;
        RECT 517.950 413.250 520.050 414.150 ;
        RECT 511.950 409.950 514.050 412.050 ;
        RECT 517.950 409.950 520.050 412.050 ;
        RECT 505.950 403.500 508.050 405.600 ;
        RECT 518.400 397.050 519.450 409.950 ;
        RECT 514.950 394.950 517.050 397.050 ;
        RECT 517.950 394.950 520.050 397.050 ;
        RECT 502.950 391.950 505.050 394.050 ;
        RECT 503.400 388.050 504.450 391.950 ;
        RECT 502.950 385.950 505.050 388.050 ;
        RECT 457.950 382.950 460.050 385.050 ;
        RECT 463.950 384.450 466.050 385.050 ;
        RECT 461.250 383.250 462.750 384.150 ;
        RECT 463.950 383.400 468.450 384.450 ;
        RECT 463.950 382.950 466.050 383.400 ;
        RECT 467.400 382.050 468.450 383.400 ;
        RECT 499.950 383.250 502.050 384.150 ;
        RECT 502.950 383.850 505.050 384.750 ;
        RECT 448.950 379.950 451.050 382.050 ;
        RECT 454.950 381.450 457.050 382.050 ;
        RECT 452.400 380.400 457.050 381.450 ;
        RECT 458.250 380.850 459.750 381.750 ;
        RECT 452.400 379.050 453.450 380.400 ;
        RECT 454.950 379.950 457.050 380.400 ;
        RECT 460.950 379.950 463.050 382.050 ;
        RECT 464.250 380.850 466.050 381.750 ;
        RECT 466.950 379.950 469.050 382.050 ;
        RECT 499.950 379.950 502.050 382.050 ;
        RECT 451.950 376.950 454.050 379.050 ;
        RECT 454.950 377.850 457.050 378.750 ;
        RECT 445.950 350.400 448.050 352.500 ;
        RECT 446.400 333.600 447.600 350.400 ;
        RECT 461.400 343.050 462.450 379.950 ;
        RECT 466.950 376.950 469.050 379.050 ;
        RECT 460.950 340.950 463.050 343.050 ;
        RECT 445.950 331.500 448.050 333.600 ;
        RECT 439.950 313.950 442.050 316.050 ;
        RECT 442.950 313.950 445.050 316.050 ;
        RECT 439.950 311.850 442.050 312.750 ;
        RECT 442.950 311.250 445.050 312.150 ;
        RECT 442.950 307.950 445.050 310.050 ;
        RECT 427.950 304.950 430.050 307.050 ;
        RECT 439.950 304.950 442.050 307.050 ;
        RECT 409.950 277.950 412.050 280.050 ;
        RECT 400.950 268.950 403.050 271.050 ;
        RECT 406.950 268.950 409.050 271.050 ;
        RECT 401.400 264.450 402.450 268.950 ;
        RECT 403.950 266.250 406.050 267.150 ;
        RECT 406.950 266.850 409.050 267.750 ;
        RECT 403.950 264.450 406.050 265.050 ;
        RECT 401.400 263.400 406.050 264.450 ;
        RECT 403.950 262.950 406.050 263.400 ;
        RECT 370.950 241.950 373.050 244.050 ;
        RECT 371.400 241.050 372.450 241.950 ;
        RECT 370.950 238.950 373.050 241.050 ;
        RECT 374.250 239.250 375.750 240.150 ;
        RECT 376.950 238.950 379.050 241.050 ;
        RECT 379.950 238.950 382.050 241.050 ;
        RECT 380.400 238.050 381.450 238.950 ;
        RECT 370.950 236.850 372.750 237.750 ;
        RECT 373.950 235.950 376.050 238.050 ;
        RECT 377.250 236.850 378.750 237.750 ;
        RECT 379.950 235.950 382.050 238.050 ;
        RECT 374.400 202.050 375.450 235.950 ;
        RECT 379.950 233.850 382.050 234.750 ;
        RECT 373.950 199.950 376.050 202.050 ;
        RECT 367.950 193.950 370.050 196.050 ;
        RECT 374.400 193.050 375.450 199.950 ;
        RECT 382.950 197.250 385.050 198.150 ;
        RECT 388.950 197.250 391.050 198.150 ;
        RECT 382.950 193.950 385.050 196.050 ;
        RECT 388.950 193.950 391.050 196.050 ;
        RECT 373.950 190.950 376.050 193.050 ;
        RECT 389.400 190.050 390.450 193.950 ;
        RECT 388.950 187.950 391.050 190.050 ;
        RECT 410.400 175.050 411.450 277.950 ;
        RECT 421.950 271.950 424.050 274.050 ;
        RECT 412.950 268.950 415.050 271.050 ;
        RECT 413.400 241.050 414.450 268.950 ;
        RECT 422.400 241.050 423.450 271.950 ;
        RECT 427.950 241.950 430.050 244.050 ;
        RECT 428.400 241.050 429.450 241.950 ;
        RECT 412.950 238.950 415.050 241.050 ;
        RECT 421.950 238.950 424.050 241.050 ;
        RECT 425.250 239.250 426.750 240.150 ;
        RECT 427.950 238.950 430.050 241.050 ;
        RECT 413.400 235.050 414.450 238.950 ;
        RECT 418.950 237.450 421.050 238.050 ;
        RECT 416.400 236.400 421.050 237.450 ;
        RECT 422.250 236.850 423.750 237.750 ;
        RECT 412.950 232.950 415.050 235.050 ;
        RECT 416.400 232.050 417.450 236.400 ;
        RECT 418.950 235.950 421.050 236.400 ;
        RECT 424.950 235.950 427.050 238.050 ;
        RECT 428.250 236.850 430.050 237.750 ;
        RECT 425.400 235.050 426.450 235.950 ;
        RECT 418.950 233.850 421.050 234.750 ;
        RECT 424.950 232.950 427.050 235.050 ;
        RECT 415.950 229.950 418.050 232.050 ;
        RECT 433.950 199.950 436.050 202.050 ;
        RECT 424.950 197.250 427.050 198.150 ;
        RECT 430.950 197.250 433.050 198.150 ;
        RECT 424.950 193.950 427.050 196.050 ;
        RECT 430.950 195.450 433.050 196.050 ;
        RECT 434.400 195.450 435.450 199.950 ;
        RECT 428.250 194.250 429.750 195.150 ;
        RECT 430.950 194.400 435.450 195.450 ;
        RECT 430.950 193.950 433.050 194.400 ;
        RECT 427.950 190.950 430.050 193.050 ;
        RECT 418.950 187.950 421.050 190.050 ;
        RECT 400.950 172.950 403.050 175.050 ;
        RECT 409.950 172.950 412.050 175.050 ;
        RECT 346.950 169.950 349.050 172.050 ;
        RECT 347.400 169.050 348.450 169.950 ;
        RECT 346.950 166.950 349.050 169.050 ;
        RECT 401.400 166.050 402.450 172.950 ;
        RECT 313.950 164.850 315.750 165.750 ;
        RECT 316.950 163.950 319.050 166.050 ;
        RECT 320.250 164.850 321.750 165.750 ;
        RECT 322.950 163.950 325.050 166.050 ;
        RECT 337.950 163.950 340.050 166.050 ;
        RECT 361.950 164.250 363.750 165.150 ;
        RECT 364.950 163.950 367.050 166.050 ;
        RECT 368.250 164.250 370.050 165.150 ;
        RECT 400.950 163.950 403.050 166.050 ;
        RECT 403.950 163.950 406.050 166.050 ;
        RECT 406.950 163.950 409.050 166.050 ;
        RECT 410.250 164.250 412.050 165.150 ;
        RECT 295.950 131.250 298.050 132.150 ;
        RECT 301.950 130.950 304.050 133.050 ;
        RECT 289.950 127.950 292.050 130.050 ;
        RECT 292.950 128.250 294.750 129.150 ;
        RECT 295.950 127.950 298.050 130.050 ;
        RECT 301.950 129.450 304.050 130.050 ;
        RECT 299.250 128.250 300.750 129.150 ;
        RECT 301.950 128.400 306.450 129.450 ;
        RECT 301.950 127.950 304.050 128.400 ;
        RECT 292.950 124.950 295.050 127.050 ;
        RECT 298.950 124.950 301.050 127.050 ;
        RECT 302.250 125.850 304.050 126.750 ;
        RECT 293.400 121.050 294.450 124.950 ;
        RECT 292.950 118.950 295.050 121.050 ;
        RECT 299.400 115.050 300.450 124.950 ;
        RECT 305.400 124.050 306.450 128.400 ;
        RECT 304.950 121.950 307.050 124.050 ;
        RECT 298.950 112.950 301.050 115.050 ;
        RECT 280.950 96.450 283.050 97.050 ;
        RECT 280.950 95.400 285.450 96.450 ;
        RECT 280.950 94.950 283.050 95.400 ;
        RECT 280.950 92.850 283.050 93.750 ;
        RECT 284.400 91.050 285.450 95.400 ;
        RECT 317.400 94.050 318.450 163.950 ;
        RECT 322.950 161.850 325.050 162.750 ;
        RECT 338.400 133.050 339.450 163.950 ;
        RECT 404.400 163.050 405.450 163.950 ;
        RECT 361.950 160.950 364.050 163.050 ;
        RECT 365.250 161.850 366.750 162.750 ;
        RECT 367.950 160.950 370.050 163.050 ;
        RECT 400.950 161.850 402.750 162.750 ;
        RECT 403.950 160.950 406.050 163.050 ;
        RECT 407.250 161.850 408.750 162.750 ;
        RECT 409.950 162.450 412.050 163.050 ;
        RECT 409.950 161.400 414.450 162.450 ;
        RECT 409.950 160.950 412.050 161.400 ;
        RECT 368.400 154.050 369.450 160.950 ;
        RECT 403.950 158.850 406.050 159.750 ;
        RECT 409.950 157.950 412.050 160.050 ;
        RECT 367.950 151.950 370.050 154.050 ;
        RECT 376.950 151.950 379.050 154.050 ;
        RECT 337.950 130.950 340.050 133.050 ;
        RECT 338.400 130.050 339.450 130.950 ;
        RECT 328.950 127.950 331.050 130.050 ;
        RECT 337.950 127.950 340.050 130.050 ;
        RECT 341.250 128.250 342.750 129.150 ;
        RECT 343.950 127.950 346.050 130.050 ;
        RECT 322.950 97.950 325.050 100.050 ;
        RECT 313.950 92.250 315.750 93.150 ;
        RECT 316.950 91.950 319.050 94.050 ;
        RECT 320.250 92.250 322.050 93.150 ;
        RECT 274.950 89.400 279.450 90.450 ;
        RECT 274.950 88.950 277.050 89.400 ;
        RECT 283.950 88.950 286.050 91.050 ;
        RECT 313.950 88.950 316.050 91.050 ;
        RECT 317.250 89.850 318.750 90.750 ;
        RECT 319.950 90.450 322.050 91.050 ;
        RECT 323.400 90.450 324.450 97.950 ;
        RECT 319.950 89.400 324.450 90.450 ;
        RECT 319.950 88.950 322.050 89.400 ;
        RECT 280.950 53.250 283.050 54.150 ;
        RECT 286.950 53.250 289.050 54.150 ;
        RECT 307.950 52.950 310.050 55.050 ;
        RECT 280.950 49.950 283.050 52.050 ;
        RECT 284.250 50.250 285.750 51.150 ;
        RECT 286.950 49.950 289.050 52.050 ;
        RECT 205.950 22.950 208.050 25.050 ;
        RECT 211.950 22.950 214.050 25.050 ;
        RECT 205.950 20.850 208.050 21.750 ;
        RECT 211.950 20.850 214.050 21.750 ;
        RECT 181.950 15.300 184.050 17.400 ;
        RECT 196.950 15.300 199.050 17.400 ;
        RECT 64.950 9.600 67.050 11.700 ;
        RECT 160.950 10.500 163.050 12.600 ;
        RECT 182.250 11.700 183.450 15.300 ;
        RECT 197.550 11.700 198.750 15.300 ;
        RECT 218.400 12.600 219.600 29.400 ;
        RECT 259.950 28.950 262.050 31.050 ;
        RECT 281.400 25.050 282.450 49.950 ;
        RECT 287.400 49.050 288.450 49.950 ;
        RECT 283.950 46.950 286.050 49.050 ;
        RECT 286.950 46.950 289.050 49.050 ;
        RECT 280.950 22.950 283.050 25.050 ;
        RECT 259.950 20.250 261.750 21.150 ;
        RECT 262.950 19.950 265.050 22.050 ;
        RECT 266.250 20.250 268.050 21.150 ;
        RECT 284.400 19.050 285.450 46.950 ;
        RECT 308.400 25.050 309.450 52.950 ;
        RECT 314.400 49.050 315.450 88.950 ;
        RECT 322.950 52.950 325.050 55.050 ;
        RECT 322.950 50.850 325.050 51.750 ;
        RECT 325.950 50.250 328.050 51.150 ;
        RECT 313.950 46.950 316.050 49.050 ;
        RECT 325.950 48.450 328.050 49.050 ;
        RECT 329.400 48.450 330.450 127.950 ;
        RECT 337.950 125.850 339.750 126.750 ;
        RECT 340.950 124.950 343.050 127.050 ;
        RECT 344.250 125.850 346.050 126.750 ;
        RECT 358.950 124.950 361.050 127.050 ;
        RECT 341.400 97.050 342.450 124.950 ;
        RECT 340.950 94.950 343.050 97.050 ;
        RECT 359.400 94.050 360.450 124.950 ;
        RECT 355.950 92.250 357.750 93.150 ;
        RECT 358.950 91.950 361.050 94.050 ;
        RECT 362.250 92.250 364.050 93.150 ;
        RECT 355.950 88.950 358.050 91.050 ;
        RECT 359.250 89.850 360.750 90.750 ;
        RECT 361.950 88.950 364.050 91.050 ;
        RECT 356.400 55.050 357.450 88.950 ;
        RECT 373.950 55.950 376.050 58.050 ;
        RECT 355.950 52.950 358.050 55.050 ;
        RECT 361.950 53.250 364.050 54.150 ;
        RECT 367.950 53.250 370.050 54.150 ;
        RECT 370.950 52.950 373.050 55.050 ;
        RECT 361.950 49.950 364.050 52.050 ;
        RECT 367.950 51.450 370.050 52.050 ;
        RECT 371.400 51.450 372.450 52.950 ;
        RECT 365.250 50.250 366.750 51.150 ;
        RECT 367.950 50.400 372.450 51.450 ;
        RECT 367.950 49.950 370.050 50.400 ;
        RECT 325.950 47.400 330.450 48.450 ;
        RECT 325.950 46.950 328.050 47.400 ;
        RECT 364.950 46.950 367.050 49.050 ;
        RECT 316.950 29.400 319.050 31.500 ;
        RECT 301.950 22.950 304.050 25.050 ;
        RECT 305.250 23.250 306.750 24.150 ;
        RECT 307.950 22.950 310.050 25.050 ;
        RECT 298.950 19.950 301.050 22.050 ;
        RECT 302.250 20.850 303.750 21.750 ;
        RECT 304.950 19.950 307.050 22.050 ;
        RECT 308.250 20.850 310.050 21.750 ;
        RECT 305.400 19.050 306.450 19.950 ;
        RECT 259.950 16.950 262.050 19.050 ;
        RECT 263.250 17.850 264.750 18.750 ;
        RECT 283.950 16.950 286.050 19.050 ;
        RECT 298.950 17.850 301.050 18.750 ;
        RECT 304.950 16.950 307.050 19.050 ;
        RECT 317.400 12.600 318.600 29.400 ;
        RECT 326.400 25.050 327.450 46.950 ;
        RECT 328.950 43.950 331.050 46.050 ;
        RECT 329.400 25.050 330.450 43.950 ;
        RECT 337.950 29.400 340.050 31.500 ;
        RECT 322.950 22.950 325.050 25.050 ;
        RECT 325.950 22.950 328.050 25.050 ;
        RECT 328.950 22.950 331.050 25.050 ;
        RECT 322.950 20.850 325.050 21.750 ;
        RECT 328.950 20.850 331.050 21.750 ;
        RECT 338.250 17.400 339.450 29.400 ;
        RECT 340.950 26.250 343.050 27.150 ;
        RECT 340.950 22.950 343.050 25.050 ;
        RECT 374.400 19.050 375.450 55.950 ;
        RECT 377.400 40.050 378.450 151.950 ;
        RECT 379.950 130.950 382.050 133.050 ;
        RECT 380.400 130.050 381.450 130.950 ;
        RECT 379.950 127.950 382.050 130.050 ;
        RECT 385.950 129.450 388.050 130.050 ;
        RECT 383.250 128.250 384.750 129.150 ;
        RECT 385.950 128.400 390.450 129.450 ;
        RECT 385.950 127.950 388.050 128.400 ;
        RECT 379.950 125.850 381.750 126.750 ;
        RECT 382.950 124.950 385.050 127.050 ;
        RECT 386.250 125.850 388.050 126.750 ;
        RECT 383.400 94.050 384.450 124.950 ;
        RECT 389.400 124.050 390.450 128.400 ;
        RECT 388.950 121.950 391.050 124.050 ;
        RECT 400.950 94.950 403.050 97.050 ;
        RECT 382.950 91.950 385.050 94.050 ;
        RECT 397.950 93.450 400.050 94.050 ;
        RECT 395.400 92.400 400.050 93.450 ;
        RECT 383.400 91.050 384.450 91.950 ;
        RECT 382.950 88.950 385.050 91.050 ;
        RECT 395.400 85.050 396.450 92.400 ;
        RECT 397.950 91.950 400.050 92.400 ;
        RECT 401.400 91.050 402.450 94.950 ;
        RECT 403.950 91.950 406.050 94.050 ;
        RECT 407.250 92.250 409.050 93.150 ;
        RECT 397.950 89.850 399.750 90.750 ;
        RECT 400.950 88.950 403.050 91.050 ;
        RECT 404.250 89.850 405.750 90.750 ;
        RECT 406.950 90.450 409.050 91.050 ;
        RECT 410.400 90.450 411.450 157.950 ;
        RECT 413.400 157.050 414.450 161.400 ;
        RECT 412.950 154.950 415.050 157.050 ;
        RECT 419.400 126.450 420.450 187.950 ;
        RECT 436.950 163.950 439.050 166.050 ;
        RECT 437.400 151.050 438.450 163.950 ;
        RECT 436.950 148.950 439.050 151.050 ;
        RECT 424.950 131.250 427.050 132.150 ;
        RECT 421.950 128.250 423.750 129.150 ;
        RECT 424.950 127.950 427.050 130.050 ;
        RECT 428.250 128.250 429.750 129.150 ;
        RECT 430.950 127.950 433.050 130.050 ;
        RECT 421.950 126.450 424.050 127.050 ;
        RECT 419.400 125.400 424.050 126.450 ;
        RECT 421.950 124.950 424.050 125.400 ;
        RECT 427.950 124.950 430.050 127.050 ;
        RECT 431.250 125.850 433.050 126.750 ;
        RECT 428.400 124.050 429.450 124.950 ;
        RECT 427.950 121.950 430.050 124.050 ;
        RECT 436.950 97.950 439.050 100.050 ;
        RECT 406.950 89.400 411.450 90.450 ;
        RECT 406.950 88.950 409.050 89.400 ;
        RECT 400.950 86.850 403.050 87.750 ;
        RECT 394.950 82.950 397.050 85.050 ;
        RECT 400.950 82.950 403.050 85.050 ;
        RECT 401.400 55.050 402.450 82.950 ;
        RECT 412.950 62.400 415.050 64.500 ;
        RECT 400.950 52.950 403.050 55.050 ;
        RECT 400.950 50.850 403.050 51.750 ;
        RECT 403.950 50.250 406.050 51.150 ;
        RECT 403.950 46.950 406.050 49.050 ;
        RECT 404.400 40.050 405.450 46.950 ;
        RECT 413.400 45.600 414.600 62.400 ;
        RECT 427.950 61.950 430.050 64.050 ;
        RECT 433.950 63.300 436.050 65.400 ;
        RECT 418.950 53.250 421.050 54.150 ;
        RECT 424.950 53.250 427.050 54.150 ;
        RECT 418.950 51.450 421.050 52.050 ;
        RECT 418.950 50.400 423.450 51.450 ;
        RECT 418.950 49.950 421.050 50.400 ;
        RECT 412.950 43.500 415.050 45.600 ;
        RECT 376.950 37.950 379.050 40.050 ;
        RECT 403.950 37.950 406.050 40.050 ;
        RECT 376.950 28.950 379.050 31.050 ;
        RECT 337.950 15.300 340.050 17.400 ;
        RECT 373.950 16.950 376.050 19.050 ;
        RECT 377.400 18.450 378.450 28.950 ;
        RECT 422.400 25.050 423.450 50.400 ;
        RECT 424.950 49.950 427.050 52.050 ;
        RECT 425.400 46.050 426.450 49.950 ;
        RECT 424.950 43.950 427.050 46.050 ;
        RECT 428.400 25.050 429.450 61.950 ;
        RECT 434.250 59.700 435.450 63.300 ;
        RECT 433.950 57.600 436.050 59.700 ;
        RECT 434.250 45.600 435.450 57.600 ;
        RECT 437.400 55.050 438.450 97.950 ;
        RECT 440.400 58.050 441.450 304.950 ;
        RECT 445.950 271.950 448.050 274.050 ;
        RECT 451.950 273.450 454.050 274.050 ;
        RECT 449.250 272.250 450.750 273.150 ;
        RECT 451.950 272.400 456.450 273.450 ;
        RECT 451.950 271.950 454.050 272.400 ;
        RECT 445.950 269.850 447.750 270.750 ;
        RECT 448.950 268.950 451.050 271.050 ;
        RECT 452.250 269.850 454.050 270.750 ;
        RECT 455.400 268.050 456.450 272.400 ;
        RECT 454.950 265.950 457.050 268.050 ;
        RECT 445.950 241.950 448.050 244.050 ;
        RECT 460.950 243.450 463.050 244.050 ;
        RECT 458.400 242.400 463.050 243.450 ;
        RECT 446.400 172.050 447.450 241.950 ;
        RECT 458.400 232.050 459.450 242.400 ;
        RECT 460.950 241.950 463.050 242.400 ;
        RECT 460.950 239.850 462.750 240.750 ;
        RECT 463.950 238.950 466.050 241.050 ;
        RECT 463.950 236.850 466.050 237.750 ;
        RECT 467.400 234.450 468.450 376.950 ;
        RECT 505.950 350.400 508.050 352.500 ;
        RECT 484.950 343.950 487.050 346.050 ;
        RECT 487.950 344.250 490.050 345.150 ;
        RECT 485.400 342.450 486.450 343.950 ;
        RECT 487.950 342.450 490.050 343.050 ;
        RECT 485.400 341.400 490.050 342.450 ;
        RECT 487.950 340.950 490.050 341.400 ;
        RECT 491.250 341.250 492.750 342.150 ;
        RECT 493.950 340.950 496.050 343.050 ;
        RECT 497.250 341.250 499.050 342.150 ;
        RECT 484.950 337.950 487.050 340.050 ;
        RECT 490.950 337.950 493.050 340.050 ;
        RECT 494.250 338.850 495.750 339.750 ;
        RECT 496.950 337.950 499.050 340.050 ;
        RECT 478.950 319.950 481.050 322.050 ;
        RECT 479.400 313.050 480.450 319.950 ;
        RECT 485.400 313.050 486.450 337.950 ;
        RECT 497.400 337.050 498.450 337.950 ;
        RECT 496.950 334.950 499.050 337.050 ;
        RECT 506.400 333.600 507.600 350.400 ;
        RECT 511.950 341.250 514.050 342.150 ;
        RECT 511.950 337.950 514.050 340.050 ;
        RECT 515.400 339.450 516.450 394.950 ;
        RECT 517.950 341.250 520.050 342.150 ;
        RECT 517.950 339.450 520.050 340.050 ;
        RECT 515.400 338.400 520.050 339.450 ;
        RECT 517.950 337.950 520.050 338.400 ;
        RECT 521.400 336.450 522.450 415.950 ;
        RECT 527.250 405.600 528.450 417.600 ;
        RECT 530.400 412.050 531.450 487.950 ;
        RECT 538.950 485.850 540.750 486.750 ;
        RECT 541.950 484.950 544.050 487.050 ;
        RECT 545.250 485.850 547.050 486.750 ;
        RECT 548.400 481.050 549.450 488.400 ;
        RECT 547.950 478.950 550.050 481.050 ;
        RECT 554.400 477.600 555.600 494.400 ;
        RECT 575.250 491.700 576.450 495.300 ;
        RECT 577.950 493.950 580.050 496.050 ;
        RECT 574.950 489.600 577.050 491.700 ;
        RECT 559.950 485.250 562.050 486.150 ;
        RECT 565.950 485.250 568.050 486.150 ;
        RECT 559.950 481.950 562.050 484.050 ;
        RECT 565.950 481.950 568.050 484.050 ;
        RECT 553.950 475.500 556.050 477.600 ;
        RECT 560.400 472.050 561.450 481.950 ;
        RECT 559.950 469.950 562.050 472.050 ;
        RECT 544.950 457.950 547.050 460.050 ;
        RECT 545.400 457.050 546.450 457.950 ;
        RECT 544.950 454.950 547.050 457.050 ;
        RECT 535.950 452.250 537.750 453.150 ;
        RECT 538.950 451.950 541.050 454.050 ;
        RECT 542.250 452.250 544.050 453.150 ;
        RECT 535.950 448.950 538.050 451.050 ;
        RECT 539.250 449.850 540.750 450.750 ;
        RECT 541.950 448.950 544.050 451.050 ;
        RECT 536.400 448.050 537.450 448.950 ;
        RECT 535.950 445.950 538.050 448.050 ;
        RECT 529.950 409.950 532.050 412.050 ;
        RECT 529.950 407.850 532.050 408.750 ;
        RECT 526.950 403.500 529.050 405.600 ;
        RECT 545.400 391.050 546.450 454.950 ;
        RECT 566.400 397.050 567.450 481.950 ;
        RECT 575.250 477.600 576.450 489.600 ;
        RECT 577.950 483.450 580.050 484.050 ;
        RECT 577.950 482.400 582.450 483.450 ;
        RECT 577.950 481.950 580.050 482.400 ;
        RECT 577.950 479.850 580.050 480.750 ;
        RECT 581.400 478.050 582.450 482.400 ;
        RECT 590.400 481.050 591.450 560.400 ;
        RECT 614.400 493.050 615.450 632.400 ;
        RECT 616.950 631.950 619.050 632.400 ;
        RECT 620.250 632.250 621.750 633.150 ;
        RECT 622.950 631.950 625.050 634.050 ;
        RECT 628.950 631.950 631.050 634.050 ;
        RECT 616.950 629.850 618.750 630.750 ;
        RECT 619.950 628.950 622.050 631.050 ;
        RECT 623.250 629.850 625.050 630.750 ;
        RECT 634.950 622.950 637.050 625.050 ;
        RECT 635.400 601.050 636.450 622.950 ;
        RECT 641.400 601.050 642.450 745.950 ;
        RECT 683.400 745.050 684.450 745.950 ;
        RECT 682.950 742.950 685.050 745.050 ;
        RECT 715.950 742.950 718.050 745.050 ;
        RECT 676.950 740.850 679.050 741.750 ;
        RECT 682.950 740.850 685.050 741.750 ;
        RECT 715.950 740.850 718.050 741.750 ;
        RECT 721.950 740.850 724.050 741.750 ;
        RECT 739.950 703.950 742.050 706.050 ;
        RECT 748.950 703.950 751.050 706.050 ;
        RECT 754.950 705.450 757.050 706.050 ;
        RECT 752.250 704.250 753.750 705.150 ;
        RECT 754.950 704.400 759.450 705.450 ;
        RECT 754.950 703.950 757.050 704.400 ;
        RECT 667.950 701.250 670.050 702.150 ;
        RECT 673.950 701.250 676.050 702.150 ;
        RECT 709.950 701.250 712.050 702.150 ;
        RECT 715.950 701.250 718.050 702.150 ;
        RECT 667.950 697.950 670.050 700.050 ;
        RECT 709.950 697.950 712.050 700.050 ;
        RECT 668.400 673.050 669.450 697.950 ;
        RECT 673.950 694.950 676.050 697.050 ;
        RECT 674.400 673.050 675.450 694.950 ;
        RECT 700.950 673.950 703.050 676.050 ;
        RECT 655.950 670.950 658.050 673.050 ;
        RECT 664.950 670.950 667.050 673.050 ;
        RECT 667.950 670.950 670.050 673.050 ;
        RECT 671.250 671.250 672.750 672.150 ;
        RECT 673.950 670.950 676.050 673.050 ;
        RECT 634.950 598.950 637.050 601.050 ;
        RECT 638.250 599.250 639.750 600.150 ;
        RECT 640.950 598.950 643.050 601.050 ;
        RECT 634.950 596.850 636.750 597.750 ;
        RECT 637.950 595.950 640.050 598.050 ;
        RECT 641.250 596.850 642.750 597.750 ;
        RECT 643.950 597.450 646.050 598.050 ;
        RECT 643.950 596.400 648.450 597.450 ;
        RECT 643.950 595.950 646.050 596.400 ;
        RECT 643.950 593.850 646.050 594.750 ;
        RECT 628.950 560.250 631.050 561.150 ;
        RECT 647.400 559.050 648.450 596.400 ;
        RECT 619.950 557.250 621.750 558.150 ;
        RECT 622.950 556.950 625.050 559.050 ;
        RECT 628.950 558.450 631.050 559.050 ;
        RECT 626.250 557.250 627.750 558.150 ;
        RECT 628.950 557.400 633.450 558.450 ;
        RECT 628.950 556.950 631.050 557.400 ;
        RECT 619.950 553.950 622.050 556.050 ;
        RECT 623.250 554.850 624.750 555.750 ;
        RECT 625.950 553.950 628.050 556.050 ;
        RECT 620.400 523.050 621.450 553.950 ;
        RECT 625.950 550.950 628.050 553.050 ;
        RECT 626.400 526.050 627.450 550.950 ;
        RECT 622.950 524.250 624.750 525.150 ;
        RECT 625.950 523.950 628.050 526.050 ;
        RECT 629.250 524.250 631.050 525.150 ;
        RECT 619.950 520.950 622.050 523.050 ;
        RECT 622.950 520.950 625.050 523.050 ;
        RECT 626.250 521.850 627.750 522.750 ;
        RECT 628.950 520.950 631.050 523.050 ;
        RECT 613.950 490.950 616.050 493.050 ;
        RECT 619.950 488.250 622.050 489.150 ;
        RECT 607.950 484.950 610.050 487.050 ;
        RECT 610.950 485.250 612.750 486.150 ;
        RECT 613.950 484.950 616.050 487.050 ;
        RECT 617.250 485.250 618.750 486.150 ;
        RECT 619.950 484.950 622.050 487.050 ;
        RECT 589.950 478.950 592.050 481.050 ;
        RECT 574.950 475.500 577.050 477.600 ;
        RECT 580.950 475.950 583.050 478.050 ;
        RECT 583.950 469.950 586.050 472.050 ;
        RECT 584.400 457.050 585.450 469.950 ;
        RECT 574.950 454.950 577.050 457.050 ;
        RECT 583.950 454.950 586.050 457.050 ;
        RECT 587.250 455.250 588.750 456.150 ;
        RECT 589.950 454.950 592.050 457.050 ;
        RECT 568.950 416.250 571.050 417.150 ;
        RECT 575.400 415.050 576.450 454.950 ;
        RECT 580.950 451.950 583.050 454.050 ;
        RECT 584.250 452.850 585.750 453.750 ;
        RECT 586.950 451.950 589.050 454.050 ;
        RECT 590.250 452.850 592.050 453.750 ;
        RECT 580.950 449.850 583.050 450.750 ;
        RECT 608.400 415.050 609.450 484.950 ;
        RECT 610.950 481.950 613.050 484.050 ;
        RECT 614.250 482.850 615.750 483.750 ;
        RECT 616.950 481.950 619.050 484.050 ;
        RECT 611.400 481.050 612.450 481.950 ;
        RECT 610.950 478.950 613.050 481.050 ;
        RECT 568.950 412.950 571.050 415.050 ;
        RECT 572.250 413.250 573.750 414.150 ;
        RECT 574.950 412.950 577.050 415.050 ;
        RECT 578.250 413.250 580.050 414.150 ;
        RECT 580.950 412.950 583.050 415.050 ;
        RECT 607.950 412.950 610.050 415.050 ;
        RECT 613.950 412.950 616.050 415.050 ;
        RECT 569.400 409.050 570.450 412.950 ;
        RECT 571.950 409.950 574.050 412.050 ;
        RECT 575.250 410.850 576.750 411.750 ;
        RECT 577.950 411.450 580.050 412.050 ;
        RECT 581.400 411.450 582.450 412.950 ;
        RECT 577.950 410.400 582.450 411.450 ;
        RECT 577.950 409.950 580.050 410.400 ;
        RECT 610.950 410.250 613.050 411.150 ;
        RECT 613.950 410.850 616.050 411.750 ;
        RECT 568.950 406.950 571.050 409.050 ;
        RECT 565.950 394.950 568.050 397.050 ;
        RECT 544.950 388.950 547.050 391.050 ;
        RECT 553.950 389.400 556.050 391.500 ;
        RECT 545.400 385.050 546.450 388.950 ;
        RECT 538.950 384.450 541.050 385.050 ;
        RECT 538.950 383.400 543.450 384.450 ;
        RECT 538.950 382.950 541.050 383.400 ;
        RECT 538.950 380.850 541.050 381.750 ;
        RECT 526.950 351.300 529.050 353.400 ;
        RECT 527.250 347.700 528.450 351.300 ;
        RECT 526.950 345.600 529.050 347.700 ;
        RECT 542.400 346.050 543.450 383.400 ;
        RECT 544.950 382.950 547.050 385.050 ;
        RECT 544.950 380.850 547.050 381.750 ;
        RECT 554.400 372.600 555.600 389.400 ;
        RECT 572.400 388.050 573.450 409.950 ;
        RECT 610.950 406.950 613.050 409.050 ;
        RECT 574.950 389.400 577.050 391.500 ;
        RECT 559.950 385.950 562.050 388.050 ;
        RECT 571.950 385.950 574.050 388.050 ;
        RECT 560.400 385.050 561.450 385.950 ;
        RECT 559.950 382.950 562.050 385.050 ;
        RECT 565.950 382.950 568.050 385.050 ;
        RECT 559.950 380.850 562.050 381.750 ;
        RECT 565.950 380.850 568.050 381.750 ;
        RECT 575.250 377.400 576.450 389.400 ;
        RECT 611.400 388.050 612.450 406.950 ;
        RECT 623.400 394.050 624.450 520.950 ;
        RECT 628.950 490.950 631.050 493.050 ;
        RECT 625.950 457.950 628.050 460.050 ;
        RECT 626.400 457.050 627.450 457.950 ;
        RECT 625.950 454.950 628.050 457.050 ;
        RECT 625.950 452.850 628.050 453.750 ;
        RECT 622.950 391.950 625.050 394.050 ;
        RECT 613.950 388.950 616.050 391.050 ;
        RECT 577.950 386.250 580.050 387.150 ;
        RECT 580.950 385.950 583.050 388.050 ;
        RECT 610.950 385.950 613.050 388.050 ;
        RECT 577.950 384.450 580.050 385.050 ;
        RECT 581.400 384.450 582.450 385.950 ;
        RECT 614.400 385.050 615.450 388.950 ;
        RECT 577.950 383.400 582.450 384.450 ;
        RECT 577.950 382.950 580.050 383.400 ;
        RECT 589.950 382.950 592.050 385.050 ;
        RECT 613.950 382.950 616.050 385.050 ;
        RECT 619.950 384.450 622.050 385.050 ;
        RECT 619.950 383.400 624.450 384.450 ;
        RECT 619.950 382.950 622.050 383.400 ;
        RECT 574.950 375.300 577.050 377.400 ;
        RECT 553.950 370.500 556.050 372.600 ;
        RECT 575.250 371.700 576.450 375.300 ;
        RECT 574.950 369.600 577.050 371.700 ;
        RECT 518.400 335.400 522.450 336.450 ;
        RECT 505.950 331.500 508.050 333.600 ;
        RECT 478.950 310.950 481.050 313.050 ;
        RECT 482.250 311.250 483.750 312.150 ;
        RECT 484.950 310.950 487.050 313.050 ;
        RECT 478.950 308.850 480.750 309.750 ;
        RECT 481.950 307.950 484.050 310.050 ;
        RECT 485.250 308.850 486.750 309.750 ;
        RECT 487.950 307.950 490.050 310.050 ;
        RECT 487.950 305.850 490.050 306.750 ;
        RECT 514.950 274.950 517.050 277.050 ;
        RECT 478.950 271.950 481.050 274.050 ;
        RECT 490.950 271.950 493.050 274.050 ;
        RECT 479.400 264.450 480.450 271.950 ;
        RECT 491.400 271.050 492.450 271.950 ;
        RECT 515.400 271.050 516.450 274.950 ;
        RECT 518.400 271.050 519.450 335.400 ;
        RECT 527.250 333.600 528.450 345.600 ;
        RECT 541.950 343.950 544.050 346.050 ;
        RECT 590.400 343.050 591.450 382.950 ;
        RECT 613.950 380.850 616.050 381.750 ;
        RECT 619.950 380.850 622.050 381.750 ;
        RECT 610.950 346.950 613.050 349.050 ;
        RECT 589.950 340.950 592.050 343.050 ;
        RECT 529.950 337.950 532.050 340.050 ;
        RECT 568.950 338.850 571.050 339.750 ;
        RECT 571.950 337.950 574.050 340.050 ;
        RECT 589.950 338.850 592.050 339.750 ;
        RECT 529.950 335.850 532.050 336.750 ;
        RECT 565.950 334.950 568.050 337.050 ;
        RECT 526.950 331.500 529.050 333.600 ;
        RECT 520.950 319.950 523.050 322.050 ;
        RECT 521.400 306.450 522.450 319.950 ;
        RECT 523.950 308.250 525.750 309.150 ;
        RECT 526.950 307.950 529.050 310.050 ;
        RECT 566.400 309.450 567.450 334.950 ;
        RECT 572.400 316.050 573.450 337.950 ;
        RECT 611.400 316.050 612.450 346.950 ;
        RECT 571.950 313.950 574.050 316.050 ;
        RECT 610.950 315.450 613.050 316.050 ;
        RECT 610.950 314.400 615.450 315.450 ;
        RECT 610.950 313.950 613.050 314.400 ;
        RECT 568.950 311.250 571.050 312.150 ;
        RECT 571.950 311.850 574.050 312.750 ;
        RECT 607.950 311.250 610.050 312.150 ;
        RECT 610.950 311.850 613.050 312.750 ;
        RECT 568.950 309.450 571.050 310.050 ;
        RECT 530.250 308.250 532.050 309.150 ;
        RECT 566.400 308.400 571.050 309.450 ;
        RECT 568.950 307.950 571.050 308.400 ;
        RECT 607.950 307.950 610.050 310.050 ;
        RECT 523.950 306.450 526.050 307.050 ;
        RECT 521.400 305.400 526.050 306.450 ;
        RECT 527.250 305.850 528.750 306.750 ;
        RECT 523.950 304.950 526.050 305.400 ;
        RECT 484.950 269.250 487.050 270.150 ;
        RECT 490.950 268.950 493.050 271.050 ;
        RECT 514.950 268.950 517.050 271.050 ;
        RECT 517.950 268.950 520.050 271.050 ;
        RECT 481.950 266.250 483.750 267.150 ;
        RECT 484.950 265.950 487.050 268.050 ;
        RECT 490.950 266.850 493.050 267.750 ;
        RECT 481.950 264.450 484.050 265.050 ;
        RECT 479.400 263.400 484.050 264.450 ;
        RECT 481.950 262.950 484.050 263.400 ;
        RECT 469.950 239.250 472.050 240.150 ;
        RECT 517.950 238.950 520.050 241.050 ;
        RECT 469.950 235.950 472.050 238.050 ;
        RECT 508.950 236.250 510.750 237.150 ;
        RECT 511.950 235.950 514.050 238.050 ;
        RECT 515.250 236.250 517.050 237.150 ;
        RECT 470.400 235.050 471.450 235.950 ;
        RECT 464.400 233.400 468.450 234.450 ;
        RECT 457.950 229.950 460.050 232.050 ;
        RECT 451.950 202.950 454.050 205.050 ;
        RECT 445.950 169.950 448.050 172.050 ;
        RECT 446.400 169.050 447.450 169.950 ;
        RECT 452.400 169.050 453.450 202.950 ;
        RECT 458.400 196.050 459.450 229.950 ;
        RECT 457.950 193.950 460.050 196.050 ;
        RECT 464.400 186.450 465.450 233.400 ;
        RECT 469.950 232.950 472.050 235.050 ;
        RECT 508.950 232.950 511.050 235.050 ;
        RECT 512.250 233.850 513.750 234.750 ;
        RECT 514.950 234.450 517.050 235.050 ;
        RECT 518.400 234.450 519.450 238.950 ;
        RECT 514.950 233.400 519.450 234.450 ;
        RECT 514.950 232.950 517.050 233.400 ;
        RECT 511.950 202.950 514.050 205.050 ;
        RECT 512.400 202.050 513.450 202.950 ;
        RECT 466.950 200.250 469.050 201.150 ;
        RECT 478.950 199.950 481.050 202.050 ;
        RECT 502.950 199.950 505.050 202.050 ;
        RECT 511.950 199.950 514.050 202.050 ;
        RECT 515.250 200.250 516.750 201.150 ;
        RECT 517.950 199.950 520.050 202.050 ;
        RECT 466.950 196.950 469.050 199.050 ;
        RECT 470.250 197.250 471.750 198.150 ;
        RECT 472.950 196.950 475.050 199.050 ;
        RECT 476.250 197.250 478.050 198.150 ;
        RECT 467.400 190.050 468.450 196.950 ;
        RECT 479.400 196.050 480.450 199.950 ;
        RECT 487.950 196.950 490.050 199.050 ;
        RECT 469.950 193.950 472.050 196.050 ;
        RECT 473.250 194.850 474.750 195.750 ;
        RECT 475.950 193.950 478.050 196.050 ;
        RECT 478.950 193.950 481.050 196.050 ;
        RECT 466.950 187.950 469.050 190.050 ;
        RECT 464.400 185.400 468.450 186.450 ;
        RECT 445.950 166.950 448.050 169.050 ;
        RECT 449.250 167.250 450.750 168.150 ;
        RECT 451.950 166.950 454.050 169.050 ;
        RECT 445.950 164.850 447.750 165.750 ;
        RECT 448.950 163.950 451.050 166.050 ;
        RECT 452.250 164.850 453.750 165.750 ;
        RECT 454.950 163.950 457.050 166.050 ;
        RECT 448.950 160.950 451.050 163.050 ;
        RECT 454.950 161.850 457.050 162.750 ;
        RECT 442.950 97.950 445.050 100.050 ;
        RECT 442.950 95.850 445.050 96.750 ;
        RECT 445.950 95.250 448.050 96.150 ;
        RECT 445.950 93.450 448.050 94.050 ;
        RECT 449.400 93.450 450.450 160.950 ;
        RECT 467.400 130.050 468.450 185.400 ;
        RECT 478.950 172.950 481.050 175.050 ;
        RECT 472.950 131.250 475.050 132.150 ;
        RECT 466.950 127.950 469.050 130.050 ;
        RECT 470.250 128.250 471.750 129.150 ;
        RECT 472.950 127.950 475.050 130.050 ;
        RECT 476.250 128.250 478.050 129.150 ;
        RECT 466.950 125.850 468.750 126.750 ;
        RECT 469.950 124.950 472.050 127.050 ;
        RECT 475.950 126.450 478.050 127.050 ;
        RECT 479.400 126.450 480.450 172.950 ;
        RECT 475.950 125.400 480.450 126.450 ;
        RECT 475.950 124.950 478.050 125.400 ;
        RECT 488.400 118.050 489.450 196.950 ;
        RECT 490.950 187.950 493.050 190.050 ;
        RECT 491.400 166.050 492.450 187.950 ;
        RECT 496.950 166.950 499.050 169.050 ;
        RECT 497.400 166.050 498.450 166.950 ;
        RECT 490.950 163.950 493.050 166.050 ;
        RECT 496.950 163.950 499.050 166.050 ;
        RECT 500.250 164.250 502.050 165.150 ;
        RECT 490.950 161.850 492.750 162.750 ;
        RECT 493.950 160.950 496.050 163.050 ;
        RECT 497.250 161.850 498.750 162.750 ;
        RECT 499.950 162.450 502.050 163.050 ;
        RECT 503.400 162.450 504.450 199.950 ;
        RECT 511.950 197.850 513.750 198.750 ;
        RECT 514.950 196.950 517.050 199.050 ;
        RECT 518.250 197.850 520.050 198.750 ;
        RECT 520.950 187.950 523.050 190.050 ;
        RECT 511.950 166.950 514.050 169.050 ;
        RECT 499.950 161.400 504.450 162.450 ;
        RECT 499.950 160.950 502.050 161.400 ;
        RECT 505.950 160.950 508.050 163.050 ;
        RECT 493.950 158.850 496.050 159.750 ;
        RECT 506.400 123.450 507.450 160.950 ;
        RECT 512.400 127.050 513.450 166.950 ;
        RECT 517.950 128.250 520.050 129.150 ;
        RECT 508.950 125.250 510.750 126.150 ;
        RECT 511.950 124.950 514.050 127.050 ;
        RECT 517.950 126.450 520.050 127.050 ;
        RECT 521.400 126.450 522.450 187.950 ;
        RECT 524.400 163.050 525.450 304.950 ;
        RECT 577.950 277.950 580.050 280.050 ;
        RECT 589.950 278.400 592.050 280.500 ;
        RECT 535.950 274.950 538.050 277.050 ;
        RECT 536.400 274.050 537.450 274.950 ;
        RECT 529.950 271.950 532.050 274.050 ;
        RECT 533.250 272.250 534.750 273.150 ;
        RECT 535.950 271.950 538.050 274.050 ;
        RECT 571.950 272.250 574.050 273.150 ;
        RECT 578.400 271.050 579.450 277.950 ;
        RECT 529.950 269.850 531.750 270.750 ;
        RECT 532.950 268.950 535.050 271.050 ;
        RECT 536.250 269.850 538.050 270.750 ;
        RECT 571.950 268.950 574.050 271.050 ;
        RECT 575.250 269.250 576.750 270.150 ;
        RECT 577.950 268.950 580.050 271.050 ;
        RECT 581.250 269.250 583.050 270.150 ;
        RECT 572.400 265.050 573.450 268.950 ;
        RECT 574.950 265.950 577.050 268.050 ;
        RECT 578.250 266.850 579.750 267.750 ;
        RECT 580.950 265.950 583.050 268.050 ;
        RECT 575.400 265.050 576.450 265.950 ;
        RECT 571.950 262.950 574.050 265.050 ;
        RECT 574.950 262.950 577.050 265.050 ;
        RECT 590.400 261.600 591.600 278.400 ;
        RECT 595.950 269.250 598.050 270.150 ;
        RECT 601.950 269.250 604.050 270.150 ;
        RECT 608.400 268.050 609.450 307.950 ;
        RECT 610.950 279.300 613.050 281.400 ;
        RECT 611.250 275.700 612.450 279.300 ;
        RECT 610.950 273.600 613.050 275.700 ;
        RECT 595.950 265.950 598.050 268.050 ;
        RECT 601.950 265.950 604.050 268.050 ;
        RECT 607.950 265.950 610.050 268.050 ;
        RECT 596.400 265.050 597.450 265.950 ;
        RECT 602.400 265.050 603.450 265.950 ;
        RECT 595.950 262.950 598.050 265.050 ;
        RECT 601.950 262.950 604.050 265.050 ;
        RECT 611.250 261.600 612.450 273.600 ;
        RECT 614.400 268.050 615.450 314.400 ;
        RECT 623.400 274.050 624.450 383.400 ;
        RECT 629.400 349.050 630.450 490.950 ;
        RECT 632.400 487.050 633.450 557.400 ;
        RECT 646.950 556.950 649.050 559.050 ;
        RECT 656.400 553.050 657.450 670.950 ;
        RECT 665.400 670.050 666.450 670.950 ;
        RECT 701.400 670.050 702.450 673.950 ;
        RECT 703.950 672.450 706.050 673.050 ;
        RECT 706.950 672.450 709.050 673.050 ;
        RECT 703.950 671.400 709.050 672.450 ;
        RECT 703.950 670.950 706.050 671.400 ;
        RECT 706.950 670.950 709.050 671.400 ;
        RECT 710.250 671.250 711.750 672.150 ;
        RECT 712.950 670.950 715.050 673.050 ;
        RECT 664.950 667.950 667.050 670.050 ;
        RECT 668.250 668.850 669.750 669.750 ;
        RECT 670.950 667.950 673.050 670.050 ;
        RECT 674.250 668.850 676.050 669.750 ;
        RECT 700.950 667.950 703.050 670.050 ;
        RECT 664.950 665.850 667.050 666.750 ;
        RECT 664.950 637.950 667.050 640.050 ;
        RECT 658.950 632.250 661.050 633.150 ;
        RECT 665.400 631.050 666.450 637.950 ;
        RECT 658.950 628.950 661.050 631.050 ;
        RECT 662.250 629.250 663.750 630.150 ;
        RECT 664.950 628.950 667.050 631.050 ;
        RECT 668.250 629.250 670.050 630.150 ;
        RECT 700.950 629.250 703.050 630.150 ;
        RECT 661.950 625.950 664.050 628.050 ;
        RECT 665.250 626.850 666.750 627.750 ;
        RECT 667.950 625.950 670.050 628.050 ;
        RECT 704.400 627.450 705.450 670.950 ;
        RECT 706.950 668.850 708.750 669.750 ;
        RECT 709.950 667.950 712.050 670.050 ;
        RECT 713.250 668.850 714.750 669.750 ;
        RECT 715.950 669.450 718.050 670.050 ;
        RECT 715.950 668.400 720.450 669.450 ;
        RECT 715.950 667.950 718.050 668.400 ;
        RECT 715.950 665.850 718.050 666.750 ;
        RECT 706.950 629.250 709.050 630.150 ;
        RECT 706.950 627.450 709.050 628.050 ;
        RECT 704.400 626.400 709.050 627.450 ;
        RECT 706.950 625.950 709.050 626.400 ;
        RECT 668.400 625.050 669.450 625.950 ;
        RECT 661.950 622.950 664.050 625.050 ;
        RECT 667.950 622.950 670.050 625.050 ;
        RECT 682.950 622.950 685.050 625.050 ;
        RECT 662.400 562.050 663.450 622.950 ;
        RECT 683.400 601.050 684.450 622.950 ;
        RECT 682.950 598.950 685.050 601.050 ;
        RECT 685.950 598.950 688.050 601.050 ;
        RECT 682.950 596.850 685.050 597.750 ;
        RECT 661.950 561.450 664.050 562.050 ;
        RECT 659.400 560.400 664.050 561.450 ;
        RECT 655.950 550.950 658.050 553.050 ;
        RECT 659.400 523.050 660.450 560.400 ;
        RECT 661.950 559.950 664.050 560.400 ;
        RECT 665.250 560.250 666.750 561.150 ;
        RECT 667.950 559.950 670.050 562.050 ;
        RECT 676.950 559.950 679.050 562.050 ;
        RECT 661.950 557.850 663.750 558.750 ;
        RECT 664.950 556.950 667.050 559.050 ;
        RECT 668.250 557.850 670.050 558.750 ;
        RECT 664.950 550.950 667.050 553.050 ;
        RECT 665.400 526.050 666.450 550.950 ;
        RECT 670.950 529.950 673.050 532.050 ;
        RECT 661.950 524.250 663.750 525.150 ;
        RECT 664.950 523.950 667.050 526.050 ;
        RECT 668.250 524.250 670.050 525.150 ;
        RECT 658.950 520.950 661.050 523.050 ;
        RECT 661.950 520.950 664.050 523.050 ;
        RECT 665.250 521.850 666.750 522.750 ;
        RECT 667.950 520.950 670.050 523.050 ;
        RECT 662.400 493.050 663.450 520.950 ;
        RECT 661.950 490.950 664.050 493.050 ;
        RECT 671.400 490.050 672.450 529.950 ;
        RECT 640.950 487.950 643.050 490.050 ;
        RECT 658.950 487.950 661.050 490.050 ;
        RECT 662.250 488.250 663.750 489.150 ;
        RECT 664.950 487.950 667.050 490.050 ;
        RECT 670.950 487.950 673.050 490.050 ;
        RECT 631.950 484.950 634.050 487.050 ;
        RECT 631.950 454.950 634.050 457.050 ;
        RECT 631.950 452.850 634.050 453.750 ;
        RECT 631.950 389.400 634.050 391.500 ;
        RECT 632.400 372.600 633.600 389.400 ;
        RECT 637.950 388.950 640.050 391.050 ;
        RECT 638.400 385.050 639.450 388.950 ;
        RECT 637.950 382.950 640.050 385.050 ;
        RECT 637.950 380.850 640.050 381.750 ;
        RECT 631.950 370.500 634.050 372.600 ;
        RECT 628.950 346.950 631.050 349.050 ;
        RECT 641.400 346.050 642.450 487.950 ;
        RECT 658.950 485.850 660.750 486.750 ;
        RECT 661.950 484.950 664.050 487.050 ;
        RECT 665.250 485.850 667.050 486.750 ;
        RECT 671.400 481.050 672.450 487.950 ;
        RECT 670.950 478.950 673.050 481.050 ;
        RECT 670.950 475.950 673.050 478.050 ;
        RECT 671.400 460.050 672.450 475.950 ;
        RECT 670.950 457.950 673.050 460.050 ;
        RECT 658.950 454.950 661.050 457.050 ;
        RECT 667.950 455.250 670.050 456.150 ;
        RECT 670.950 455.850 673.050 456.750 ;
        RECT 649.950 421.950 652.050 424.050 ;
        RECT 650.400 414.450 651.450 421.950 ;
        RECT 652.950 416.250 655.050 417.150 ;
        RECT 659.400 415.050 660.450 454.950 ;
        RECT 667.950 451.950 670.050 454.050 ;
        RECT 668.400 451.050 669.450 451.950 ;
        RECT 667.950 448.950 670.050 451.050 ;
        RECT 652.950 414.450 655.050 415.050 ;
        RECT 650.400 413.400 655.050 414.450 ;
        RECT 652.950 412.950 655.050 413.400 ;
        RECT 656.250 413.250 657.750 414.150 ;
        RECT 658.950 412.950 661.050 415.050 ;
        RECT 662.250 413.250 664.050 414.150 ;
        RECT 655.950 409.950 658.050 412.050 ;
        RECT 659.250 410.850 660.750 411.750 ;
        RECT 661.950 409.950 664.050 412.050 ;
        RECT 652.950 389.400 655.050 391.500 ;
        RECT 656.400 391.050 657.450 409.950 ;
        RECT 643.950 382.950 646.050 385.050 ;
        RECT 649.950 382.950 652.050 385.050 ;
        RECT 643.950 380.850 646.050 381.750 ;
        RECT 643.950 351.300 646.050 353.400 ;
        RECT 644.550 347.700 645.750 351.300 ;
        RECT 625.950 343.950 628.050 346.050 ;
        RECT 628.950 343.950 631.050 346.050 ;
        RECT 632.250 344.250 633.750 345.150 ;
        RECT 634.950 343.950 637.050 346.050 ;
        RECT 640.950 343.950 643.050 346.050 ;
        RECT 643.950 345.600 646.050 347.700 ;
        RECT 626.400 313.050 627.450 343.950 ;
        RECT 628.950 341.850 630.750 342.750 ;
        RECT 631.950 340.950 634.050 343.050 ;
        RECT 635.250 341.850 637.050 342.750 ;
        RECT 625.950 310.950 628.050 313.050 ;
        RECT 622.950 271.950 625.050 274.050 ;
        RECT 626.400 271.050 627.450 310.950 ;
        RECT 632.400 310.050 633.450 340.950 ;
        RECT 641.400 340.050 642.450 343.950 ;
        RECT 640.950 337.950 643.050 340.050 ;
        RECT 640.950 335.850 643.050 336.750 ;
        RECT 644.550 333.600 645.750 345.600 ;
        RECT 646.950 337.950 649.050 340.050 ;
        RECT 650.400 339.450 651.450 382.950 ;
        RECT 653.250 377.400 654.450 389.400 ;
        RECT 655.950 388.950 658.050 391.050 ;
        RECT 655.950 386.250 658.050 387.150 ;
        RECT 658.950 385.950 661.050 388.050 ;
        RECT 655.950 384.450 658.050 385.050 ;
        RECT 659.400 384.450 660.450 385.950 ;
        RECT 655.950 383.400 660.450 384.450 ;
        RECT 655.950 382.950 658.050 383.400 ;
        RECT 662.400 379.050 663.450 409.950 ;
        RECT 652.950 375.300 655.050 377.400 ;
        RECT 661.950 376.950 664.050 379.050 ;
        RECT 653.250 371.700 654.450 375.300 ;
        RECT 652.950 369.600 655.050 371.700 ;
        RECT 664.950 350.400 667.050 352.500 ;
        RECT 652.950 341.250 655.050 342.150 ;
        RECT 658.950 341.250 661.050 342.150 ;
        RECT 652.950 339.450 655.050 340.050 ;
        RECT 650.400 338.400 655.050 339.450 ;
        RECT 652.950 337.950 655.050 338.400 ;
        RECT 658.950 337.950 661.050 340.050 ;
        RECT 643.950 331.500 646.050 333.600 ;
        RECT 647.400 313.050 648.450 337.950 ;
        RECT 653.400 316.050 654.450 337.950 ;
        RECT 665.400 333.600 666.600 350.400 ;
        RECT 664.950 331.500 667.050 333.600 ;
        RECT 661.950 317.400 664.050 319.500 ;
        RECT 652.950 313.950 655.050 316.050 ;
        RECT 646.950 310.950 649.050 313.050 ;
        RECT 650.250 311.250 651.750 312.150 ;
        RECT 652.950 310.950 655.050 313.050 ;
        RECT 658.950 310.950 661.050 313.050 ;
        RECT 631.950 307.950 634.050 310.050 ;
        RECT 643.950 307.950 646.050 310.050 ;
        RECT 647.250 308.850 648.750 309.750 ;
        RECT 649.950 307.950 652.050 310.050 ;
        RECT 653.250 308.850 655.050 309.750 ;
        RECT 643.950 305.850 646.050 306.750 ;
        RECT 650.400 304.050 651.450 307.950 ;
        RECT 643.950 301.950 646.050 304.050 ;
        RECT 649.950 301.950 652.050 304.050 ;
        RECT 625.950 268.950 628.050 271.050 ;
        RECT 613.950 265.950 616.050 268.050 ;
        RECT 613.950 263.850 616.050 264.750 ;
        RECT 589.950 259.500 592.050 261.600 ;
        RECT 610.950 259.500 613.050 261.600 ;
        RECT 626.400 244.050 627.450 268.950 ;
        RECT 547.950 241.950 550.050 244.050 ;
        RECT 568.950 241.950 571.050 244.050 ;
        RECT 586.950 241.950 589.050 244.050 ;
        RECT 625.950 241.950 628.050 244.050 ;
        RECT 547.950 239.850 550.050 240.750 ;
        RECT 550.950 239.250 553.050 240.150 ;
        RECT 550.950 235.950 553.050 238.050 ;
        RECT 551.400 232.050 552.450 235.950 ;
        RECT 550.950 229.950 553.050 232.050 ;
        RECT 547.950 226.950 550.050 229.050 ;
        RECT 548.400 199.050 549.450 226.950 ;
        RECT 553.950 203.250 556.050 204.150 ;
        RECT 550.950 200.250 552.750 201.150 ;
        RECT 553.950 199.950 556.050 202.050 ;
        RECT 557.250 200.250 558.750 201.150 ;
        RECT 559.950 199.950 562.050 202.050 ;
        RECT 554.400 199.050 555.450 199.950 ;
        RECT 569.400 199.050 570.450 241.950 ;
        RECT 587.400 241.050 588.450 241.950 ;
        RECT 586.950 238.950 589.050 241.050 ;
        RECT 590.250 239.250 591.750 240.150 ;
        RECT 592.950 238.950 595.050 241.050 ;
        RECT 586.950 236.850 588.750 237.750 ;
        RECT 589.950 235.950 592.050 238.050 ;
        RECT 593.250 236.850 594.750 237.750 ;
        RECT 595.950 235.950 598.050 238.050 ;
        RECT 626.400 235.050 627.450 241.950 ;
        RECT 631.950 236.250 633.750 237.150 ;
        RECT 634.950 235.950 637.050 238.050 ;
        RECT 638.250 236.250 640.050 237.150 ;
        RECT 595.950 233.850 598.050 234.750 ;
        RECT 625.950 232.950 628.050 235.050 ;
        RECT 631.950 232.950 634.050 235.050 ;
        RECT 635.250 233.850 636.750 234.750 ;
        RECT 637.950 232.950 640.050 235.050 ;
        RECT 574.950 229.950 577.050 232.050 ;
        RECT 571.950 207.300 574.050 209.400 ;
        RECT 572.550 203.700 573.750 207.300 ;
        RECT 571.950 201.600 574.050 203.700 ;
        RECT 547.950 196.950 550.050 199.050 ;
        RECT 550.950 196.950 553.050 199.050 ;
        RECT 553.950 196.950 556.050 199.050 ;
        RECT 556.950 196.950 559.050 199.050 ;
        RECT 560.250 197.850 562.050 198.750 ;
        RECT 568.950 196.950 571.050 199.050 ;
        RECT 551.400 190.050 552.450 196.950 ;
        RECT 554.400 196.050 555.450 196.950 ;
        RECT 553.950 193.950 556.050 196.050 ;
        RECT 550.950 187.950 553.050 190.050 ;
        RECT 538.950 166.950 541.050 169.050 ;
        RECT 539.400 166.050 540.450 166.950 ;
        RECT 535.950 164.250 537.750 165.150 ;
        RECT 538.950 163.950 541.050 166.050 ;
        RECT 542.250 164.250 544.050 165.150 ;
        RECT 523.950 160.950 526.050 163.050 ;
        RECT 539.250 161.850 540.750 162.750 ;
        RECT 541.950 160.950 544.050 163.050 ;
        RECT 515.250 125.250 516.750 126.150 ;
        RECT 517.950 125.400 522.450 126.450 ;
        RECT 517.950 124.950 520.050 125.400 ;
        RECT 508.950 123.450 511.050 124.050 ;
        RECT 506.400 122.400 511.050 123.450 ;
        RECT 512.250 122.850 513.750 123.750 ;
        RECT 487.950 115.950 490.050 118.050 ;
        RECT 484.950 109.950 487.050 112.050 ;
        RECT 460.950 100.950 463.050 103.050 ;
        RECT 445.950 92.400 450.450 93.450 ;
        RECT 445.950 91.950 448.050 92.400 ;
        RECT 446.400 64.050 447.450 91.950 ;
        RECT 445.950 61.950 448.050 64.050 ;
        RECT 448.950 63.300 451.050 65.400 ;
        RECT 449.550 59.700 450.750 63.300 ;
        RECT 439.950 55.950 442.050 58.050 ;
        RECT 448.950 57.600 451.050 59.700 ;
        RECT 436.950 52.950 439.050 55.050 ;
        RECT 437.400 52.050 438.450 52.950 ;
        RECT 436.950 49.950 439.050 52.050 ;
        RECT 445.950 49.950 448.050 52.050 ;
        RECT 436.950 47.850 439.050 48.750 ;
        RECT 445.950 47.850 448.050 48.750 ;
        RECT 449.550 45.600 450.750 57.600 ;
        RECT 457.950 53.250 460.050 54.150 ;
        RECT 457.950 51.450 460.050 52.050 ;
        RECT 461.400 51.450 462.450 100.950 ;
        RECT 478.950 95.850 481.050 96.750 ;
        RECT 481.950 95.250 484.050 96.150 ;
        RECT 481.950 93.450 484.050 94.050 ;
        RECT 485.400 93.450 486.450 109.950 ;
        RECT 488.400 96.450 489.450 115.950 ;
        RECT 493.950 101.400 496.050 103.500 ;
        RECT 490.950 98.250 493.050 99.150 ;
        RECT 490.950 96.450 493.050 97.050 ;
        RECT 488.400 95.400 493.050 96.450 ;
        RECT 490.950 94.950 493.050 95.400 ;
        RECT 481.950 92.400 486.450 93.450 ;
        RECT 481.950 91.950 484.050 92.400 ;
        RECT 494.550 89.400 495.750 101.400 ;
        RECT 502.950 100.950 505.050 103.050 ;
        RECT 503.400 97.050 504.450 100.950 ;
        RECT 506.400 100.050 507.450 122.400 ;
        RECT 508.950 121.950 511.050 122.400 ;
        RECT 514.950 121.950 517.050 124.050 ;
        RECT 515.400 121.050 516.450 121.950 ;
        RECT 514.950 118.950 517.050 121.050 ;
        RECT 514.950 101.400 517.050 103.500 ;
        RECT 505.950 97.950 508.050 100.050 ;
        RECT 502.950 94.950 505.050 97.050 ;
        RECT 508.950 96.450 511.050 97.050 ;
        RECT 508.950 95.400 513.450 96.450 ;
        RECT 508.950 94.950 511.050 95.400 ;
        RECT 502.950 92.850 505.050 93.750 ;
        RECT 508.950 92.850 511.050 93.750 ;
        RECT 512.400 91.050 513.450 95.400 ;
        RECT 493.950 87.300 496.050 89.400 ;
        RECT 511.950 88.950 514.050 91.050 ;
        RECT 494.550 83.700 495.750 87.300 ;
        RECT 515.400 84.600 516.600 101.400 ;
        RECT 542.400 97.050 543.450 160.950 ;
        RECT 553.950 124.950 556.050 127.050 ;
        RECT 550.950 122.250 553.050 123.150 ;
        RECT 553.950 122.850 556.050 123.750 ;
        RECT 550.950 118.950 553.050 121.050 ;
        RECT 551.400 118.050 552.450 118.950 ;
        RECT 557.400 118.050 558.450 196.950 ;
        RECT 569.400 196.050 570.450 196.950 ;
        RECT 568.950 193.950 571.050 196.050 ;
        RECT 568.950 191.850 571.050 192.750 ;
        RECT 572.550 189.600 573.750 201.600 ;
        RECT 571.950 187.500 574.050 189.600 ;
        RECT 575.400 166.050 576.450 229.950 ;
        RECT 592.950 206.400 595.050 208.500 ;
        RECT 580.950 197.250 583.050 198.150 ;
        RECT 586.950 197.250 589.050 198.150 ;
        RECT 580.950 193.950 583.050 196.050 ;
        RECT 586.950 193.950 589.050 196.050 ;
        RECT 587.400 193.050 588.450 193.950 ;
        RECT 580.950 190.950 583.050 193.050 ;
        RECT 586.950 190.950 589.050 193.050 ;
        RECT 581.400 169.050 582.450 190.950 ;
        RECT 593.400 189.600 594.600 206.400 ;
        RECT 625.950 202.950 628.050 205.050 ;
        RECT 637.950 202.950 640.050 205.050 ;
        RECT 592.950 187.500 595.050 189.600 ;
        RECT 619.950 169.950 622.050 172.050 ;
        RECT 620.400 169.050 621.450 169.950 ;
        RECT 626.400 169.050 627.450 202.950 ;
        RECT 638.400 202.050 639.450 202.950 ;
        RECT 631.950 199.950 634.050 202.050 ;
        RECT 635.250 200.250 636.750 201.150 ;
        RECT 637.950 199.950 640.050 202.050 ;
        RECT 631.950 197.850 633.750 198.750 ;
        RECT 634.950 196.950 637.050 199.050 ;
        RECT 638.250 197.850 640.050 198.750 ;
        RECT 577.950 166.950 580.050 169.050 ;
        RECT 580.950 166.950 583.050 169.050 ;
        RECT 586.950 168.450 589.050 169.050 ;
        RECT 584.250 167.250 585.750 168.150 ;
        RECT 586.950 167.400 591.450 168.450 ;
        RECT 586.950 166.950 589.050 167.400 ;
        RECT 578.400 166.050 579.450 166.950 ;
        RECT 574.950 163.950 577.050 166.050 ;
        RECT 577.950 163.950 580.050 166.050 ;
        RECT 581.250 164.850 582.750 165.750 ;
        RECT 583.950 163.950 586.050 166.050 ;
        RECT 587.250 164.850 589.050 165.750 ;
        RECT 590.400 163.050 591.450 167.400 ;
        RECT 619.950 166.950 622.050 169.050 ;
        RECT 623.250 167.250 624.750 168.150 ;
        RECT 625.950 166.950 628.050 169.050 ;
        RECT 619.950 164.850 621.750 165.750 ;
        RECT 622.950 163.950 625.050 166.050 ;
        RECT 626.250 164.850 627.750 165.750 ;
        RECT 628.950 165.450 631.050 166.050 ;
        RECT 628.950 164.400 633.450 165.450 ;
        RECT 628.950 163.950 631.050 164.400 ;
        RECT 577.950 161.850 580.050 162.750 ;
        RECT 589.950 160.950 592.050 163.050 ;
        RECT 610.950 160.950 613.050 163.050 ;
        RECT 628.950 161.850 631.050 162.750 ;
        RECT 559.950 157.950 562.050 160.050 ;
        RECT 560.400 127.050 561.450 157.950 ;
        RECT 589.950 129.450 592.050 130.050 ;
        RECT 587.400 128.400 592.050 129.450 ;
        RECT 595.950 129.450 598.050 130.050 ;
        RECT 559.950 124.950 562.050 127.050 ;
        RECT 550.950 115.950 553.050 118.050 ;
        RECT 556.950 115.950 559.050 118.050 ;
        RECT 560.400 100.050 561.450 124.950 ;
        RECT 587.400 124.050 588.450 128.400 ;
        RECT 589.950 127.950 592.050 128.400 ;
        RECT 593.250 128.250 594.750 129.150 ;
        RECT 595.950 128.400 600.450 129.450 ;
        RECT 595.950 127.950 598.050 128.400 ;
        RECT 589.950 125.850 591.750 126.750 ;
        RECT 592.950 124.950 595.050 127.050 ;
        RECT 596.250 125.850 598.050 126.750 ;
        RECT 586.950 121.950 589.050 124.050 ;
        RECT 559.950 97.950 562.050 100.050 ;
        RECT 541.950 94.950 544.050 97.050 ;
        RECT 553.950 94.950 556.050 97.050 ;
        RECT 557.250 95.250 558.750 96.150 ;
        RECT 559.950 94.950 562.050 97.050 ;
        RECT 565.950 94.950 568.050 97.050 ;
        RECT 553.950 92.850 555.750 93.750 ;
        RECT 556.950 91.950 559.050 94.050 ;
        RECT 560.250 92.850 561.750 93.750 ;
        RECT 562.950 91.950 565.050 94.050 ;
        RECT 566.400 91.050 567.450 94.950 ;
        RECT 562.950 89.850 565.050 90.750 ;
        RECT 565.950 88.950 568.050 91.050 ;
        RECT 493.950 81.600 496.050 83.700 ;
        RECT 514.950 82.500 517.050 84.600 ;
        RECT 587.400 79.050 588.450 121.950 ;
        RECT 599.400 121.050 600.450 128.400 ;
        RECT 598.950 118.950 601.050 121.050 ;
        RECT 601.950 92.250 603.750 93.150 ;
        RECT 604.950 91.950 607.050 94.050 ;
        RECT 608.250 92.250 610.050 93.150 ;
        RECT 605.250 89.850 606.750 90.750 ;
        RECT 607.950 90.450 610.050 91.050 ;
        RECT 611.400 90.450 612.450 160.950 ;
        RECT 632.400 160.050 633.450 164.400 ;
        RECT 631.950 157.950 634.050 160.050 ;
        RECT 637.950 127.950 640.050 130.050 ;
        RECT 638.400 127.050 639.450 127.950 ;
        RECT 631.950 125.250 634.050 126.150 ;
        RECT 637.950 124.950 640.050 127.050 ;
        RECT 644.400 124.050 645.450 301.950 ;
        RECT 659.400 294.450 660.450 310.950 ;
        RECT 662.400 300.600 663.600 317.400 ;
        RECT 664.950 313.950 667.050 316.050 ;
        RECT 673.950 313.950 676.050 316.050 ;
        RECT 661.950 298.500 664.050 300.600 ;
        RECT 659.400 293.400 663.450 294.450 ;
        RECT 658.950 272.250 661.050 273.150 ;
        RECT 649.950 269.250 651.750 270.150 ;
        RECT 652.950 268.950 655.050 271.050 ;
        RECT 656.250 269.250 657.750 270.150 ;
        RECT 658.950 268.950 661.050 271.050 ;
        RECT 662.400 268.050 663.450 293.400 ;
        RECT 665.400 268.050 666.450 313.950 ;
        RECT 674.400 313.050 675.450 313.950 ;
        RECT 667.950 310.950 670.050 313.050 ;
        RECT 673.950 310.950 676.050 313.050 ;
        RECT 667.950 308.850 670.050 309.750 ;
        RECT 673.950 308.850 676.050 309.750 ;
        RECT 649.950 265.950 652.050 268.050 ;
        RECT 653.250 266.850 654.750 267.750 ;
        RECT 655.950 265.950 658.050 268.050 ;
        RECT 661.950 265.950 664.050 268.050 ;
        RECT 664.950 265.950 667.050 268.050 ;
        RECT 646.950 245.400 649.050 247.500 ;
        RECT 647.400 228.600 648.600 245.400 ;
        RECT 650.400 232.050 651.450 265.950 ;
        RECT 665.400 265.050 666.450 265.950 ;
        RECT 664.950 262.950 667.050 265.050 ;
        RECT 665.400 241.050 666.450 262.950 ;
        RECT 667.950 245.400 670.050 247.500 ;
        RECT 652.950 238.950 655.050 241.050 ;
        RECT 658.950 238.950 661.050 241.050 ;
        RECT 664.950 238.950 667.050 241.050 ;
        RECT 652.950 236.850 655.050 237.750 ;
        RECT 658.950 236.850 661.050 237.750 ;
        RECT 668.250 233.400 669.450 245.400 ;
        RECT 670.950 242.250 673.050 243.150 ;
        RECT 670.950 238.950 673.050 241.050 ;
        RECT 671.400 235.050 672.450 238.950 ;
        RECT 649.950 229.950 652.050 232.050 ;
        RECT 667.950 231.300 670.050 233.400 ;
        RECT 670.950 232.950 673.050 235.050 ;
        RECT 646.950 226.500 649.050 228.600 ;
        RECT 668.250 227.700 669.450 231.300 ;
        RECT 667.950 225.600 670.050 227.700 ;
        RECT 649.950 206.400 652.050 208.500 ;
        RECT 670.950 207.300 673.050 209.400 ;
        RECT 650.400 189.600 651.600 206.400 ;
        RECT 671.250 203.700 672.450 207.300 ;
        RECT 670.950 201.600 673.050 203.700 ;
        RECT 655.950 197.250 658.050 198.150 ;
        RECT 661.950 197.250 664.050 198.150 ;
        RECT 655.950 193.950 658.050 196.050 ;
        RECT 661.950 193.950 664.050 196.050 ;
        RECT 656.400 193.050 657.450 193.950 ;
        RECT 655.950 190.950 658.050 193.050 ;
        RECT 649.950 187.500 652.050 189.600 ;
        RECT 628.950 122.250 630.750 123.150 ;
        RECT 631.950 121.950 634.050 124.050 ;
        RECT 637.950 122.850 640.050 123.750 ;
        RECT 643.950 121.950 646.050 124.050 ;
        RECT 628.950 118.950 631.050 121.050 ;
        RECT 662.400 103.050 663.450 193.950 ;
        RECT 667.950 190.950 670.050 193.050 ;
        RECT 668.400 166.050 669.450 190.950 ;
        RECT 671.250 189.600 672.450 201.600 ;
        RECT 673.950 195.450 676.050 196.050 ;
        RECT 677.400 195.450 678.450 559.950 ;
        RECT 686.400 556.050 687.450 598.950 ;
        RECT 688.950 596.850 691.050 597.750 ;
        RECT 700.950 557.250 703.050 558.150 ;
        RECT 706.950 557.250 709.050 558.150 ;
        RECT 685.950 553.950 688.050 556.050 ;
        RECT 706.950 553.950 709.050 556.050 ;
        RECT 709.950 553.950 712.050 556.050 ;
        RECT 707.400 532.050 708.450 553.950 ;
        RECT 700.950 529.950 703.050 532.050 ;
        RECT 706.950 529.950 709.050 532.050 ;
        RECT 701.400 529.050 702.450 529.950 ;
        RECT 700.950 526.950 703.050 529.050 ;
        RECT 706.950 528.450 709.050 529.050 ;
        RECT 710.400 528.450 711.450 553.950 ;
        RECT 719.400 553.050 720.450 668.400 ;
        RECT 721.950 598.950 724.050 601.050 ;
        RECT 721.950 596.850 724.050 597.750 ;
        RECT 727.950 596.850 730.050 597.750 ;
        RECT 718.950 550.950 721.050 553.050 ;
        RECT 704.250 527.250 705.750 528.150 ;
        RECT 706.950 527.400 711.450 528.450 ;
        RECT 706.950 526.950 709.050 527.400 ;
        RECT 733.950 526.950 736.050 529.050 ;
        RECT 700.950 524.850 702.750 525.750 ;
        RECT 703.950 523.950 706.050 526.050 ;
        RECT 707.250 524.850 708.750 525.750 ;
        RECT 709.950 523.950 712.050 526.050 ;
        RECT 715.950 523.950 718.050 526.050 ;
        RECT 709.950 521.850 712.050 522.750 ;
        RECT 688.950 514.950 691.050 517.050 ;
        RECT 682.950 317.400 685.050 319.500 ;
        RECT 683.250 305.400 684.450 317.400 ;
        RECT 685.950 314.250 688.050 315.150 ;
        RECT 685.950 310.950 688.050 313.050 ;
        RECT 682.950 303.300 685.050 305.400 ;
        RECT 683.250 299.700 684.450 303.300 ;
        RECT 682.950 297.600 685.050 299.700 ;
        RECT 673.950 194.400 678.450 195.450 ;
        RECT 673.950 193.950 676.050 194.400 ;
        RECT 673.950 191.850 676.050 192.750 ;
        RECT 670.950 187.500 673.050 189.600 ;
        RECT 664.950 164.250 666.750 165.150 ;
        RECT 667.950 163.950 670.050 166.050 ;
        RECT 671.250 164.250 673.050 165.150 ;
        RECT 673.950 163.950 676.050 166.050 ;
        RECT 664.950 160.950 667.050 163.050 ;
        RECT 668.250 161.850 669.750 162.750 ;
        RECT 670.950 162.450 673.050 163.050 ;
        RECT 674.400 162.450 675.450 163.950 ;
        RECT 677.400 163.050 678.450 194.400 ;
        RECT 670.950 161.400 675.450 162.450 ;
        RECT 670.950 160.950 673.050 161.400 ;
        RECT 676.950 160.950 679.050 163.050 ;
        RECT 665.400 157.050 666.450 160.950 ;
        RECT 664.950 154.950 667.050 157.050 ;
        RECT 673.950 129.450 676.050 130.050 ;
        RECT 671.400 128.400 676.050 129.450 ;
        RECT 671.400 127.050 672.450 128.400 ;
        RECT 673.950 127.950 676.050 128.400 ;
        RECT 677.250 128.250 678.750 129.150 ;
        RECT 679.950 127.950 682.050 130.050 ;
        RECT 689.400 127.050 690.450 514.950 ;
        RECT 697.950 485.250 700.050 486.150 ;
        RECT 703.950 485.250 706.050 486.150 ;
        RECT 697.950 483.450 700.050 484.050 ;
        RECT 697.950 482.400 702.450 483.450 ;
        RECT 697.950 481.950 700.050 482.400 ;
        RECT 691.950 413.250 694.050 414.150 ;
        RECT 697.950 413.250 700.050 414.150 ;
        RECT 697.950 409.950 700.050 412.050 ;
        RECT 698.400 391.050 699.450 409.950 ;
        RECT 701.400 409.050 702.450 482.400 ;
        RECT 703.950 478.950 706.050 481.050 ;
        RECT 704.400 450.450 705.450 478.950 ;
        RECT 706.950 452.250 708.750 453.150 ;
        RECT 709.950 451.950 712.050 454.050 ;
        RECT 713.250 452.250 715.050 453.150 ;
        RECT 706.950 450.450 709.050 451.050 ;
        RECT 704.400 449.400 709.050 450.450 ;
        RECT 710.250 449.850 711.750 450.750 ;
        RECT 706.950 448.950 709.050 449.400 ;
        RECT 712.950 448.950 715.050 451.050 ;
        RECT 700.950 406.950 703.050 409.050 ;
        RECT 713.400 394.050 714.450 448.950 ;
        RECT 703.950 391.950 706.050 394.050 ;
        RECT 712.950 391.950 715.050 394.050 ;
        RECT 697.950 388.950 700.050 391.050 ;
        RECT 691.950 385.950 694.050 388.050 ;
        RECT 691.950 383.850 694.050 384.750 ;
        RECT 694.950 383.250 697.050 384.150 ;
        RECT 694.950 379.950 697.050 382.050 ;
        RECT 695.400 379.050 696.450 379.950 ;
        RECT 694.950 376.950 697.050 379.050 ;
        RECT 704.400 313.050 705.450 391.950 ;
        RECT 712.950 388.950 715.050 391.050 ;
        RECT 706.950 346.950 709.050 349.050 ;
        RECT 707.400 346.050 708.450 346.950 ;
        RECT 713.400 346.050 714.450 388.950 ;
        RECT 706.950 343.950 709.050 346.050 ;
        RECT 710.250 344.250 711.750 345.150 ;
        RECT 712.950 343.950 715.050 346.050 ;
        RECT 716.400 343.050 717.450 523.950 ;
        RECT 734.400 484.050 735.450 526.950 ;
        RECT 740.400 522.450 741.450 703.950 ;
        RECT 748.950 701.850 750.750 702.750 ;
        RECT 751.950 700.950 754.050 703.050 ;
        RECT 755.250 701.850 757.050 702.750 ;
        RECT 748.950 670.950 751.050 673.050 ;
        RECT 748.950 668.850 751.050 669.750 ;
        RECT 742.950 629.250 745.050 630.150 ;
        RECT 748.950 629.250 751.050 630.150 ;
        RECT 742.950 625.950 745.050 628.050 ;
        RECT 743.400 625.050 744.450 625.950 ;
        RECT 742.950 622.950 745.050 625.050 ;
        RECT 742.950 557.250 745.050 558.150 ;
        RECT 748.950 557.250 751.050 558.150 ;
        RECT 742.950 553.950 745.050 556.050 ;
        RECT 742.950 526.950 745.050 529.050 ;
        RECT 742.950 524.850 745.050 525.750 ;
        RECT 748.950 524.850 751.050 525.750 ;
        RECT 740.400 521.400 744.450 522.450 ;
        RECT 739.950 485.250 742.050 486.150 ;
        RECT 733.950 481.950 736.050 484.050 ;
        RECT 739.950 481.950 742.050 484.050 ;
        RECT 740.400 457.050 741.450 481.950 ;
        RECT 743.400 460.050 744.450 521.400 ;
        RECT 745.950 485.250 748.050 486.150 ;
        RECT 752.400 466.050 753.450 700.950 ;
        RECT 754.950 668.850 757.050 669.750 ;
        RECT 751.950 463.950 754.050 466.050 ;
        RECT 758.400 463.050 759.450 704.400 ;
        RECT 760.950 463.950 763.050 466.050 ;
        RECT 745.950 460.950 748.050 463.050 ;
        RECT 757.950 460.950 760.050 463.050 ;
        RECT 742.950 457.950 745.050 460.050 ;
        RECT 739.950 454.950 742.050 457.050 ;
        RECT 733.950 413.250 736.050 414.150 ;
        RECT 739.950 413.250 742.050 414.150 ;
        RECT 739.950 409.950 742.050 412.050 ;
        RECT 736.950 406.950 739.050 409.050 ;
        RECT 730.950 400.950 733.050 403.050 ;
        RECT 724.950 379.950 727.050 382.050 ;
        RECT 706.950 341.850 708.750 342.750 ;
        RECT 709.950 340.950 712.050 343.050 ;
        RECT 713.250 341.850 715.050 342.750 ;
        RECT 715.950 340.950 718.050 343.050 ;
        RECT 703.950 310.950 706.050 313.050 ;
        RECT 704.400 274.050 705.450 310.950 ;
        RECT 725.400 310.050 726.450 379.950 ;
        RECT 731.400 340.050 732.450 400.950 ;
        RECT 737.400 385.050 738.450 406.950 ;
        RECT 740.400 403.050 741.450 409.950 ;
        RECT 739.950 400.950 742.050 403.050 ;
        RECT 743.400 391.050 744.450 457.950 ;
        RECT 742.950 388.950 745.050 391.050 ;
        RECT 743.400 385.050 744.450 388.950 ;
        RECT 736.950 382.950 739.050 385.050 ;
        RECT 740.250 383.250 741.750 384.150 ;
        RECT 742.950 382.950 745.050 385.050 ;
        RECT 733.950 379.950 736.050 382.050 ;
        RECT 737.250 380.850 738.750 381.750 ;
        RECT 739.950 379.950 742.050 382.050 ;
        RECT 743.250 380.850 745.050 381.750 ;
        RECT 740.400 379.050 741.450 379.950 ;
        RECT 733.950 377.850 736.050 378.750 ;
        RECT 739.950 376.950 742.050 379.050 ;
        RECT 736.950 346.950 739.050 349.050 ;
        RECT 730.950 337.950 733.050 340.050 ;
        RECT 721.950 308.250 723.750 309.150 ;
        RECT 724.950 307.950 727.050 310.050 ;
        RECT 728.250 308.250 730.050 309.150 ;
        RECT 721.950 304.950 724.050 307.050 ;
        RECT 725.250 305.850 726.750 306.750 ;
        RECT 727.950 304.950 730.050 307.050 ;
        RECT 712.950 278.400 715.050 280.500 ;
        RECT 697.950 271.950 700.050 274.050 ;
        RECT 701.250 272.250 702.750 273.150 ;
        RECT 703.950 271.950 706.050 274.050 ;
        RECT 706.950 271.950 709.050 274.050 ;
        RECT 697.950 269.850 699.750 270.750 ;
        RECT 700.950 268.950 703.050 271.050 ;
        RECT 704.250 269.850 706.050 270.750 ;
        RECT 707.400 241.050 708.450 271.950 ;
        RECT 713.400 261.600 714.600 278.400 ;
        RECT 718.950 269.250 721.050 270.150 ;
        RECT 718.950 265.950 721.050 268.050 ;
        RECT 712.950 259.500 715.050 261.600 ;
        RECT 719.400 256.050 720.450 265.950 ;
        RECT 712.950 253.950 715.050 256.050 ;
        RECT 718.950 253.950 721.050 256.050 ;
        RECT 713.400 241.050 714.450 253.950 ;
        RECT 722.400 241.050 723.450 304.950 ;
        RECT 733.950 279.300 736.050 281.400 ;
        RECT 734.250 275.700 735.450 279.300 ;
        RECT 733.950 273.600 736.050 275.700 ;
        RECT 724.950 269.250 727.050 270.150 ;
        RECT 724.950 265.950 727.050 268.050 ;
        RECT 706.950 240.450 709.050 241.050 ;
        RECT 704.400 239.400 709.050 240.450 ;
        RECT 704.400 235.050 705.450 239.400 ;
        RECT 706.950 238.950 709.050 239.400 ;
        RECT 710.250 239.250 711.750 240.150 ;
        RECT 712.950 238.950 715.050 241.050 ;
        RECT 721.950 238.950 724.050 241.050 ;
        RECT 706.950 236.850 708.750 237.750 ;
        RECT 709.950 235.950 712.050 238.050 ;
        RECT 713.250 236.850 714.750 237.750 ;
        RECT 715.950 235.950 718.050 238.050 ;
        RECT 703.950 232.950 706.050 235.050 ;
        RECT 704.400 195.450 705.450 232.950 ;
        RECT 710.400 229.050 711.450 235.950 ;
        RECT 715.950 233.850 718.050 234.750 ;
        RECT 709.950 226.950 712.050 229.050 ;
        RECT 715.950 200.250 718.050 201.150 ;
        RECT 706.950 197.250 708.750 198.150 ;
        RECT 709.950 196.950 712.050 199.050 ;
        RECT 713.250 197.250 714.750 198.150 ;
        RECT 715.950 196.950 718.050 199.050 ;
        RECT 706.950 195.450 709.050 196.050 ;
        RECT 704.400 194.400 709.050 195.450 ;
        RECT 710.250 194.850 711.750 195.750 ;
        RECT 706.950 193.950 709.050 194.400 ;
        RECT 712.950 193.950 715.050 196.050 ;
        RECT 707.400 169.050 708.450 193.950 ;
        RECT 716.400 187.050 717.450 196.950 ;
        RECT 725.400 193.050 726.450 265.950 ;
        RECT 734.250 261.600 735.450 273.600 ;
        RECT 737.400 268.050 738.450 346.950 ;
        RECT 746.400 346.050 747.450 460.950 ;
        RECT 757.950 457.950 760.050 460.050 ;
        RECT 758.400 457.050 759.450 457.950 ;
        RECT 751.950 454.950 754.050 457.050 ;
        RECT 755.250 455.250 756.750 456.150 ;
        RECT 757.950 454.950 760.050 457.050 ;
        RECT 748.950 451.950 751.050 454.050 ;
        RECT 752.250 452.850 753.750 453.750 ;
        RECT 754.950 451.950 757.050 454.050 ;
        RECT 758.250 452.850 760.050 453.750 ;
        RECT 755.400 451.050 756.450 451.950 ;
        RECT 748.950 449.850 751.050 450.750 ;
        RECT 754.950 448.950 757.050 451.050 ;
        RECT 742.950 343.950 745.050 346.050 ;
        RECT 745.950 343.950 748.050 346.050 ;
        RECT 754.950 344.250 757.050 345.150 ;
        RECT 757.950 343.950 760.050 346.050 ;
        RECT 739.950 340.950 742.050 343.050 ;
        RECT 740.400 337.050 741.450 340.950 ;
        RECT 743.400 339.450 744.450 343.950 ;
        RECT 745.950 341.250 747.750 342.150 ;
        RECT 748.950 340.950 751.050 343.050 ;
        RECT 752.250 341.250 753.750 342.150 ;
        RECT 754.950 340.950 757.050 343.050 ;
        RECT 745.950 339.450 748.050 340.050 ;
        RECT 743.400 338.400 748.050 339.450 ;
        RECT 749.250 338.850 750.750 339.750 ;
        RECT 739.950 334.950 742.050 337.050 ;
        RECT 743.400 307.050 744.450 338.400 ;
        RECT 745.950 337.950 748.050 338.400 ;
        RECT 751.950 337.950 754.050 340.050 ;
        RECT 742.950 304.950 745.050 307.050 ;
        RECT 736.950 265.950 739.050 268.050 ;
        RECT 745.950 265.950 748.050 268.050 ;
        RECT 736.950 263.850 739.050 264.750 ;
        RECT 733.950 259.500 736.050 261.600 ;
        RECT 746.400 234.450 747.450 265.950 ;
        RECT 748.950 236.250 750.750 237.150 ;
        RECT 751.950 235.950 754.050 238.050 ;
        RECT 755.250 236.250 757.050 237.150 ;
        RECT 748.950 234.450 751.050 235.050 ;
        RECT 746.400 233.400 751.050 234.450 ;
        RECT 752.250 233.850 753.750 234.750 ;
        RECT 748.950 232.950 751.050 233.400 ;
        RECT 754.950 232.950 757.050 235.050 ;
        RECT 727.950 206.400 730.050 208.500 ;
        RECT 748.950 207.300 751.050 209.400 ;
        RECT 724.950 190.950 727.050 193.050 ;
        RECT 728.400 189.600 729.600 206.400 ;
        RECT 749.250 203.700 750.450 207.300 ;
        RECT 748.950 201.600 751.050 203.700 ;
        RECT 733.950 197.250 736.050 198.150 ;
        RECT 739.950 197.250 742.050 198.150 ;
        RECT 733.950 193.950 736.050 196.050 ;
        RECT 739.950 193.950 742.050 196.050 ;
        RECT 740.400 193.050 741.450 193.950 ;
        RECT 739.950 190.950 742.050 193.050 ;
        RECT 749.250 189.600 750.450 201.600 ;
        RECT 758.400 196.050 759.450 343.950 ;
        RECT 761.400 343.050 762.450 463.950 ;
        RECT 760.950 340.950 763.050 343.050 ;
        RECT 751.950 193.950 754.050 196.050 ;
        RECT 757.950 193.950 760.050 196.050 ;
        RECT 751.950 191.850 754.050 192.750 ;
        RECT 727.950 187.500 730.050 189.600 ;
        RECT 748.950 187.500 751.050 189.600 ;
        RECT 715.950 184.950 718.050 187.050 ;
        RECT 751.950 184.950 754.050 187.050 ;
        RECT 706.950 166.950 709.050 169.050 ;
        RECT 712.950 166.950 715.050 169.050 ;
        RECT 703.950 164.250 705.750 165.150 ;
        RECT 706.950 163.950 709.050 166.050 ;
        RECT 710.250 164.250 712.050 165.150 ;
        RECT 713.400 163.050 714.450 166.950 ;
        RECT 752.400 166.050 753.450 184.950 ;
        RECT 748.950 164.250 750.750 165.150 ;
        RECT 751.950 163.950 754.050 166.050 ;
        RECT 755.250 164.250 757.050 165.150 ;
        RECT 703.950 160.950 706.050 163.050 ;
        RECT 707.250 161.850 708.750 162.750 ;
        RECT 709.950 162.450 712.050 163.050 ;
        RECT 712.950 162.450 715.050 163.050 ;
        RECT 709.950 161.400 715.050 162.450 ;
        RECT 709.950 160.950 712.050 161.400 ;
        RECT 712.950 160.950 715.050 161.400 ;
        RECT 748.950 160.950 751.050 163.050 ;
        RECT 752.250 161.850 753.750 162.750 ;
        RECT 754.950 162.450 757.050 163.050 ;
        RECT 758.400 162.450 759.450 193.950 ;
        RECT 754.950 161.400 759.450 162.450 ;
        RECT 754.950 160.950 757.050 161.400 ;
        RECT 718.950 129.450 721.050 130.050 ;
        RECT 716.400 128.400 721.050 129.450 ;
        RECT 670.950 124.950 673.050 127.050 ;
        RECT 673.950 125.850 675.750 126.750 ;
        RECT 676.950 124.950 679.050 127.050 ;
        RECT 680.250 125.850 682.050 126.750 ;
        RECT 688.950 124.950 691.050 127.050 ;
        RECT 677.400 124.050 678.450 124.950 ;
        RECT 676.950 121.950 679.050 124.050 ;
        RECT 716.400 123.450 717.450 128.400 ;
        RECT 718.950 127.950 721.050 128.400 ;
        RECT 722.250 128.250 723.750 129.150 ;
        RECT 724.950 127.950 727.050 130.050 ;
        RECT 745.950 127.950 748.050 130.050 ;
        RECT 718.950 125.850 720.750 126.750 ;
        RECT 721.950 124.950 724.050 127.050 ;
        RECT 725.250 125.850 727.050 126.750 ;
        RECT 716.400 122.400 720.450 123.450 ;
        RECT 661.950 100.950 664.050 103.050 ;
        RECT 643.950 95.250 646.050 96.150 ;
        RECT 662.400 93.450 663.450 100.950 ;
        RECT 700.950 97.950 703.050 100.050 ;
        RECT 709.950 97.950 712.050 100.050 ;
        RECT 664.950 95.250 667.050 96.150 ;
        RECT 700.950 95.850 703.050 96.750 ;
        RECT 703.950 95.250 706.050 96.150 ;
        RECT 664.950 93.450 667.050 94.050 ;
        RECT 662.400 92.400 667.050 93.450 ;
        RECT 664.950 91.950 667.050 92.400 ;
        RECT 703.950 91.950 706.050 94.050 ;
        RECT 607.950 89.400 612.450 90.450 ;
        RECT 607.950 88.950 610.050 89.400 ;
        RECT 613.950 88.950 616.050 91.050 ;
        RECT 514.950 76.950 517.050 79.050 ;
        RECT 586.950 76.950 589.050 79.050 ;
        RECT 469.950 62.400 472.050 64.500 ;
        RECT 463.950 53.250 466.050 54.150 ;
        RECT 457.950 50.400 462.450 51.450 ;
        RECT 457.950 49.950 460.050 50.400 ;
        RECT 463.950 49.950 466.050 52.050 ;
        RECT 458.400 46.050 459.450 49.950 ;
        RECT 464.400 46.050 465.450 49.950 ;
        RECT 433.950 43.500 436.050 45.600 ;
        RECT 448.950 43.500 451.050 45.600 ;
        RECT 457.950 43.950 460.050 46.050 ;
        RECT 463.950 43.950 466.050 46.050 ;
        RECT 470.400 45.600 471.600 62.400 ;
        RECT 511.950 54.450 514.050 55.050 ;
        RECT 515.400 54.450 516.450 76.950 ;
        RECT 610.950 62.400 613.050 64.500 ;
        RECT 547.950 55.950 550.050 58.050 ;
        RECT 550.950 55.950 553.050 58.050 ;
        RECT 554.250 56.250 555.750 57.150 ;
        RECT 592.950 56.250 595.050 57.150 ;
        RECT 598.950 55.950 601.050 58.050 ;
        RECT 511.950 53.400 516.450 54.450 ;
        RECT 511.950 52.950 514.050 53.400 ;
        RECT 508.950 50.250 511.050 51.150 ;
        RECT 511.950 50.850 514.050 51.750 ;
        RECT 508.950 46.950 511.050 49.050 ;
        RECT 469.950 43.500 472.050 45.600 ;
        RECT 508.950 43.950 511.050 46.050 ;
        RECT 509.400 25.050 510.450 43.950 ;
        RECT 515.400 25.050 516.450 53.400 ;
        RECT 421.950 22.950 424.050 25.050 ;
        RECT 425.250 23.250 426.750 24.150 ;
        RECT 427.950 22.950 430.050 25.050 ;
        RECT 508.950 22.950 511.050 25.050 ;
        RECT 512.250 23.250 513.750 24.150 ;
        RECT 514.950 22.950 517.050 25.050 ;
        RECT 379.950 20.250 381.750 21.150 ;
        RECT 382.950 19.950 385.050 22.050 ;
        RECT 386.250 20.250 388.050 21.150 ;
        RECT 418.950 19.950 421.050 22.050 ;
        RECT 422.250 20.850 423.750 21.750 ;
        RECT 424.950 19.950 427.050 22.050 ;
        RECT 428.250 20.850 430.050 21.750 ;
        RECT 463.950 20.250 465.750 21.150 ;
        RECT 466.950 19.950 469.050 22.050 ;
        RECT 470.250 20.250 472.050 21.150 ;
        RECT 505.950 19.950 508.050 22.050 ;
        RECT 509.250 20.850 510.750 21.750 ;
        RECT 511.950 19.950 514.050 22.050 ;
        RECT 515.250 20.850 517.050 21.750 ;
        RECT 425.400 19.050 426.450 19.950 ;
        RECT 512.400 19.050 513.450 19.950 ;
        RECT 379.950 18.450 382.050 19.050 ;
        RECT 377.400 17.400 382.050 18.450 ;
        RECT 383.250 17.850 384.750 18.750 ;
        RECT 418.950 17.850 421.050 18.750 ;
        RECT 379.950 16.950 382.050 17.400 ;
        RECT 424.950 16.950 427.050 19.050 ;
        RECT 463.950 16.950 466.050 19.050 ;
        RECT 467.250 17.850 468.750 18.750 ;
        RECT 505.950 17.850 508.050 18.750 ;
        RECT 511.950 16.950 514.050 19.050 ;
        RECT 548.400 18.450 549.450 55.950 ;
        RECT 599.400 55.050 600.450 55.950 ;
        RECT 550.950 53.850 552.750 54.750 ;
        RECT 553.950 52.950 556.050 55.050 ;
        RECT 557.250 53.850 559.050 54.750 ;
        RECT 592.950 52.950 595.050 55.050 ;
        RECT 596.250 53.250 597.750 54.150 ;
        RECT 598.950 52.950 601.050 55.050 ;
        RECT 602.250 53.250 604.050 54.150 ;
        RECT 595.950 49.950 598.050 52.050 ;
        RECT 599.250 50.850 600.750 51.750 ;
        RECT 601.950 49.950 604.050 52.050 ;
        RECT 596.400 49.050 597.450 49.950 ;
        RECT 595.950 46.950 598.050 49.050 ;
        RECT 611.400 45.600 612.600 62.400 ;
        RECT 614.400 52.050 615.450 88.950 ;
        RECT 631.950 63.300 634.050 65.400 ;
        RECT 632.250 59.700 633.450 63.300 ;
        RECT 631.950 57.600 634.050 59.700 ;
        RECT 634.950 58.950 637.050 61.050 ;
        RECT 616.950 53.250 619.050 54.150 ;
        RECT 622.950 53.250 625.050 54.150 ;
        RECT 613.950 49.950 616.050 52.050 ;
        RECT 616.950 49.950 619.050 52.050 ;
        RECT 622.950 49.950 625.050 52.050 ;
        RECT 617.400 49.050 618.450 49.950 ;
        RECT 616.950 46.950 619.050 49.050 ;
        RECT 610.950 43.500 613.050 45.600 ;
        RECT 610.950 29.400 613.050 31.500 ;
        RECT 595.950 22.950 598.050 25.050 ;
        RECT 601.950 24.450 604.050 25.050 ;
        RECT 599.250 23.250 600.750 24.150 ;
        RECT 601.950 23.400 606.450 24.450 ;
        RECT 601.950 22.950 604.050 23.400 ;
        RECT 605.400 22.050 606.450 23.400 ;
        RECT 550.950 20.250 552.750 21.150 ;
        RECT 553.950 19.950 556.050 22.050 ;
        RECT 557.250 20.250 559.050 21.150 ;
        RECT 592.950 19.950 595.050 22.050 ;
        RECT 596.250 20.850 597.750 21.750 ;
        RECT 598.950 19.950 601.050 22.050 ;
        RECT 602.250 20.850 604.050 21.750 ;
        RECT 604.950 19.950 607.050 22.050 ;
        RECT 599.400 19.050 600.450 19.950 ;
        RECT 550.950 18.450 553.050 19.050 ;
        RECT 548.400 17.400 553.050 18.450 ;
        RECT 554.250 17.850 555.750 18.750 ;
        RECT 592.950 17.850 595.050 18.750 ;
        RECT 550.950 16.950 553.050 17.400 ;
        RECT 598.950 16.950 601.050 19.050 ;
        RECT 181.950 9.600 184.050 11.700 ;
        RECT 196.950 9.600 199.050 11.700 ;
        RECT 217.950 10.500 220.050 12.600 ;
        RECT 316.950 10.500 319.050 12.600 ;
        RECT 338.250 11.700 339.450 15.300 ;
        RECT 611.400 12.600 612.600 29.400 ;
        RECT 623.400 25.050 624.450 49.950 ;
        RECT 632.250 45.600 633.450 57.600 ;
        RECT 635.400 52.050 636.450 58.950 ;
        RECT 665.400 52.050 666.450 91.950 ;
        RECT 704.400 91.050 705.450 91.950 ;
        RECT 703.950 88.950 706.050 91.050 ;
        RECT 710.400 61.050 711.450 97.950 ;
        RECT 709.950 58.950 712.050 61.050 ;
        RECT 710.400 58.050 711.450 58.950 ;
        RECT 670.950 57.450 673.050 58.050 ;
        RECT 668.400 56.400 673.050 57.450 ;
        RECT 634.950 49.950 637.050 52.050 ;
        RECT 664.950 49.950 667.050 52.050 ;
        RECT 668.400 51.450 669.450 56.400 ;
        RECT 670.950 55.950 673.050 56.400 ;
        RECT 674.250 56.250 675.750 57.150 ;
        RECT 676.950 55.950 679.050 58.050 ;
        RECT 709.950 55.950 712.050 58.050 ;
        RECT 713.250 56.250 714.750 57.150 ;
        RECT 715.950 55.950 718.050 58.050 ;
        RECT 719.400 55.050 720.450 122.400 ;
        RECT 746.400 94.050 747.450 127.950 ;
        RECT 742.950 92.250 744.750 93.150 ;
        RECT 745.950 91.950 748.050 94.050 ;
        RECT 749.250 92.250 751.050 93.150 ;
        RECT 742.950 88.950 745.050 91.050 ;
        RECT 746.250 89.850 747.750 90.750 ;
        RECT 754.950 55.950 757.050 58.050 ;
        RECT 755.400 55.050 756.450 55.950 ;
        RECT 670.950 53.850 672.750 54.750 ;
        RECT 673.950 52.950 676.050 55.050 ;
        RECT 677.250 53.850 679.050 54.750 ;
        RECT 709.950 53.850 711.750 54.750 ;
        RECT 712.950 52.950 715.050 55.050 ;
        RECT 716.250 53.850 718.050 54.750 ;
        RECT 718.950 52.950 721.050 55.050 ;
        RECT 754.950 52.950 757.050 55.050 ;
        RECT 668.400 50.400 672.450 51.450 ;
        RECT 634.950 47.850 637.050 48.750 ;
        RECT 631.950 43.500 634.050 45.600 ;
        RECT 631.950 29.400 634.050 31.500 ;
        RECT 616.950 22.950 619.050 25.050 ;
        RECT 622.950 22.950 625.050 25.050 ;
        RECT 616.950 20.850 619.050 21.750 ;
        RECT 622.950 20.850 625.050 21.750 ;
        RECT 632.250 17.400 633.450 29.400 ;
        RECT 634.950 26.250 637.050 27.150 ;
        RECT 668.400 25.050 669.450 50.400 ;
        RECT 671.400 28.050 672.450 50.400 ;
        RECT 670.950 25.950 673.050 28.050 ;
        RECT 674.400 27.450 675.450 52.950 ;
        RECT 751.950 50.250 754.050 51.150 ;
        RECT 754.950 50.850 757.050 51.750 ;
        RECT 715.950 37.950 718.050 40.050 ;
        RECT 674.400 26.400 678.450 27.450 ;
        RECT 634.950 22.950 637.050 25.050 ;
        RECT 667.950 22.950 670.050 25.050 ;
        RECT 670.950 23.850 673.050 24.750 ;
        RECT 673.950 23.250 676.050 24.150 ;
        RECT 673.950 19.950 676.050 22.050 ;
        RECT 677.400 19.050 678.450 26.400 ;
        RECT 716.400 22.050 717.450 37.950 ;
        RECT 712.950 20.250 714.750 21.150 ;
        RECT 715.950 19.950 718.050 22.050 ;
        RECT 719.250 20.250 721.050 21.150 ;
        RECT 721.950 19.950 724.050 22.050 ;
        RECT 748.950 20.250 750.750 21.150 ;
        RECT 751.950 19.950 754.050 22.050 ;
        RECT 755.250 20.250 757.050 21.150 ;
        RECT 631.950 15.300 634.050 17.400 ;
        RECT 676.950 16.950 679.050 19.050 ;
        RECT 712.950 16.950 715.050 19.050 ;
        RECT 716.250 17.850 717.750 18.750 ;
        RECT 718.950 18.450 721.050 19.050 ;
        RECT 722.400 18.450 723.450 19.950 ;
        RECT 718.950 17.400 723.450 18.450 ;
        RECT 752.250 17.850 753.750 18.750 ;
        RECT 718.950 16.950 721.050 17.400 ;
        RECT 754.950 16.950 757.050 19.050 ;
        RECT 337.950 9.600 340.050 11.700 ;
        RECT 610.950 10.500 613.050 12.600 ;
        RECT 632.250 11.700 633.450 15.300 ;
        RECT 631.950 9.600 634.050 11.700 ;
      LAYER metal3 ;
        RECT 103.950 747.600 106.050 748.050 ;
        RECT 181.950 747.600 184.050 748.050 ;
        RECT 103.950 746.400 184.050 747.600 ;
        RECT 103.950 745.950 106.050 746.400 ;
        RECT 181.950 745.950 184.050 746.400 ;
        RECT 196.950 747.600 199.050 748.050 ;
        RECT 229.950 747.600 232.050 748.050 ;
        RECT 196.950 746.400 232.050 747.600 ;
        RECT 196.950 745.950 199.050 746.400 ;
        RECT 229.950 745.950 232.050 746.400 ;
        RECT 268.950 747.600 271.050 748.050 ;
        RECT 283.950 747.600 286.050 748.050 ;
        RECT 268.950 746.400 286.050 747.600 ;
        RECT 268.950 745.950 271.050 746.400 ;
        RECT 283.950 745.950 286.050 746.400 ;
        RECT 562.950 747.600 565.050 748.050 ;
        RECT 595.950 747.600 598.050 748.050 ;
        RECT 634.950 747.600 637.050 748.050 ;
        RECT 562.950 746.400 598.050 747.600 ;
        RECT 562.950 745.950 565.050 746.400 ;
        RECT 595.950 745.950 598.050 746.400 ;
        RECT 599.400 746.400 637.050 747.600 ;
        RECT 76.950 744.600 79.050 745.050 ;
        RECT 97.950 744.600 100.050 745.050 ;
        RECT 76.950 743.400 100.050 744.600 ;
        RECT 76.950 742.950 79.050 743.400 ;
        RECT 97.950 742.950 100.050 743.400 ;
        RECT 154.950 744.600 157.050 745.050 ;
        RECT 175.950 744.600 178.050 745.050 ;
        RECT 154.950 743.400 178.050 744.600 ;
        RECT 154.950 742.950 157.050 743.400 ;
        RECT 175.950 742.950 178.050 743.400 ;
        RECT 271.950 744.600 274.050 745.050 ;
        RECT 292.950 744.600 295.050 745.050 ;
        RECT 271.950 743.400 295.050 744.600 ;
        RECT 271.950 742.950 274.050 743.400 ;
        RECT 292.950 742.950 295.050 743.400 ;
        RECT 391.950 744.600 394.050 745.050 ;
        RECT 397.950 744.600 400.050 745.050 ;
        RECT 391.950 743.400 400.050 744.600 ;
        RECT 391.950 742.950 394.050 743.400 ;
        RECT 397.950 742.950 400.050 743.400 ;
        RECT 403.950 744.600 406.050 745.050 ;
        RECT 463.950 744.600 466.050 745.050 ;
        RECT 403.950 743.400 466.050 744.600 ;
        RECT 403.950 742.950 406.050 743.400 ;
        RECT 463.950 742.950 466.050 743.400 ;
        RECT 481.950 744.600 484.050 745.050 ;
        RECT 599.400 744.600 600.600 746.400 ;
        RECT 634.950 745.950 637.050 746.400 ;
        RECT 640.950 747.600 643.050 748.050 ;
        RECT 682.950 747.600 685.050 748.050 ;
        RECT 640.950 746.400 685.050 747.600 ;
        RECT 640.950 745.950 643.050 746.400 ;
        RECT 682.950 745.950 685.050 746.400 ;
        RECT 481.950 743.400 600.600 744.600 ;
        RECT 622.950 744.600 625.050 745.050 ;
        RECT 715.950 744.600 718.050 745.050 ;
        RECT 622.950 743.400 718.050 744.600 ;
        RECT 481.950 742.950 484.050 743.400 ;
        RECT 622.950 742.950 625.050 743.400 ;
        RECT 715.950 742.950 718.050 743.400 ;
        RECT 31.950 741.600 34.050 742.050 ;
        RECT 73.950 741.600 76.050 742.050 ;
        RECT 31.950 740.400 76.050 741.600 ;
        RECT 31.950 739.950 34.050 740.400 ;
        RECT 73.950 739.950 76.050 740.400 ;
        RECT 127.950 741.600 130.050 742.050 ;
        RECT 151.950 741.600 154.050 742.050 ;
        RECT 127.950 740.400 154.050 741.600 ;
        RECT 127.950 739.950 130.050 740.400 ;
        RECT 151.950 739.950 154.050 740.400 ;
        RECT 163.950 741.600 166.050 742.050 ;
        RECT 232.950 741.600 235.050 742.050 ;
        RECT 235.950 741.600 238.050 742.050 ;
        RECT 163.950 740.400 238.050 741.600 ;
        RECT 163.950 739.950 166.050 740.400 ;
        RECT 232.950 739.950 235.050 740.400 ;
        RECT 235.950 739.950 238.050 740.400 ;
        RECT 316.950 741.600 319.050 742.050 ;
        RECT 352.950 741.600 355.050 742.050 ;
        RECT 316.950 740.400 355.050 741.600 ;
        RECT 316.950 739.950 319.050 740.400 ;
        RECT 352.950 739.950 355.050 740.400 ;
        RECT 358.950 741.600 361.050 742.050 ;
        RECT 400.950 741.600 403.050 742.050 ;
        RECT 358.950 740.400 403.050 741.600 ;
        RECT 358.950 739.950 361.050 740.400 ;
        RECT 400.950 739.950 403.050 740.400 ;
        RECT 406.950 741.600 409.050 742.050 ;
        RECT 442.950 741.600 445.050 742.050 ;
        RECT 406.950 740.400 445.050 741.600 ;
        RECT 406.950 739.950 409.050 740.400 ;
        RECT 442.950 739.950 445.050 740.400 ;
        RECT 34.950 738.600 37.050 739.050 ;
        RECT 85.950 738.600 88.050 739.050 ;
        RECT 34.950 737.400 88.050 738.600 ;
        RECT 34.950 736.950 37.050 737.400 ;
        RECT 85.950 736.950 88.050 737.400 ;
        RECT 277.950 738.600 280.050 739.050 ;
        RECT 361.950 738.600 364.050 739.050 ;
        RECT 277.950 737.400 364.050 738.600 ;
        RECT 277.950 736.950 280.050 737.400 ;
        RECT 361.950 736.950 364.050 737.400 ;
        RECT 439.950 738.600 442.050 739.050 ;
        RECT 481.950 738.600 484.050 739.050 ;
        RECT 439.950 737.400 484.050 738.600 ;
        RECT 439.950 736.950 442.050 737.400 ;
        RECT 481.950 736.950 484.050 737.400 ;
        RECT 34.950 735.600 37.050 736.050 ;
        RECT 79.950 735.600 82.050 736.050 ;
        RECT 259.950 735.600 262.050 736.050 ;
        RECT 34.950 734.400 262.050 735.600 ;
        RECT 34.950 733.950 37.050 734.400 ;
        RECT 79.950 733.950 82.050 734.400 ;
        RECT 259.950 733.950 262.050 734.400 ;
        RECT 283.950 732.600 286.050 733.050 ;
        RECT 319.950 732.600 322.050 733.050 ;
        RECT 283.950 731.400 322.050 732.600 ;
        RECT 283.950 730.950 286.050 731.400 ;
        RECT 319.950 730.950 322.050 731.400 ;
        RECT 76.950 708.600 79.050 709.050 ;
        RECT 535.950 708.600 538.050 709.050 ;
        RECT 76.950 707.400 538.050 708.600 ;
        RECT 76.950 706.950 79.050 707.400 ;
        RECT 535.950 706.950 538.050 707.400 ;
        RECT 115.950 705.600 118.050 706.050 ;
        RECT 220.950 705.600 223.050 706.050 ;
        RECT 115.950 704.400 223.050 705.600 ;
        RECT 115.950 703.950 118.050 704.400 ;
        RECT 220.950 703.950 223.050 704.400 ;
        RECT 376.950 705.600 379.050 706.050 ;
        RECT 391.950 705.600 394.050 706.050 ;
        RECT 427.950 705.600 430.050 706.050 ;
        RECT 445.950 705.600 448.050 706.050 ;
        RECT 376.950 704.400 448.050 705.600 ;
        RECT 376.950 703.950 379.050 704.400 ;
        RECT 391.950 703.950 394.050 704.400 ;
        RECT 427.950 703.950 430.050 704.400 ;
        RECT 445.950 703.950 448.050 704.400 ;
        RECT 484.950 705.600 487.050 706.050 ;
        RECT 520.950 705.600 523.050 706.050 ;
        RECT 544.950 705.600 547.050 706.050 ;
        RECT 484.950 704.400 547.050 705.600 ;
        RECT 484.950 703.950 487.050 704.400 ;
        RECT 520.950 703.950 523.050 704.400 ;
        RECT 544.950 703.950 547.050 704.400 ;
        RECT 739.950 705.600 742.050 706.050 ;
        RECT 748.950 705.600 751.050 706.050 ;
        RECT 739.950 704.400 751.050 705.600 ;
        RECT 739.950 703.950 742.050 704.400 ;
        RECT 748.950 703.950 751.050 704.400 ;
        RECT 115.950 702.600 118.050 703.050 ;
        RECT 121.950 702.600 124.050 703.050 ;
        RECT 115.950 701.400 124.050 702.600 ;
        RECT 115.950 700.950 118.050 701.400 ;
        RECT 121.950 700.950 124.050 701.400 ;
        RECT 208.950 702.600 211.050 703.050 ;
        RECT 292.950 702.600 295.050 703.050 ;
        RECT 313.950 702.600 316.050 703.050 ;
        RECT 208.950 701.400 316.050 702.600 ;
        RECT 208.950 700.950 211.050 701.400 ;
        RECT 292.950 700.950 295.050 701.400 ;
        RECT 313.950 700.950 316.050 701.400 ;
        RECT 334.950 702.600 337.050 703.050 ;
        RECT 415.950 702.600 418.050 703.050 ;
        RECT 334.950 701.400 418.050 702.600 ;
        RECT 334.950 700.950 337.050 701.400 ;
        RECT 415.950 700.950 418.050 701.400 ;
        RECT 421.950 700.950 424.050 703.050 ;
        RECT 433.950 702.600 436.050 703.050 ;
        RECT 502.950 702.600 505.050 703.050 ;
        RECT 589.950 702.600 592.050 703.050 ;
        RECT 433.950 701.400 592.050 702.600 ;
        RECT 433.950 700.950 436.050 701.400 ;
        RECT 502.950 700.950 505.050 701.400 ;
        RECT 589.950 700.950 592.050 701.400 ;
        RECT 631.950 702.600 634.050 703.050 ;
        RECT 637.950 702.600 640.050 703.050 ;
        RECT 631.950 701.400 640.050 702.600 ;
        RECT 631.950 700.950 634.050 701.400 ;
        RECT 637.950 700.950 640.050 701.400 ;
        RECT 85.950 699.600 88.050 700.050 ;
        RECT 88.950 699.600 91.050 700.050 ;
        RECT 118.950 699.600 121.050 700.050 ;
        RECT 157.950 699.600 160.050 700.050 ;
        RECT 166.950 699.600 169.050 700.050 ;
        RECT 85.950 698.400 169.050 699.600 ;
        RECT 85.950 697.950 88.050 698.400 ;
        RECT 88.950 697.950 91.050 698.400 ;
        RECT 118.950 697.950 121.050 698.400 ;
        RECT 157.950 697.950 160.050 698.400 ;
        RECT 166.950 697.950 169.050 698.400 ;
        RECT 289.950 699.600 292.050 700.050 ;
        RECT 322.950 699.600 325.050 700.050 ;
        RECT 367.950 699.600 370.050 700.050 ;
        RECT 289.950 698.400 370.050 699.600 ;
        RECT 289.950 697.950 292.050 698.400 ;
        RECT 322.950 697.950 325.050 698.400 ;
        RECT 367.950 697.950 370.050 698.400 ;
        RECT 379.950 699.600 382.050 700.050 ;
        RECT 422.400 699.600 423.600 700.950 ;
        RECT 379.950 698.400 423.600 699.600 ;
        RECT 424.950 699.600 427.050 700.050 ;
        RECT 445.950 699.600 448.050 700.050 ;
        RECT 424.950 698.400 448.050 699.600 ;
        RECT 379.950 697.950 382.050 698.400 ;
        RECT 424.950 697.950 427.050 698.400 ;
        RECT 445.950 697.950 448.050 698.400 ;
        RECT 586.950 699.600 589.050 700.050 ;
        RECT 622.950 699.600 625.050 700.050 ;
        RECT 586.950 698.400 625.050 699.600 ;
        RECT 586.950 697.950 589.050 698.400 ;
        RECT 622.950 697.950 625.050 698.400 ;
        RECT 628.950 699.600 631.050 700.050 ;
        RECT 709.950 699.600 712.050 700.050 ;
        RECT 628.950 698.400 712.050 699.600 ;
        RECT 628.950 697.950 631.050 698.400 ;
        RECT 709.950 697.950 712.050 698.400 ;
        RECT 82.950 696.600 85.050 697.050 ;
        RECT 169.950 696.600 172.050 697.050 ;
        RECT 82.950 695.400 172.050 696.600 ;
        RECT 82.950 694.950 85.050 695.400 ;
        RECT 169.950 694.950 172.050 695.400 ;
        RECT 250.950 696.600 253.050 697.050 ;
        RECT 328.950 696.600 331.050 697.050 ;
        RECT 373.950 696.600 376.050 697.050 ;
        RECT 250.950 695.400 376.050 696.600 ;
        RECT 250.950 694.950 253.050 695.400 ;
        RECT 328.950 694.950 331.050 695.400 ;
        RECT 373.950 694.950 376.050 695.400 ;
        RECT 466.950 696.600 469.050 697.050 ;
        RECT 499.950 696.600 502.050 697.050 ;
        RECT 466.950 695.400 502.050 696.600 ;
        RECT 466.950 694.950 469.050 695.400 ;
        RECT 499.950 694.950 502.050 695.400 ;
        RECT 547.950 696.600 550.050 697.050 ;
        RECT 598.950 696.600 601.050 697.050 ;
        RECT 547.950 695.400 601.050 696.600 ;
        RECT 547.950 694.950 550.050 695.400 ;
        RECT 598.950 694.950 601.050 695.400 ;
        RECT 634.950 696.600 637.050 697.050 ;
        RECT 673.950 696.600 676.050 697.050 ;
        RECT 634.950 695.400 676.050 696.600 ;
        RECT 634.950 694.950 637.050 695.400 ;
        RECT 673.950 694.950 676.050 695.400 ;
        RECT 259.950 693.600 262.050 694.050 ;
        RECT 295.950 693.600 298.050 694.050 ;
        RECT 259.950 692.400 298.050 693.600 ;
        RECT 259.950 691.950 262.050 692.400 ;
        RECT 295.950 691.950 298.050 692.400 ;
        RECT 451.950 693.600 454.050 694.050 ;
        RECT 472.950 693.600 475.050 694.050 ;
        RECT 541.950 693.600 544.050 694.050 ;
        RECT 550.950 693.600 553.050 694.050 ;
        RECT 451.950 692.400 553.050 693.600 ;
        RECT 451.950 691.950 454.050 692.400 ;
        RECT 472.950 691.950 475.050 692.400 ;
        RECT 541.950 691.950 544.050 692.400 ;
        RECT 550.950 691.950 553.050 692.400 ;
        RECT 592.950 693.600 595.050 694.050 ;
        RECT 634.950 693.600 637.050 694.050 ;
        RECT 592.950 692.400 637.050 693.600 ;
        RECT 592.950 691.950 595.050 692.400 ;
        RECT 634.950 691.950 637.050 692.400 ;
        RECT 172.950 690.600 175.050 691.050 ;
        RECT 451.950 690.600 454.050 691.050 ;
        RECT 172.950 689.400 454.050 690.600 ;
        RECT 172.950 688.950 175.050 689.400 ;
        RECT 451.950 688.950 454.050 689.400 ;
        RECT 211.950 681.600 214.050 682.050 ;
        RECT 232.950 681.600 235.050 682.050 ;
        RECT 241.950 681.600 244.050 682.050 ;
        RECT 211.950 680.400 244.050 681.600 ;
        RECT 211.950 679.950 214.050 680.400 ;
        RECT 232.950 679.950 235.050 680.400 ;
        RECT 241.950 679.950 244.050 680.400 ;
        RECT 205.950 678.600 208.050 679.050 ;
        RECT 253.950 678.600 256.050 679.050 ;
        RECT 205.950 677.400 256.050 678.600 ;
        RECT 205.950 676.950 208.050 677.400 ;
        RECT 253.950 676.950 256.050 677.400 ;
        RECT 283.950 678.600 286.050 679.050 ;
        RECT 382.950 678.600 385.050 679.050 ;
        RECT 283.950 677.400 385.050 678.600 ;
        RECT 283.950 676.950 286.050 677.400 ;
        RECT 382.950 676.950 385.050 677.400 ;
        RECT 37.950 675.600 40.050 676.050 ;
        RECT 46.950 675.600 49.050 676.050 ;
        RECT 37.950 674.400 49.050 675.600 ;
        RECT 37.950 673.950 40.050 674.400 ;
        RECT 46.950 673.950 49.050 674.400 ;
        RECT 109.950 675.600 112.050 676.050 ;
        RECT 157.950 675.600 160.050 676.050 ;
        RECT 205.950 675.600 208.050 676.050 ;
        RECT 109.950 674.400 208.050 675.600 ;
        RECT 109.950 673.950 112.050 674.400 ;
        RECT 157.950 673.950 160.050 674.400 ;
        RECT 205.950 673.950 208.050 674.400 ;
        RECT 220.950 675.600 223.050 676.050 ;
        RECT 289.950 675.600 292.050 676.050 ;
        RECT 220.950 674.400 292.050 675.600 ;
        RECT 220.950 673.950 223.050 674.400 ;
        RECT 289.950 673.950 292.050 674.400 ;
        RECT 433.950 675.600 436.050 676.050 ;
        RECT 469.950 675.600 472.050 676.050 ;
        RECT 484.950 675.600 487.050 676.050 ;
        RECT 433.950 674.400 487.050 675.600 ;
        RECT 433.950 673.950 436.050 674.400 ;
        RECT 469.950 673.950 472.050 674.400 ;
        RECT 484.950 673.950 487.050 674.400 ;
        RECT 550.950 675.600 553.050 676.050 ;
        RECT 580.950 675.600 583.050 676.050 ;
        RECT 550.950 674.400 583.050 675.600 ;
        RECT 550.950 673.950 553.050 674.400 ;
        RECT 580.950 673.950 583.050 674.400 ;
        RECT 598.950 675.600 601.050 676.050 ;
        RECT 700.950 675.600 703.050 676.050 ;
        RECT 598.950 674.400 703.050 675.600 ;
        RECT 598.950 673.950 601.050 674.400 ;
        RECT 700.950 673.950 703.050 674.400 ;
        RECT 64.950 672.600 67.050 673.050 ;
        RECT 73.950 672.600 76.050 673.050 ;
        RECT 64.950 671.400 76.050 672.600 ;
        RECT 64.950 670.950 67.050 671.400 ;
        RECT 73.950 670.950 76.050 671.400 ;
        RECT 76.950 672.600 79.050 673.050 ;
        RECT 85.950 672.600 88.050 673.050 ;
        RECT 76.950 671.400 88.050 672.600 ;
        RECT 76.950 670.950 79.050 671.400 ;
        RECT 85.950 670.950 88.050 671.400 ;
        RECT 154.950 672.600 157.050 673.050 ;
        RECT 163.950 672.600 166.050 673.050 ;
        RECT 154.950 671.400 166.050 672.600 ;
        RECT 154.950 670.950 157.050 671.400 ;
        RECT 163.950 670.950 166.050 671.400 ;
        RECT 211.950 672.600 214.050 673.050 ;
        RECT 220.950 672.600 223.050 673.050 ;
        RECT 211.950 671.400 223.050 672.600 ;
        RECT 211.950 670.950 214.050 671.400 ;
        RECT 220.950 670.950 223.050 671.400 ;
        RECT 250.950 672.600 253.050 673.050 ;
        RECT 376.950 672.600 379.050 673.050 ;
        RECT 250.950 671.400 379.050 672.600 ;
        RECT 250.950 670.950 253.050 671.400 ;
        RECT 376.950 670.950 379.050 671.400 ;
        RECT 400.950 672.600 403.050 673.050 ;
        RECT 427.950 672.600 430.050 673.050 ;
        RECT 400.950 671.400 430.050 672.600 ;
        RECT 400.950 670.950 403.050 671.400 ;
        RECT 427.950 670.950 430.050 671.400 ;
        RECT 451.950 672.600 454.050 673.050 ;
        RECT 463.950 672.600 466.050 673.050 ;
        RECT 505.950 672.600 508.050 673.050 ;
        RECT 451.950 671.400 466.050 672.600 ;
        RECT 451.950 670.950 454.050 671.400 ;
        RECT 463.950 670.950 466.050 671.400 ;
        RECT 482.400 671.400 508.050 672.600 ;
        RECT 46.950 669.600 49.050 670.050 ;
        RECT 160.950 669.600 163.050 670.050 ;
        RECT 46.950 668.400 163.050 669.600 ;
        RECT 46.950 667.950 49.050 668.400 ;
        RECT 160.950 667.950 163.050 668.400 ;
        RECT 238.950 669.600 241.050 670.050 ;
        RECT 247.950 669.600 250.050 670.050 ;
        RECT 238.950 668.400 250.050 669.600 ;
        RECT 238.950 667.950 241.050 668.400 ;
        RECT 247.950 667.950 250.050 668.400 ;
        RECT 292.950 669.600 295.050 670.050 ;
        RECT 331.950 669.600 334.050 670.050 ;
        RECT 421.950 669.600 424.050 670.050 ;
        RECT 482.400 669.600 483.600 671.400 ;
        RECT 505.950 670.950 508.050 671.400 ;
        RECT 508.950 672.600 511.050 673.050 ;
        RECT 529.950 672.600 532.050 673.050 ;
        RECT 508.950 671.400 532.050 672.600 ;
        RECT 508.950 670.950 511.050 671.400 ;
        RECT 529.950 670.950 532.050 671.400 ;
        RECT 535.950 672.600 538.050 673.050 ;
        RECT 541.950 672.600 544.050 673.050 ;
        RECT 535.950 671.400 544.050 672.600 ;
        RECT 535.950 670.950 538.050 671.400 ;
        RECT 541.950 670.950 544.050 671.400 ;
        RECT 655.950 672.600 658.050 673.050 ;
        RECT 664.950 672.600 667.050 673.050 ;
        RECT 655.950 671.400 667.050 672.600 ;
        RECT 655.950 670.950 658.050 671.400 ;
        RECT 664.950 670.950 667.050 671.400 ;
        RECT 673.950 672.600 676.050 673.050 ;
        RECT 703.950 672.600 706.050 673.050 ;
        RECT 673.950 671.400 706.050 672.600 ;
        RECT 673.950 670.950 676.050 671.400 ;
        RECT 703.950 670.950 706.050 671.400 ;
        RECT 712.950 672.600 715.050 673.050 ;
        RECT 748.950 672.600 751.050 673.050 ;
        RECT 712.950 671.400 751.050 672.600 ;
        RECT 712.950 670.950 715.050 671.400 ;
        RECT 748.950 670.950 751.050 671.400 ;
        RECT 292.950 668.400 334.050 669.600 ;
        RECT 292.950 667.950 295.050 668.400 ;
        RECT 331.950 667.950 334.050 668.400 ;
        RECT 377.400 668.400 424.050 669.600 ;
        RECT 34.950 666.600 37.050 667.050 ;
        RECT 67.950 666.600 70.050 667.050 ;
        RECT 34.950 665.400 70.050 666.600 ;
        RECT 34.950 664.950 37.050 665.400 ;
        RECT 67.950 664.950 70.050 665.400 ;
        RECT 85.950 666.600 88.050 667.050 ;
        RECT 118.950 666.600 121.050 667.050 ;
        RECT 85.950 665.400 121.050 666.600 ;
        RECT 85.950 664.950 88.050 665.400 ;
        RECT 118.950 664.950 121.050 665.400 ;
        RECT 328.950 666.600 331.050 667.050 ;
        RECT 334.950 666.600 337.050 667.050 ;
        RECT 328.950 665.400 337.050 666.600 ;
        RECT 328.950 664.950 331.050 665.400 ;
        RECT 334.950 664.950 337.050 665.400 ;
        RECT 340.950 666.600 343.050 667.050 ;
        RECT 377.400 666.600 378.600 668.400 ;
        RECT 421.950 667.950 424.050 668.400 ;
        RECT 428.400 668.400 483.600 669.600 ;
        RECT 484.950 669.600 487.050 670.050 ;
        RECT 511.950 669.600 514.050 670.050 ;
        RECT 484.950 668.400 514.050 669.600 ;
        RECT 340.950 665.400 378.600 666.600 ;
        RECT 340.950 664.950 343.050 665.400 ;
        RECT 379.950 664.950 382.050 667.050 ;
        RECT 424.950 666.600 427.050 667.050 ;
        RECT 428.400 666.600 429.600 668.400 ;
        RECT 484.950 667.950 487.050 668.400 ;
        RECT 511.950 667.950 514.050 668.400 ;
        RECT 517.950 669.600 520.050 670.050 ;
        RECT 583.950 669.600 586.050 670.050 ;
        RECT 670.950 669.600 673.050 670.050 ;
        RECT 517.950 668.400 673.050 669.600 ;
        RECT 517.950 667.950 520.050 668.400 ;
        RECT 583.950 667.950 586.050 668.400 ;
        RECT 670.950 667.950 673.050 668.400 ;
        RECT 700.950 669.600 703.050 670.050 ;
        RECT 709.950 669.600 712.050 670.050 ;
        RECT 700.950 668.400 712.050 669.600 ;
        RECT 700.950 667.950 703.050 668.400 ;
        RECT 709.950 667.950 712.050 668.400 ;
        RECT 424.950 665.400 429.600 666.600 ;
        RECT 424.950 664.950 427.050 665.400 ;
        RECT 430.950 664.950 433.050 667.050 ;
        RECT 628.950 666.600 631.050 667.050 ;
        RECT 634.950 666.600 637.050 667.050 ;
        RECT 628.950 665.400 637.050 666.600 ;
        RECT 628.950 664.950 631.050 665.400 ;
        RECT 634.950 664.950 637.050 665.400 ;
        RECT 115.950 663.600 118.050 664.050 ;
        RECT 121.950 663.600 124.050 664.050 ;
        RECT 115.950 662.400 124.050 663.600 ;
        RECT 115.950 661.950 118.050 662.400 ;
        RECT 121.950 661.950 124.050 662.400 ;
        RECT 346.950 663.600 349.050 664.050 ;
        RECT 380.400 663.600 381.600 664.950 ;
        RECT 403.950 663.600 406.050 664.050 ;
        RECT 346.950 662.400 406.050 663.600 ;
        RECT 346.950 661.950 349.050 662.400 ;
        RECT 403.950 661.950 406.050 662.400 ;
        RECT 421.950 663.600 424.050 664.050 ;
        RECT 431.400 663.600 432.600 664.950 ;
        RECT 421.950 662.400 432.600 663.600 ;
        RECT 421.950 661.950 424.050 662.400 ;
        RECT 484.950 648.600 487.050 649.050 ;
        RECT 622.950 648.600 625.050 649.050 ;
        RECT 484.950 647.400 625.050 648.600 ;
        RECT 484.950 646.950 487.050 647.400 ;
        RECT 622.950 646.950 625.050 647.400 ;
        RECT 235.950 639.600 238.050 640.050 ;
        RECT 664.950 639.600 667.050 640.050 ;
        RECT 235.950 638.400 667.050 639.600 ;
        RECT 235.950 637.950 238.050 638.400 ;
        RECT 664.950 637.950 667.050 638.400 ;
        RECT 37.950 636.600 40.050 637.050 ;
        RECT 43.950 636.600 46.050 637.050 ;
        RECT 79.950 636.600 82.050 637.050 ;
        RECT 109.950 636.600 112.050 637.050 ;
        RECT 37.950 635.400 112.050 636.600 ;
        RECT 37.950 634.950 40.050 635.400 ;
        RECT 43.950 634.950 46.050 635.400 ;
        RECT 79.950 634.950 82.050 635.400 ;
        RECT 109.950 634.950 112.050 635.400 ;
        RECT 169.950 636.600 172.050 637.050 ;
        RECT 208.950 636.600 211.050 637.050 ;
        RECT 169.950 635.400 211.050 636.600 ;
        RECT 169.950 634.950 172.050 635.400 ;
        RECT 208.950 634.950 211.050 635.400 ;
        RECT 286.950 636.600 289.050 637.050 ;
        RECT 295.950 636.600 298.050 637.050 ;
        RECT 310.950 636.600 313.050 637.050 ;
        RECT 286.950 635.400 313.050 636.600 ;
        RECT 286.950 634.950 289.050 635.400 ;
        RECT 295.950 634.950 298.050 635.400 ;
        RECT 310.950 634.950 313.050 635.400 ;
        RECT 364.950 636.600 367.050 637.050 ;
        RECT 373.950 636.600 376.050 637.050 ;
        RECT 364.950 635.400 376.050 636.600 ;
        RECT 364.950 634.950 367.050 635.400 ;
        RECT 373.950 634.950 376.050 635.400 ;
        RECT 385.950 636.600 388.050 637.050 ;
        RECT 490.950 636.600 493.050 637.050 ;
        RECT 385.950 635.400 493.050 636.600 ;
        RECT 385.950 634.950 388.050 635.400 ;
        RECT 490.950 634.950 493.050 635.400 ;
        RECT 538.950 636.600 541.050 637.050 ;
        RECT 577.950 636.600 580.050 637.050 ;
        RECT 538.950 635.400 580.050 636.600 ;
        RECT 538.950 634.950 541.050 635.400 ;
        RECT 577.950 634.950 580.050 635.400 ;
        RECT 31.950 633.600 34.050 634.050 ;
        RECT 40.950 633.600 43.050 634.050 ;
        RECT 31.950 632.400 43.050 633.600 ;
        RECT 31.950 631.950 34.050 632.400 ;
        RECT 40.950 631.950 43.050 632.400 ;
        RECT 73.950 633.600 76.050 634.050 ;
        RECT 151.950 633.600 154.050 634.050 ;
        RECT 160.950 633.600 163.050 634.050 ;
        RECT 73.950 632.400 96.600 633.600 ;
        RECT 73.950 631.950 76.050 632.400 ;
        RECT 34.950 630.600 37.050 631.050 ;
        RECT 64.950 630.600 67.050 631.050 ;
        RECT 34.950 629.400 67.050 630.600 ;
        RECT 34.950 628.950 37.050 629.400 ;
        RECT 64.950 628.950 67.050 629.400 ;
        RECT 76.950 630.600 79.050 631.050 ;
        RECT 85.950 630.600 88.050 631.050 ;
        RECT 76.950 629.400 88.050 630.600 ;
        RECT 95.400 630.600 96.600 632.400 ;
        RECT 151.950 632.400 163.050 633.600 ;
        RECT 151.950 631.950 154.050 632.400 ;
        RECT 160.950 631.950 163.050 632.400 ;
        RECT 190.950 633.600 193.050 634.050 ;
        RECT 202.950 633.600 205.050 634.050 ;
        RECT 190.950 632.400 205.050 633.600 ;
        RECT 190.950 631.950 193.050 632.400 ;
        RECT 202.950 631.950 205.050 632.400 ;
        RECT 292.950 633.600 295.050 634.050 ;
        RECT 316.950 633.600 319.050 634.050 ;
        RECT 322.950 633.600 325.050 634.050 ;
        RECT 292.950 632.400 325.050 633.600 ;
        RECT 292.950 631.950 295.050 632.400 ;
        RECT 316.950 631.950 319.050 632.400 ;
        RECT 322.950 631.950 325.050 632.400 ;
        RECT 361.950 633.600 364.050 634.050 ;
        RECT 367.950 633.600 370.050 634.050 ;
        RECT 361.950 632.400 370.050 633.600 ;
        RECT 361.950 631.950 364.050 632.400 ;
        RECT 367.950 631.950 370.050 632.400 ;
        RECT 403.950 633.600 406.050 634.050 ;
        RECT 415.950 633.600 418.050 634.050 ;
        RECT 403.950 632.400 418.050 633.600 ;
        RECT 403.950 631.950 406.050 632.400 ;
        RECT 415.950 631.950 418.050 632.400 ;
        RECT 523.950 633.600 526.050 634.050 ;
        RECT 583.950 633.600 586.050 634.050 ;
        RECT 523.950 632.400 586.050 633.600 ;
        RECT 523.950 631.950 526.050 632.400 ;
        RECT 583.950 631.950 586.050 632.400 ;
        RECT 622.950 633.600 625.050 634.050 ;
        RECT 628.950 633.600 631.050 634.050 ;
        RECT 622.950 632.400 631.050 633.600 ;
        RECT 622.950 631.950 625.050 632.400 ;
        RECT 628.950 631.950 631.050 632.400 ;
        RECT 118.950 630.600 121.050 631.050 ;
        RECT 163.950 630.600 166.050 631.050 ;
        RECT 95.400 629.400 166.050 630.600 ;
        RECT 76.950 628.950 79.050 629.400 ;
        RECT 85.950 628.950 88.050 629.400 ;
        RECT 118.950 628.950 121.050 629.400 ;
        RECT 163.950 628.950 166.050 629.400 ;
        RECT 205.950 630.600 208.050 631.050 ;
        RECT 247.950 630.600 250.050 631.050 ;
        RECT 205.950 629.400 250.050 630.600 ;
        RECT 205.950 628.950 208.050 629.400 ;
        RECT 247.950 628.950 250.050 629.400 ;
        RECT 325.950 630.600 328.050 631.050 ;
        RECT 346.950 630.600 349.050 631.050 ;
        RECT 325.950 629.400 349.050 630.600 ;
        RECT 325.950 628.950 328.050 629.400 ;
        RECT 346.950 628.950 349.050 629.400 ;
        RECT 370.950 630.600 373.050 631.050 ;
        RECT 400.950 630.600 403.050 631.050 ;
        RECT 370.950 629.400 403.050 630.600 ;
        RECT 370.950 628.950 373.050 629.400 ;
        RECT 400.950 628.950 403.050 629.400 ;
        RECT 406.950 630.600 409.050 631.050 ;
        RECT 418.950 630.600 421.050 631.050 ;
        RECT 454.950 630.600 457.050 631.050 ;
        RECT 406.950 629.400 417.600 630.600 ;
        RECT 406.950 628.950 409.050 629.400 ;
        RECT 244.950 627.600 247.050 628.050 ;
        RECT 283.950 627.600 286.050 628.050 ;
        RECT 244.950 626.400 286.050 627.600 ;
        RECT 244.950 625.950 247.050 626.400 ;
        RECT 283.950 625.950 286.050 626.400 ;
        RECT 289.950 627.600 292.050 628.050 ;
        RECT 361.950 627.600 364.050 628.050 ;
        RECT 412.950 627.600 415.050 628.050 ;
        RECT 289.950 626.400 415.050 627.600 ;
        RECT 416.400 627.600 417.600 629.400 ;
        RECT 418.950 629.400 457.050 630.600 ;
        RECT 418.950 628.950 421.050 629.400 ;
        RECT 454.950 628.950 457.050 629.400 ;
        RECT 493.950 630.600 496.050 631.050 ;
        RECT 508.950 630.600 511.050 631.050 ;
        RECT 493.950 629.400 511.050 630.600 ;
        RECT 493.950 628.950 496.050 629.400 ;
        RECT 508.950 628.950 511.050 629.400 ;
        RECT 511.950 630.600 514.050 631.050 ;
        RECT 529.950 630.600 532.050 631.050 ;
        RECT 511.950 629.400 532.050 630.600 ;
        RECT 511.950 628.950 514.050 629.400 ;
        RECT 529.950 628.950 532.050 629.400 ;
        RECT 619.950 630.600 622.050 631.050 ;
        RECT 658.950 630.600 661.050 631.050 ;
        RECT 619.950 629.400 661.050 630.600 ;
        RECT 619.950 628.950 622.050 629.400 ;
        RECT 658.950 628.950 661.050 629.400 ;
        RECT 535.950 627.600 538.050 628.050 ;
        RECT 416.400 626.400 538.050 627.600 ;
        RECT 289.950 625.950 292.050 626.400 ;
        RECT 361.950 625.950 364.050 626.400 ;
        RECT 412.950 625.950 415.050 626.400 ;
        RECT 535.950 625.950 538.050 626.400 ;
        RECT 661.950 627.600 664.050 628.050 ;
        RECT 661.950 626.400 690.600 627.600 ;
        RECT 661.950 625.950 664.050 626.400 ;
        RECT 457.950 624.600 460.050 625.050 ;
        RECT 499.950 624.600 502.050 625.050 ;
        RECT 457.950 623.400 502.050 624.600 ;
        RECT 457.950 622.950 460.050 623.400 ;
        RECT 499.950 622.950 502.050 623.400 ;
        RECT 634.950 624.600 637.050 625.050 ;
        RECT 661.950 624.600 664.050 625.050 ;
        RECT 667.950 624.600 670.050 625.050 ;
        RECT 682.950 624.600 685.050 625.050 ;
        RECT 634.950 623.400 685.050 624.600 ;
        RECT 689.400 624.600 690.600 626.400 ;
        RECT 742.950 624.600 745.050 625.050 ;
        RECT 689.400 623.400 745.050 624.600 ;
        RECT 634.950 622.950 637.050 623.400 ;
        RECT 661.950 622.950 664.050 623.400 ;
        RECT 667.950 622.950 670.050 623.400 ;
        RECT 682.950 622.950 685.050 623.400 ;
        RECT 742.950 622.950 745.050 623.400 ;
        RECT 241.950 621.600 244.050 622.050 ;
        RECT 316.950 621.600 319.050 622.050 ;
        RECT 241.950 620.400 319.050 621.600 ;
        RECT 241.950 619.950 244.050 620.400 ;
        RECT 316.950 619.950 319.050 620.400 ;
        RECT 550.950 615.600 553.050 616.050 ;
        RECT 580.950 615.600 583.050 616.050 ;
        RECT 550.950 614.400 583.050 615.600 ;
        RECT 550.950 613.950 553.050 614.400 ;
        RECT 580.950 613.950 583.050 614.400 ;
        RECT 40.950 606.600 43.050 607.050 ;
        RECT 76.950 606.600 79.050 607.050 ;
        RECT 79.950 606.600 82.050 607.050 ;
        RECT 115.950 606.600 118.050 607.050 ;
        RECT 40.950 605.400 118.050 606.600 ;
        RECT 40.950 604.950 43.050 605.400 ;
        RECT 76.950 604.950 79.050 605.400 ;
        RECT 79.950 604.950 82.050 605.400 ;
        RECT 115.950 604.950 118.050 605.400 ;
        RECT 37.950 603.600 40.050 604.050 ;
        RECT 190.950 603.600 193.050 604.050 ;
        RECT 37.950 602.400 193.050 603.600 ;
        RECT 37.950 601.950 40.050 602.400 ;
        RECT 190.950 601.950 193.050 602.400 ;
        RECT 235.950 603.600 238.050 604.050 ;
        RECT 274.950 603.600 277.050 604.050 ;
        RECT 235.950 602.400 277.050 603.600 ;
        RECT 235.950 601.950 238.050 602.400 ;
        RECT 274.950 601.950 277.050 602.400 ;
        RECT 313.950 603.600 316.050 604.050 ;
        RECT 331.950 603.600 334.050 604.050 ;
        RECT 364.950 603.600 367.050 604.050 ;
        RECT 313.950 602.400 367.050 603.600 ;
        RECT 313.950 601.950 316.050 602.400 ;
        RECT 331.950 601.950 334.050 602.400 ;
        RECT 364.950 601.950 367.050 602.400 ;
        RECT 529.950 603.600 532.050 604.050 ;
        RECT 595.950 603.600 598.050 604.050 ;
        RECT 529.950 602.400 598.050 603.600 ;
        RECT 529.950 601.950 532.050 602.400 ;
        RECT 595.950 601.950 598.050 602.400 ;
        RECT 34.950 600.600 37.050 601.050 ;
        RECT 46.950 600.600 49.050 601.050 ;
        RECT 34.950 599.400 49.050 600.600 ;
        RECT 34.950 598.950 37.050 599.400 ;
        RECT 46.950 598.950 49.050 599.400 ;
        RECT 148.950 600.600 151.050 601.050 ;
        RECT 169.950 600.600 172.050 601.050 ;
        RECT 184.950 600.600 187.050 601.050 ;
        RECT 148.950 599.400 187.050 600.600 ;
        RECT 148.950 598.950 151.050 599.400 ;
        RECT 169.950 598.950 172.050 599.400 ;
        RECT 184.950 598.950 187.050 599.400 ;
        RECT 196.950 600.600 199.050 601.050 ;
        RECT 280.950 600.600 283.050 601.050 ;
        RECT 196.950 599.400 283.050 600.600 ;
        RECT 196.950 598.950 199.050 599.400 ;
        RECT 280.950 598.950 283.050 599.400 ;
        RECT 400.950 600.600 403.050 601.050 ;
        RECT 463.950 600.600 466.050 601.050 ;
        RECT 400.950 599.400 466.050 600.600 ;
        RECT 400.950 598.950 403.050 599.400 ;
        RECT 463.950 598.950 466.050 599.400 ;
        RECT 469.950 600.600 472.050 601.050 ;
        RECT 541.950 600.600 544.050 601.050 ;
        RECT 544.950 600.600 547.050 601.050 ;
        RECT 469.950 599.400 547.050 600.600 ;
        RECT 469.950 598.950 472.050 599.400 ;
        RECT 541.950 598.950 544.050 599.400 ;
        RECT 544.950 598.950 547.050 599.400 ;
        RECT 685.950 600.600 688.050 601.050 ;
        RECT 721.950 600.600 724.050 601.050 ;
        RECT 685.950 599.400 724.050 600.600 ;
        RECT 685.950 598.950 688.050 599.400 ;
        RECT 721.950 598.950 724.050 599.400 ;
        RECT 73.950 597.600 76.050 598.050 ;
        RECT 124.950 597.600 127.050 598.050 ;
        RECT 145.950 597.600 148.050 598.050 ;
        RECT 73.950 596.400 148.050 597.600 ;
        RECT 73.950 595.950 76.050 596.400 ;
        RECT 124.950 595.950 127.050 596.400 ;
        RECT 145.950 595.950 148.050 596.400 ;
        RECT 151.950 597.600 154.050 598.050 ;
        RECT 277.950 597.600 280.050 598.050 ;
        RECT 151.950 596.400 280.050 597.600 ;
        RECT 151.950 595.950 154.050 596.400 ;
        RECT 277.950 595.950 280.050 596.400 ;
        RECT 322.950 597.600 325.050 598.050 ;
        RECT 328.950 597.600 331.050 598.050 ;
        RECT 322.950 596.400 331.050 597.600 ;
        RECT 322.950 595.950 325.050 596.400 ;
        RECT 328.950 595.950 331.050 596.400 ;
        RECT 361.950 597.600 364.050 598.050 ;
        RECT 367.950 597.600 370.050 598.050 ;
        RECT 361.950 596.400 370.050 597.600 ;
        RECT 361.950 595.950 364.050 596.400 ;
        RECT 367.950 595.950 370.050 596.400 ;
        RECT 403.950 597.600 406.050 598.050 ;
        RECT 445.950 597.600 448.050 598.050 ;
        RECT 403.950 596.400 448.050 597.600 ;
        RECT 403.950 595.950 406.050 596.400 ;
        RECT 445.950 595.950 448.050 596.400 ;
        RECT 598.950 597.600 601.050 598.050 ;
        RECT 637.950 597.600 640.050 598.050 ;
        RECT 598.950 596.400 640.050 597.600 ;
        RECT 598.950 595.950 601.050 596.400 ;
        RECT 637.950 595.950 640.050 596.400 ;
        RECT 277.950 592.950 280.050 595.050 ;
        RECT 283.950 594.600 286.050 595.050 ;
        RECT 295.950 594.600 298.050 595.050 ;
        RECT 283.950 593.400 298.050 594.600 ;
        RECT 283.950 592.950 286.050 593.400 ;
        RECT 295.950 592.950 298.050 593.400 ;
        RECT 307.950 594.600 310.050 595.050 ;
        RECT 397.950 594.600 400.050 595.050 ;
        RECT 307.950 593.400 400.050 594.600 ;
        RECT 307.950 592.950 310.050 593.400 ;
        RECT 397.950 592.950 400.050 593.400 ;
        RECT 448.950 594.600 451.050 595.050 ;
        RECT 481.950 594.600 484.050 595.050 ;
        RECT 448.950 593.400 484.050 594.600 ;
        RECT 448.950 592.950 451.050 593.400 ;
        RECT 481.950 592.950 484.050 593.400 ;
        RECT 278.400 591.600 279.600 592.950 ;
        RECT 280.950 591.600 283.050 592.050 ;
        RECT 278.400 590.400 283.050 591.600 ;
        RECT 280.950 589.950 283.050 590.400 ;
        RECT 250.950 588.600 253.050 589.050 ;
        RECT 271.950 588.600 274.050 589.050 ;
        RECT 325.950 588.600 328.050 589.050 ;
        RECT 250.950 587.400 328.050 588.600 ;
        RECT 250.950 586.950 253.050 587.400 ;
        RECT 271.950 586.950 274.050 587.400 ;
        RECT 325.950 586.950 328.050 587.400 ;
        RECT 109.950 567.600 112.050 568.050 ;
        RECT 160.950 567.600 163.050 568.050 ;
        RECT 229.950 567.600 232.050 568.050 ;
        RECT 109.950 566.400 232.050 567.600 ;
        RECT 109.950 565.950 112.050 566.400 ;
        RECT 160.950 565.950 163.050 566.400 ;
        RECT 229.950 565.950 232.050 566.400 ;
        RECT 121.950 564.600 124.050 565.050 ;
        RECT 166.950 564.600 169.050 565.050 ;
        RECT 121.950 563.400 169.050 564.600 ;
        RECT 121.950 562.950 124.050 563.400 ;
        RECT 166.950 562.950 169.050 563.400 ;
        RECT 586.950 562.950 589.050 565.050 ;
        RECT 40.950 561.600 43.050 562.050 ;
        RECT 64.950 561.600 67.050 562.050 ;
        RECT 82.950 561.600 85.050 562.050 ;
        RECT 40.950 560.400 85.050 561.600 ;
        RECT 40.950 559.950 43.050 560.400 ;
        RECT 64.950 559.950 67.050 560.400 ;
        RECT 82.950 559.950 85.050 560.400 ;
        RECT 421.950 561.600 424.050 562.050 ;
        RECT 442.950 561.600 445.050 562.050 ;
        RECT 469.950 561.600 472.050 562.050 ;
        RECT 478.950 561.600 481.050 562.050 ;
        RECT 520.950 561.600 523.050 562.050 ;
        RECT 421.950 560.400 523.050 561.600 ;
        RECT 421.950 559.950 424.050 560.400 ;
        RECT 442.950 559.950 445.050 560.400 ;
        RECT 469.950 559.950 472.050 560.400 ;
        RECT 478.950 559.950 481.050 560.400 ;
        RECT 520.950 559.950 523.050 560.400 ;
        RECT 34.950 558.600 37.050 559.050 ;
        RECT 79.950 558.600 82.050 559.050 ;
        RECT 34.950 557.400 82.050 558.600 ;
        RECT 34.950 556.950 37.050 557.400 ;
        RECT 79.950 556.950 82.050 557.400 ;
        RECT 112.950 558.600 115.050 559.050 ;
        RECT 121.950 558.600 124.050 559.050 ;
        RECT 112.950 557.400 124.050 558.600 ;
        RECT 112.950 556.950 115.050 557.400 ;
        RECT 121.950 556.950 124.050 557.400 ;
        RECT 127.950 558.600 130.050 559.050 ;
        RECT 163.950 558.600 166.050 559.050 ;
        RECT 127.950 557.400 166.050 558.600 ;
        RECT 127.950 556.950 130.050 557.400 ;
        RECT 163.950 556.950 166.050 557.400 ;
        RECT 280.950 558.600 283.050 559.050 ;
        RECT 286.950 558.600 289.050 559.050 ;
        RECT 280.950 557.400 289.050 558.600 ;
        RECT 280.950 556.950 283.050 557.400 ;
        RECT 286.950 556.950 289.050 557.400 ;
        RECT 316.950 558.600 319.050 559.050 ;
        RECT 334.950 558.600 337.050 559.050 ;
        RECT 316.950 557.400 337.050 558.600 ;
        RECT 316.950 556.950 319.050 557.400 ;
        RECT 334.950 556.950 337.050 557.400 ;
        RECT 379.950 558.600 382.050 559.050 ;
        RECT 457.950 558.600 460.050 559.050 ;
        RECT 379.950 557.400 460.050 558.600 ;
        RECT 379.950 556.950 382.050 557.400 ;
        RECT 457.950 556.950 460.050 557.400 ;
        RECT 463.950 556.950 466.050 559.050 ;
        RECT 475.950 558.600 478.050 559.050 ;
        RECT 541.950 558.600 544.050 559.050 ;
        RECT 583.950 558.600 586.050 559.050 ;
        RECT 587.400 558.600 588.600 562.950 ;
        RECT 667.950 561.600 670.050 562.050 ;
        RECT 676.950 561.600 679.050 562.050 ;
        RECT 667.950 560.400 679.050 561.600 ;
        RECT 667.950 559.950 670.050 560.400 ;
        RECT 676.950 559.950 679.050 560.400 ;
        RECT 475.950 557.400 582.600 558.600 ;
        RECT 475.950 556.950 478.050 557.400 ;
        RECT 541.950 556.950 544.050 557.400 ;
        RECT 43.950 555.600 46.050 556.050 ;
        RECT 118.950 555.600 121.050 556.050 ;
        RECT 43.950 554.400 121.050 555.600 ;
        RECT 43.950 553.950 46.050 554.400 ;
        RECT 118.950 553.950 121.050 554.400 ;
        RECT 193.950 555.600 196.050 556.050 ;
        RECT 208.950 555.600 211.050 556.050 ;
        RECT 232.950 555.600 235.050 556.050 ;
        RECT 193.950 554.400 235.050 555.600 ;
        RECT 193.950 553.950 196.050 554.400 ;
        RECT 208.950 553.950 211.050 554.400 ;
        RECT 232.950 553.950 235.050 554.400 ;
        RECT 259.950 555.600 262.050 556.050 ;
        RECT 283.950 555.600 286.050 556.050 ;
        RECT 304.950 555.600 307.050 556.050 ;
        RECT 337.950 555.600 340.050 556.050 ;
        RECT 259.950 554.400 340.050 555.600 ;
        RECT 259.950 553.950 262.050 554.400 ;
        RECT 283.950 553.950 286.050 554.400 ;
        RECT 304.950 553.950 307.050 554.400 ;
        RECT 337.950 553.950 340.050 554.400 ;
        RECT 424.950 555.600 427.050 556.050 ;
        RECT 464.400 555.600 465.600 556.950 ;
        RECT 424.950 554.400 465.600 555.600 ;
        RECT 466.950 555.600 469.050 556.050 ;
        RECT 487.950 555.600 490.050 556.050 ;
        RECT 466.950 554.400 490.050 555.600 ;
        RECT 581.400 555.600 582.600 557.400 ;
        RECT 583.950 557.400 588.600 558.600 ;
        RECT 583.950 556.950 586.050 557.400 ;
        RECT 622.950 556.950 625.050 559.050 ;
        RECT 646.950 558.600 649.050 559.050 ;
        RECT 664.950 558.600 667.050 559.050 ;
        RECT 646.950 557.400 667.050 558.600 ;
        RECT 646.950 556.950 649.050 557.400 ;
        RECT 664.950 556.950 667.050 557.400 ;
        RECT 623.400 555.600 624.600 556.950 ;
        RECT 581.400 554.400 624.600 555.600 ;
        RECT 625.950 555.600 628.050 556.050 ;
        RECT 685.950 555.600 688.050 556.050 ;
        RECT 625.950 554.400 688.050 555.600 ;
        RECT 424.950 553.950 427.050 554.400 ;
        RECT 466.950 553.950 469.050 554.400 ;
        RECT 487.950 553.950 490.050 554.400 ;
        RECT 625.950 553.950 628.050 554.400 ;
        RECT 685.950 553.950 688.050 554.400 ;
        RECT 709.950 555.600 712.050 556.050 ;
        RECT 742.950 555.600 745.050 556.050 ;
        RECT 709.950 554.400 745.050 555.600 ;
        RECT 709.950 553.950 712.050 554.400 ;
        RECT 742.950 553.950 745.050 554.400 ;
        RECT 94.950 552.600 97.050 553.050 ;
        RECT 124.950 552.600 127.050 553.050 ;
        RECT 94.950 551.400 127.050 552.600 ;
        RECT 94.950 550.950 97.050 551.400 ;
        RECT 124.950 550.950 127.050 551.400 ;
        RECT 184.950 552.600 187.050 553.050 ;
        RECT 205.950 552.600 208.050 553.050 ;
        RECT 184.950 551.400 208.050 552.600 ;
        RECT 184.950 550.950 187.050 551.400 ;
        RECT 205.950 550.950 208.050 551.400 ;
        RECT 250.950 552.600 253.050 553.050 ;
        RECT 292.950 552.600 295.050 553.050 ;
        RECT 316.950 552.600 319.050 553.050 ;
        RECT 250.950 551.400 319.050 552.600 ;
        RECT 250.950 550.950 253.050 551.400 ;
        RECT 292.950 550.950 295.050 551.400 ;
        RECT 316.950 550.950 319.050 551.400 ;
        RECT 331.950 552.600 334.050 553.050 ;
        RECT 370.950 552.600 373.050 553.050 ;
        RECT 412.950 552.600 415.050 553.050 ;
        RECT 331.950 551.400 415.050 552.600 ;
        RECT 331.950 550.950 334.050 551.400 ;
        RECT 370.950 550.950 373.050 551.400 ;
        RECT 412.950 550.950 415.050 551.400 ;
        RECT 508.950 552.600 511.050 553.050 ;
        RECT 538.950 552.600 541.050 553.050 ;
        RECT 508.950 551.400 541.050 552.600 ;
        RECT 508.950 550.950 511.050 551.400 ;
        RECT 538.950 550.950 541.050 551.400 ;
        RECT 625.950 552.600 628.050 553.050 ;
        RECT 655.950 552.600 658.050 553.050 ;
        RECT 625.950 551.400 658.050 552.600 ;
        RECT 625.950 550.950 628.050 551.400 ;
        RECT 655.950 550.950 658.050 551.400 ;
        RECT 664.950 552.600 667.050 553.050 ;
        RECT 718.950 552.600 721.050 553.050 ;
        RECT 664.950 551.400 721.050 552.600 ;
        RECT 664.950 550.950 667.050 551.400 ;
        RECT 718.950 550.950 721.050 551.400 ;
        RECT 202.950 549.600 205.050 550.050 ;
        RECT 244.950 549.600 247.050 550.050 ;
        RECT 202.950 548.400 247.050 549.600 ;
        RECT 202.950 547.950 205.050 548.400 ;
        RECT 244.950 547.950 247.050 548.400 ;
        RECT 373.950 549.600 376.050 550.050 ;
        RECT 418.950 549.600 421.050 550.050 ;
        RECT 373.950 548.400 421.050 549.600 ;
        RECT 373.950 547.950 376.050 548.400 ;
        RECT 418.950 547.950 421.050 548.400 ;
        RECT 13.950 540.600 16.050 541.050 ;
        RECT 37.950 540.600 40.050 541.050 ;
        RECT 13.950 539.400 40.050 540.600 ;
        RECT 13.950 538.950 16.050 539.400 ;
        RECT 37.950 538.950 40.050 539.400 ;
        RECT 391.950 540.600 394.050 541.050 ;
        RECT 448.950 540.600 451.050 541.050 ;
        RECT 391.950 539.400 451.050 540.600 ;
        RECT 391.950 538.950 394.050 539.400 ;
        RECT 448.950 538.950 451.050 539.400 ;
        RECT 157.950 534.600 160.050 535.050 ;
        RECT 250.950 534.600 253.050 535.050 ;
        RECT 157.950 533.400 253.050 534.600 ;
        RECT 157.950 532.950 160.050 533.400 ;
        RECT 250.950 532.950 253.050 533.400 ;
        RECT 22.950 531.600 25.050 532.050 ;
        RECT 97.950 531.600 100.050 532.050 ;
        RECT 100.950 531.600 103.050 532.050 ;
        RECT 175.950 531.600 178.050 532.050 ;
        RECT 178.950 531.600 181.050 532.050 ;
        RECT 22.950 530.400 181.050 531.600 ;
        RECT 22.950 529.950 25.050 530.400 ;
        RECT 97.950 529.950 100.050 530.400 ;
        RECT 100.950 529.950 103.050 530.400 ;
        RECT 175.950 529.950 178.050 530.400 ;
        RECT 178.950 529.950 181.050 530.400 ;
        RECT 319.950 531.600 322.050 532.050 ;
        RECT 325.950 531.600 328.050 532.050 ;
        RECT 319.950 530.400 328.050 531.600 ;
        RECT 319.950 529.950 322.050 530.400 ;
        RECT 325.950 529.950 328.050 530.400 ;
        RECT 472.950 531.600 475.050 532.050 ;
        RECT 493.950 531.600 496.050 532.050 ;
        RECT 520.950 531.600 523.050 532.050 ;
        RECT 472.950 530.400 496.050 531.600 ;
        RECT 472.950 529.950 475.050 530.400 ;
        RECT 493.950 529.950 496.050 530.400 ;
        RECT 497.400 530.400 523.050 531.600 ;
        RECT 31.950 528.600 34.050 529.050 ;
        RECT 73.950 528.600 76.050 529.050 ;
        RECT 31.950 527.400 76.050 528.600 ;
        RECT 31.950 526.950 34.050 527.400 ;
        RECT 73.950 526.950 76.050 527.400 ;
        RECT 151.950 528.600 154.050 529.050 ;
        RECT 172.950 528.600 175.050 529.050 ;
        RECT 151.950 527.400 175.050 528.600 ;
        RECT 151.950 526.950 154.050 527.400 ;
        RECT 172.950 526.950 175.050 527.400 ;
        RECT 190.950 528.600 193.050 529.050 ;
        RECT 202.950 528.600 205.050 529.050 ;
        RECT 190.950 527.400 205.050 528.600 ;
        RECT 190.950 526.950 193.050 527.400 ;
        RECT 202.950 526.950 205.050 527.400 ;
        RECT 352.950 528.600 355.050 529.050 ;
        RECT 403.950 528.600 406.050 529.050 ;
        RECT 466.950 528.600 469.050 529.050 ;
        RECT 352.950 527.400 363.600 528.600 ;
        RECT 352.950 526.950 355.050 527.400 ;
        RECT 70.950 525.600 73.050 526.050 ;
        RECT 76.950 525.600 79.050 526.050 ;
        RECT 70.950 524.400 79.050 525.600 ;
        RECT 70.950 523.950 73.050 524.400 ;
        RECT 76.950 523.950 79.050 524.400 ;
        RECT 133.950 525.600 136.050 526.050 ;
        RECT 148.950 525.600 151.050 526.050 ;
        RECT 133.950 524.400 151.050 525.600 ;
        RECT 133.950 523.950 136.050 524.400 ;
        RECT 148.950 523.950 151.050 524.400 ;
        RECT 310.950 525.600 313.050 526.050 ;
        RECT 358.950 525.600 361.050 526.050 ;
        RECT 310.950 524.400 361.050 525.600 ;
        RECT 362.400 525.600 363.600 527.400 ;
        RECT 403.950 527.400 469.050 528.600 ;
        RECT 403.950 526.950 406.050 527.400 ;
        RECT 466.950 526.950 469.050 527.400 ;
        RECT 484.950 528.600 487.050 529.050 ;
        RECT 497.400 528.600 498.600 530.400 ;
        RECT 520.950 529.950 523.050 530.400 ;
        RECT 670.950 531.600 673.050 532.050 ;
        RECT 700.950 531.600 703.050 532.050 ;
        RECT 706.950 531.600 709.050 532.050 ;
        RECT 670.950 530.400 709.050 531.600 ;
        RECT 670.950 529.950 673.050 530.400 ;
        RECT 700.950 529.950 703.050 530.400 ;
        RECT 706.950 529.950 709.050 530.400 ;
        RECT 484.950 527.400 498.600 528.600 ;
        RECT 733.950 528.600 736.050 529.050 ;
        RECT 742.950 528.600 745.050 529.050 ;
        RECT 733.950 527.400 745.050 528.600 ;
        RECT 484.950 526.950 487.050 527.400 ;
        RECT 733.950 526.950 736.050 527.400 ;
        RECT 742.950 526.950 745.050 527.400 ;
        RECT 406.950 525.600 409.050 526.050 ;
        RECT 362.400 524.400 409.050 525.600 ;
        RECT 310.950 523.950 313.050 524.400 ;
        RECT 358.950 523.950 361.050 524.400 ;
        RECT 406.950 523.950 409.050 524.400 ;
        RECT 412.950 525.600 415.050 526.050 ;
        RECT 523.950 525.600 526.050 526.050 ;
        RECT 703.950 525.600 706.050 526.050 ;
        RECT 412.950 524.400 706.050 525.600 ;
        RECT 412.950 523.950 415.050 524.400 ;
        RECT 523.950 523.950 526.050 524.400 ;
        RECT 703.950 523.950 706.050 524.400 ;
        RECT 709.950 525.600 712.050 526.050 ;
        RECT 715.950 525.600 718.050 526.050 ;
        RECT 709.950 524.400 718.050 525.600 ;
        RECT 709.950 523.950 712.050 524.400 ;
        RECT 715.950 523.950 718.050 524.400 ;
        RECT 289.950 522.600 292.050 523.050 ;
        RECT 355.950 522.600 358.050 523.050 ;
        RECT 289.950 521.400 358.050 522.600 ;
        RECT 289.950 520.950 292.050 521.400 ;
        RECT 355.950 520.950 358.050 521.400 ;
        RECT 361.950 522.600 364.050 523.050 ;
        RECT 397.950 522.600 400.050 523.050 ;
        RECT 361.950 521.400 400.050 522.600 ;
        RECT 361.950 520.950 364.050 521.400 ;
        RECT 397.950 520.950 400.050 521.400 ;
        RECT 493.950 522.600 496.050 523.050 ;
        RECT 547.950 522.600 550.050 523.050 ;
        RECT 562.950 522.600 565.050 523.050 ;
        RECT 493.950 521.400 565.050 522.600 ;
        RECT 493.950 520.950 496.050 521.400 ;
        RECT 547.950 520.950 550.050 521.400 ;
        RECT 562.950 520.950 565.050 521.400 ;
        RECT 619.950 522.600 622.050 523.050 ;
        RECT 628.950 522.600 631.050 523.050 ;
        RECT 658.950 522.600 661.050 523.050 ;
        RECT 667.950 522.600 670.050 523.050 ;
        RECT 619.950 521.400 670.050 522.600 ;
        RECT 619.950 520.950 622.050 521.400 ;
        RECT 628.950 520.950 631.050 521.400 ;
        RECT 658.950 520.950 661.050 521.400 ;
        RECT 667.950 520.950 670.050 521.400 ;
        RECT 31.950 519.600 34.050 520.050 ;
        RECT 46.950 519.600 49.050 520.050 ;
        RECT 67.950 519.600 70.050 520.050 ;
        RECT 31.950 518.400 70.050 519.600 ;
        RECT 31.950 517.950 34.050 518.400 ;
        RECT 46.950 517.950 49.050 518.400 ;
        RECT 67.950 517.950 70.050 518.400 ;
        RECT 229.950 519.600 232.050 520.050 ;
        RECT 373.950 519.600 376.050 520.050 ;
        RECT 229.950 518.400 376.050 519.600 ;
        RECT 229.950 517.950 232.050 518.400 ;
        RECT 373.950 517.950 376.050 518.400 ;
        RECT 64.950 516.600 67.050 517.050 ;
        RECT 67.950 516.600 70.050 517.050 ;
        RECT 73.950 516.600 76.050 517.050 ;
        RECT 64.950 515.400 76.050 516.600 ;
        RECT 64.950 514.950 67.050 515.400 ;
        RECT 67.950 514.950 70.050 515.400 ;
        RECT 73.950 514.950 76.050 515.400 ;
        RECT 499.950 516.600 502.050 517.050 ;
        RECT 688.950 516.600 691.050 517.050 ;
        RECT 499.950 515.400 691.050 516.600 ;
        RECT 499.950 514.950 502.050 515.400 ;
        RECT 688.950 514.950 691.050 515.400 ;
        RECT 109.950 495.600 112.050 496.050 ;
        RECT 160.950 495.600 163.050 496.050 ;
        RECT 241.950 495.600 244.050 496.050 ;
        RECT 109.950 494.400 244.050 495.600 ;
        RECT 109.950 493.950 112.050 494.400 ;
        RECT 160.950 493.950 163.050 494.400 ;
        RECT 241.950 493.950 244.050 494.400 ;
        RECT 382.950 495.600 385.050 496.050 ;
        RECT 577.950 495.600 580.050 496.050 ;
        RECT 382.950 494.400 580.050 495.600 ;
        RECT 382.950 493.950 385.050 494.400 ;
        RECT 577.950 493.950 580.050 494.400 ;
        RECT 166.950 492.600 169.050 493.050 ;
        RECT 613.950 492.600 616.050 493.050 ;
        RECT 166.950 491.400 616.050 492.600 ;
        RECT 166.950 490.950 169.050 491.400 ;
        RECT 613.950 490.950 616.050 491.400 ;
        RECT 628.950 492.600 631.050 493.050 ;
        RECT 661.950 492.600 664.050 493.050 ;
        RECT 628.950 491.400 664.050 492.600 ;
        RECT 628.950 490.950 631.050 491.400 ;
        RECT 661.950 490.950 664.050 491.400 ;
        RECT 109.950 489.600 112.050 490.050 ;
        RECT 112.950 489.600 115.050 490.050 ;
        RECT 154.950 489.600 157.050 490.050 ;
        RECT 163.950 489.600 166.050 490.050 ;
        RECT 229.950 489.600 232.050 490.050 ;
        RECT 109.950 488.400 166.050 489.600 ;
        RECT 109.950 487.950 112.050 488.400 ;
        RECT 112.950 487.950 115.050 488.400 ;
        RECT 154.950 487.950 157.050 488.400 ;
        RECT 163.950 487.950 166.050 488.400 ;
        RECT 227.400 488.400 232.050 489.600 ;
        RECT 61.950 486.600 64.050 487.050 ;
        RECT 67.950 486.600 70.050 487.050 ;
        RECT 61.950 485.400 70.050 486.600 ;
        RECT 61.950 484.950 64.050 485.400 ;
        RECT 67.950 484.950 70.050 485.400 ;
        RECT 115.950 486.600 118.050 487.050 ;
        RECT 157.950 486.600 160.050 487.050 ;
        RECT 115.950 485.400 160.050 486.600 ;
        RECT 115.950 484.950 118.050 485.400 ;
        RECT 157.950 484.950 160.050 485.400 ;
        RECT 227.400 484.050 228.600 488.400 ;
        RECT 229.950 487.950 232.050 488.400 ;
        RECT 262.950 489.600 265.050 490.050 ;
        RECT 268.950 489.600 271.050 490.050 ;
        RECT 274.950 489.600 277.050 490.050 ;
        RECT 262.950 488.400 277.050 489.600 ;
        RECT 262.950 487.950 265.050 488.400 ;
        RECT 268.950 487.950 271.050 488.400 ;
        RECT 274.950 487.950 277.050 488.400 ;
        RECT 358.950 489.600 361.050 490.050 ;
        RECT 427.950 489.600 430.050 490.050 ;
        RECT 358.950 488.400 430.050 489.600 ;
        RECT 358.950 487.950 361.050 488.400 ;
        RECT 427.950 487.950 430.050 488.400 ;
        RECT 457.950 489.600 460.050 490.050 ;
        RECT 478.950 489.600 481.050 490.050 ;
        RECT 496.950 489.600 499.050 490.050 ;
        RECT 457.950 488.400 499.050 489.600 ;
        RECT 457.950 487.950 460.050 488.400 ;
        RECT 478.950 487.950 481.050 488.400 ;
        RECT 496.950 487.950 499.050 488.400 ;
        RECT 502.950 489.600 505.050 490.050 ;
        RECT 529.950 489.600 532.050 490.050 ;
        RECT 538.950 489.600 541.050 490.050 ;
        RECT 640.950 489.600 643.050 490.050 ;
        RECT 658.950 489.600 661.050 490.050 ;
        RECT 502.950 488.400 541.050 489.600 ;
        RECT 502.950 487.950 505.050 488.400 ;
        RECT 529.950 487.950 532.050 488.400 ;
        RECT 538.950 487.950 541.050 488.400 ;
        RECT 605.400 488.400 621.600 489.600 ;
        RECT 229.950 486.600 232.050 487.050 ;
        RECT 259.950 486.600 262.050 487.050 ;
        RECT 229.950 485.400 262.050 486.600 ;
        RECT 229.950 484.950 232.050 485.400 ;
        RECT 259.950 484.950 262.050 485.400 ;
        RECT 370.950 486.600 373.050 487.050 ;
        RECT 415.950 486.600 418.050 487.050 ;
        RECT 370.950 485.400 418.050 486.600 ;
        RECT 370.950 484.950 373.050 485.400 ;
        RECT 415.950 484.950 418.050 485.400 ;
        RECT 541.950 486.600 544.050 487.050 ;
        RECT 605.400 486.600 606.600 488.400 ;
        RECT 620.400 487.050 621.600 488.400 ;
        RECT 640.950 488.400 661.050 489.600 ;
        RECT 640.950 487.950 643.050 488.400 ;
        RECT 658.950 487.950 661.050 488.400 ;
        RECT 664.950 489.600 667.050 490.050 ;
        RECT 670.950 489.600 673.050 490.050 ;
        RECT 664.950 488.400 673.050 489.600 ;
        RECT 664.950 487.950 667.050 488.400 ;
        RECT 670.950 487.950 673.050 488.400 ;
        RECT 541.950 485.400 606.600 486.600 ;
        RECT 607.950 486.600 610.050 487.050 ;
        RECT 613.950 486.600 616.050 487.050 ;
        RECT 607.950 485.400 616.050 486.600 ;
        RECT 541.950 484.950 544.050 485.400 ;
        RECT 607.950 484.950 610.050 485.400 ;
        RECT 613.950 484.950 616.050 485.400 ;
        RECT 619.950 484.950 622.050 487.050 ;
        RECT 631.950 486.600 634.050 487.050 ;
        RECT 661.950 486.600 664.050 487.050 ;
        RECT 631.950 485.400 664.050 486.600 ;
        RECT 631.950 484.950 634.050 485.400 ;
        RECT 661.950 484.950 664.050 485.400 ;
        RECT 64.950 483.600 67.050 484.050 ;
        RECT 106.950 483.600 109.050 484.050 ;
        RECT 64.950 482.400 109.050 483.600 ;
        RECT 64.950 481.950 67.050 482.400 ;
        RECT 106.950 481.950 109.050 482.400 ;
        RECT 226.950 481.950 229.050 484.050 ;
        RECT 235.950 483.600 238.050 484.050 ;
        RECT 253.950 483.600 256.050 484.050 ;
        RECT 235.950 482.400 256.050 483.600 ;
        RECT 235.950 481.950 238.050 482.400 ;
        RECT 253.950 481.950 256.050 482.400 ;
        RECT 295.950 483.600 298.050 484.050 ;
        RECT 355.950 483.600 358.050 484.050 ;
        RECT 295.950 482.400 358.050 483.600 ;
        RECT 295.950 481.950 298.050 482.400 ;
        RECT 355.950 481.950 358.050 482.400 ;
        RECT 361.950 483.600 364.050 484.050 ;
        RECT 367.950 483.600 370.050 484.050 ;
        RECT 361.950 482.400 370.050 483.600 ;
        RECT 361.950 481.950 364.050 482.400 ;
        RECT 367.950 481.950 370.050 482.400 ;
        RECT 445.950 483.600 448.050 484.050 ;
        RECT 460.950 483.600 463.050 484.050 ;
        RECT 502.950 483.600 505.050 484.050 ;
        RECT 445.950 482.400 505.050 483.600 ;
        RECT 445.950 481.950 448.050 482.400 ;
        RECT 460.950 481.950 463.050 482.400 ;
        RECT 502.950 481.950 505.050 482.400 ;
        RECT 616.950 483.600 619.050 484.050 ;
        RECT 733.950 483.600 736.050 484.050 ;
        RECT 616.950 482.400 736.050 483.600 ;
        RECT 616.950 481.950 619.050 482.400 ;
        RECT 733.950 481.950 736.050 482.400 ;
        RECT 13.950 480.600 16.050 481.050 ;
        RECT 70.950 480.600 73.050 481.050 ;
        RECT 13.950 479.400 73.050 480.600 ;
        RECT 13.950 478.950 16.050 479.400 ;
        RECT 70.950 478.950 73.050 479.400 ;
        RECT 94.950 480.600 97.050 481.050 ;
        RECT 112.950 480.600 115.050 481.050 ;
        RECT 94.950 479.400 115.050 480.600 ;
        RECT 94.950 478.950 97.050 479.400 ;
        RECT 112.950 478.950 115.050 479.400 ;
        RECT 175.950 480.600 178.050 481.050 ;
        RECT 232.950 480.600 235.050 481.050 ;
        RECT 175.950 479.400 235.050 480.600 ;
        RECT 175.950 478.950 178.050 479.400 ;
        RECT 232.950 478.950 235.050 479.400 ;
        RECT 301.950 480.600 304.050 481.050 ;
        RECT 370.950 480.600 373.050 481.050 ;
        RECT 301.950 479.400 373.050 480.600 ;
        RECT 301.950 478.950 304.050 479.400 ;
        RECT 370.950 478.950 373.050 479.400 ;
        RECT 547.950 480.600 550.050 481.050 ;
        RECT 589.950 480.600 592.050 481.050 ;
        RECT 610.950 480.600 613.050 481.050 ;
        RECT 670.950 480.600 673.050 481.050 ;
        RECT 703.950 480.600 706.050 481.050 ;
        RECT 547.950 479.400 706.050 480.600 ;
        RECT 547.950 478.950 550.050 479.400 ;
        RECT 589.950 478.950 592.050 479.400 ;
        RECT 610.950 478.950 613.050 479.400 ;
        RECT 670.950 478.950 673.050 479.400 ;
        RECT 703.950 478.950 706.050 479.400 ;
        RECT 268.950 477.600 271.050 478.050 ;
        RECT 271.950 477.600 274.050 478.050 ;
        RECT 313.950 477.600 316.050 478.050 ;
        RECT 268.950 476.400 316.050 477.600 ;
        RECT 268.950 475.950 271.050 476.400 ;
        RECT 271.950 475.950 274.050 476.400 ;
        RECT 313.950 475.950 316.050 476.400 ;
        RECT 352.950 477.600 355.050 478.050 ;
        RECT 415.950 477.600 418.050 478.050 ;
        RECT 352.950 476.400 418.050 477.600 ;
        RECT 352.950 475.950 355.050 476.400 ;
        RECT 415.950 475.950 418.050 476.400 ;
        RECT 580.950 477.600 583.050 478.050 ;
        RECT 670.950 477.600 673.050 478.050 ;
        RECT 580.950 476.400 673.050 477.600 ;
        RECT 580.950 475.950 583.050 476.400 ;
        RECT 670.950 475.950 673.050 476.400 ;
        RECT 19.950 474.600 22.050 475.050 ;
        RECT 22.950 474.600 25.050 475.050 ;
        RECT 52.950 474.600 55.050 475.050 ;
        RECT 19.950 473.400 55.050 474.600 ;
        RECT 19.950 472.950 22.050 473.400 ;
        RECT 22.950 472.950 25.050 473.400 ;
        RECT 52.950 472.950 55.050 473.400 ;
        RECT 406.950 474.600 409.050 475.050 ;
        RECT 460.950 474.600 463.050 475.050 ;
        RECT 406.950 473.400 463.050 474.600 ;
        RECT 406.950 472.950 409.050 473.400 ;
        RECT 460.950 472.950 463.050 473.400 ;
        RECT 559.950 471.600 562.050 472.050 ;
        RECT 583.950 471.600 586.050 472.050 ;
        RECT 559.950 470.400 586.050 471.600 ;
        RECT 559.950 469.950 562.050 470.400 ;
        RECT 583.950 469.950 586.050 470.400 ;
        RECT 751.950 465.600 754.050 466.050 ;
        RECT 760.950 465.600 763.050 466.050 ;
        RECT 751.950 464.400 763.050 465.600 ;
        RECT 751.950 463.950 754.050 464.400 ;
        RECT 760.950 463.950 763.050 464.400 ;
        RECT 217.950 462.600 220.050 463.050 ;
        RECT 382.950 462.600 385.050 463.050 ;
        RECT 217.950 461.400 385.050 462.600 ;
        RECT 217.950 460.950 220.050 461.400 ;
        RECT 382.950 460.950 385.050 461.400 ;
        RECT 745.950 462.600 748.050 463.050 ;
        RECT 757.950 462.600 760.050 463.050 ;
        RECT 745.950 461.400 760.050 462.600 ;
        RECT 745.950 460.950 748.050 461.400 ;
        RECT 757.950 460.950 760.050 461.400 ;
        RECT 292.950 459.600 295.050 460.050 ;
        RECT 304.950 459.600 307.050 460.050 ;
        RECT 292.950 458.400 307.050 459.600 ;
        RECT 292.950 457.950 295.050 458.400 ;
        RECT 304.950 457.950 307.050 458.400 ;
        RECT 313.950 459.600 316.050 460.050 ;
        RECT 343.950 459.600 346.050 460.050 ;
        RECT 313.950 458.400 346.050 459.600 ;
        RECT 313.950 457.950 316.050 458.400 ;
        RECT 343.950 457.950 346.050 458.400 ;
        RECT 544.950 459.600 547.050 460.050 ;
        RECT 625.950 459.600 628.050 460.050 ;
        RECT 544.950 458.400 628.050 459.600 ;
        RECT 544.950 457.950 547.050 458.400 ;
        RECT 625.950 457.950 628.050 458.400 ;
        RECT 742.950 459.600 745.050 460.050 ;
        RECT 757.950 459.600 760.050 460.050 ;
        RECT 742.950 458.400 760.050 459.600 ;
        RECT 742.950 457.950 745.050 458.400 ;
        RECT 757.950 457.950 760.050 458.400 ;
        RECT 298.950 456.600 301.050 457.050 ;
        RECT 310.950 456.600 313.050 457.050 ;
        RECT 298.950 455.400 313.050 456.600 ;
        RECT 298.950 454.950 301.050 455.400 ;
        RECT 310.950 454.950 313.050 455.400 ;
        RECT 340.950 454.950 343.050 457.050 ;
        RECT 445.950 456.600 448.050 457.050 ;
        RECT 451.950 456.600 454.050 457.050 ;
        RECT 454.950 456.600 457.050 457.050 ;
        RECT 445.950 455.400 457.050 456.600 ;
        RECT 445.950 454.950 448.050 455.400 ;
        RECT 451.950 454.950 454.050 455.400 ;
        RECT 454.950 454.950 457.050 455.400 ;
        RECT 502.950 456.600 505.050 457.050 ;
        RECT 544.950 456.600 547.050 457.050 ;
        RECT 502.950 455.400 547.050 456.600 ;
        RECT 502.950 454.950 505.050 455.400 ;
        RECT 544.950 454.950 547.050 455.400 ;
        RECT 574.950 456.600 577.050 457.050 ;
        RECT 589.950 456.600 592.050 457.050 ;
        RECT 631.950 456.600 634.050 457.050 ;
        RECT 658.950 456.600 661.050 457.050 ;
        RECT 574.950 455.400 661.050 456.600 ;
        RECT 574.950 454.950 577.050 455.400 ;
        RECT 589.950 454.950 592.050 455.400 ;
        RECT 631.950 454.950 634.050 455.400 ;
        RECT 658.950 454.950 661.050 455.400 ;
        RECT 739.950 456.600 742.050 457.050 ;
        RECT 751.950 456.600 754.050 457.050 ;
        RECT 739.950 455.400 754.050 456.600 ;
        RECT 739.950 454.950 742.050 455.400 ;
        RECT 751.950 454.950 754.050 455.400 ;
        RECT 94.950 453.600 97.050 454.050 ;
        RECT 118.950 453.600 121.050 454.050 ;
        RECT 94.950 452.400 121.050 453.600 ;
        RECT 94.950 451.950 97.050 452.400 ;
        RECT 118.950 451.950 121.050 452.400 ;
        RECT 139.950 453.600 142.050 454.050 ;
        RECT 172.950 453.600 175.050 454.050 ;
        RECT 139.950 452.400 175.050 453.600 ;
        RECT 139.950 451.950 142.050 452.400 ;
        RECT 172.950 451.950 175.050 452.400 ;
        RECT 277.950 453.600 280.050 454.050 ;
        RECT 295.950 453.600 298.050 454.050 ;
        RECT 277.950 452.400 298.050 453.600 ;
        RECT 277.950 451.950 280.050 452.400 ;
        RECT 295.950 451.950 298.050 452.400 ;
        RECT 301.950 453.600 304.050 454.050 ;
        RECT 313.950 453.600 316.050 454.050 ;
        RECT 301.950 452.400 316.050 453.600 ;
        RECT 341.400 453.600 342.600 454.950 ;
        RECT 343.950 453.600 346.050 454.050 ;
        RECT 341.400 452.400 346.050 453.600 ;
        RECT 301.950 451.950 304.050 452.400 ;
        RECT 313.950 451.950 316.050 452.400 ;
        RECT 343.950 451.950 346.050 452.400 ;
        RECT 538.950 453.600 541.050 454.050 ;
        RECT 580.950 453.600 583.050 454.050 ;
        RECT 538.950 452.400 583.050 453.600 ;
        RECT 538.950 451.950 541.050 452.400 ;
        RECT 580.950 451.950 583.050 452.400 ;
        RECT 586.950 453.600 589.050 454.050 ;
        RECT 667.950 453.600 670.050 454.050 ;
        RECT 586.950 452.400 670.050 453.600 ;
        RECT 586.950 451.950 589.050 452.400 ;
        RECT 667.950 451.950 670.050 452.400 ;
        RECT 709.950 453.600 712.050 454.050 ;
        RECT 748.950 453.600 751.050 454.050 ;
        RECT 709.950 452.400 751.050 453.600 ;
        RECT 709.950 451.950 712.050 452.400 ;
        RECT 748.950 451.950 751.050 452.400 ;
        RECT 271.950 450.600 274.050 451.050 ;
        RECT 358.950 450.600 361.050 451.050 ;
        RECT 271.950 449.400 361.050 450.600 ;
        RECT 271.950 448.950 274.050 449.400 ;
        RECT 358.950 448.950 361.050 449.400 ;
        RECT 418.950 450.600 421.050 451.050 ;
        RECT 427.950 450.600 430.050 451.050 ;
        RECT 418.950 449.400 430.050 450.600 ;
        RECT 418.950 448.950 421.050 449.400 ;
        RECT 427.950 448.950 430.050 449.400 ;
        RECT 463.950 450.600 466.050 451.050 ;
        RECT 541.950 450.600 544.050 451.050 ;
        RECT 463.950 449.400 544.050 450.600 ;
        RECT 463.950 448.950 466.050 449.400 ;
        RECT 541.950 448.950 544.050 449.400 ;
        RECT 667.950 450.600 670.050 451.050 ;
        RECT 754.950 450.600 757.050 451.050 ;
        RECT 667.950 449.400 757.050 450.600 ;
        RECT 667.950 448.950 670.050 449.400 ;
        RECT 754.950 448.950 757.050 449.400 ;
        RECT 130.950 447.600 133.050 448.050 ;
        RECT 151.950 447.600 154.050 448.050 ;
        RECT 256.950 447.600 259.050 448.050 ;
        RECT 130.950 446.400 259.050 447.600 ;
        RECT 130.950 445.950 133.050 446.400 ;
        RECT 151.950 445.950 154.050 446.400 ;
        RECT 256.950 445.950 259.050 446.400 ;
        RECT 340.950 447.600 343.050 448.050 ;
        RECT 349.950 447.600 352.050 448.050 ;
        RECT 535.950 447.600 538.050 448.050 ;
        RECT 340.950 446.400 538.050 447.600 ;
        RECT 340.950 445.950 343.050 446.400 ;
        RECT 349.950 445.950 352.050 446.400 ;
        RECT 535.950 445.950 538.050 446.400 ;
        RECT 484.950 426.600 487.050 427.050 ;
        RECT 499.950 426.600 502.050 427.050 ;
        RECT 484.950 425.400 502.050 426.600 ;
        RECT 484.950 424.950 487.050 425.400 ;
        RECT 499.950 424.950 502.050 425.400 ;
        RECT 322.950 423.600 325.050 424.050 ;
        RECT 649.950 423.600 652.050 424.050 ;
        RECT 322.950 422.400 652.050 423.600 ;
        RECT 322.950 421.950 325.050 422.400 ;
        RECT 649.950 421.950 652.050 422.400 ;
        RECT 175.950 420.600 178.050 421.050 ;
        RECT 196.950 420.600 199.050 421.050 ;
        RECT 493.950 420.600 496.050 421.050 ;
        RECT 499.950 420.600 502.050 421.050 ;
        RECT 175.950 419.400 502.050 420.600 ;
        RECT 175.950 418.950 178.050 419.400 ;
        RECT 196.950 418.950 199.050 419.400 ;
        RECT 493.950 418.950 496.050 419.400 ;
        RECT 499.950 418.950 502.050 419.400 ;
        RECT 103.950 417.600 106.050 418.050 ;
        RECT 166.950 417.600 169.050 418.050 ;
        RECT 103.950 416.400 169.050 417.600 ;
        RECT 103.950 415.950 106.050 416.400 ;
        RECT 166.950 415.950 169.050 416.400 ;
        RECT 190.950 417.600 193.050 418.050 ;
        RECT 208.950 417.600 211.050 418.050 ;
        RECT 190.950 416.400 211.050 417.600 ;
        RECT 190.950 415.950 193.050 416.400 ;
        RECT 208.950 415.950 211.050 416.400 ;
        RECT 310.950 417.600 313.050 418.050 ;
        RECT 316.950 417.600 319.050 418.050 ;
        RECT 310.950 416.400 319.050 417.600 ;
        RECT 310.950 415.950 313.050 416.400 ;
        RECT 316.950 415.950 319.050 416.400 ;
        RECT 493.950 417.600 496.050 418.050 ;
        RECT 520.950 417.600 523.050 418.050 ;
        RECT 493.950 416.400 523.050 417.600 ;
        RECT 493.950 415.950 496.050 416.400 ;
        RECT 520.950 415.950 523.050 416.400 ;
        RECT 67.950 414.600 70.050 415.050 ;
        RECT 127.950 414.600 130.050 415.050 ;
        RECT 67.950 413.400 130.050 414.600 ;
        RECT 67.950 412.950 70.050 413.400 ;
        RECT 127.950 412.950 130.050 413.400 ;
        RECT 148.950 414.600 151.050 415.050 ;
        RECT 154.950 414.600 157.050 415.050 ;
        RECT 271.950 414.600 274.050 415.050 ;
        RECT 148.950 413.400 157.050 414.600 ;
        RECT 148.950 412.950 151.050 413.400 ;
        RECT 154.950 412.950 157.050 413.400 ;
        RECT 197.400 413.400 274.050 414.600 ;
        RECT 22.950 411.600 25.050 412.050 ;
        RECT 55.950 411.600 58.050 412.050 ;
        RECT 22.950 410.400 58.050 411.600 ;
        RECT 22.950 409.950 25.050 410.400 ;
        RECT 55.950 409.950 58.050 410.400 ;
        RECT 85.950 411.600 88.050 412.050 ;
        RECT 145.950 411.600 148.050 412.050 ;
        RECT 85.950 410.400 148.050 411.600 ;
        RECT 85.950 409.950 88.050 410.400 ;
        RECT 145.950 409.950 148.050 410.400 ;
        RECT 151.950 411.600 154.050 412.050 ;
        RECT 175.950 411.600 178.050 412.050 ;
        RECT 151.950 410.400 178.050 411.600 ;
        RECT 151.950 409.950 154.050 410.400 ;
        RECT 175.950 409.950 178.050 410.400 ;
        RECT 193.950 411.600 196.050 412.050 ;
        RECT 197.400 411.600 198.600 413.400 ;
        RECT 271.950 412.950 274.050 413.400 ;
        RECT 274.950 414.600 277.050 415.050 ;
        RECT 319.950 414.600 322.050 415.050 ;
        RECT 274.950 413.400 322.050 414.600 ;
        RECT 274.950 412.950 277.050 413.400 ;
        RECT 319.950 412.950 322.050 413.400 ;
        RECT 358.950 414.600 361.050 415.050 ;
        RECT 400.950 414.600 403.050 415.050 ;
        RECT 358.950 413.400 403.050 414.600 ;
        RECT 358.950 412.950 361.050 413.400 ;
        RECT 400.950 412.950 403.050 413.400 ;
        RECT 451.950 414.600 454.050 415.050 ;
        RECT 574.950 414.600 577.050 415.050 ;
        RECT 451.950 413.400 577.050 414.600 ;
        RECT 451.950 412.950 454.050 413.400 ;
        RECT 574.950 412.950 577.050 413.400 ;
        RECT 580.950 414.600 583.050 415.050 ;
        RECT 607.950 414.600 610.050 415.050 ;
        RECT 613.950 414.600 616.050 415.050 ;
        RECT 580.950 413.400 616.050 414.600 ;
        RECT 580.950 412.950 583.050 413.400 ;
        RECT 607.950 412.950 610.050 413.400 ;
        RECT 613.950 412.950 616.050 413.400 ;
        RECT 193.950 410.400 198.600 411.600 ;
        RECT 199.950 411.600 202.050 412.050 ;
        RECT 214.950 411.600 217.050 412.050 ;
        RECT 199.950 410.400 217.050 411.600 ;
        RECT 193.950 409.950 196.050 410.400 ;
        RECT 199.950 409.950 202.050 410.400 ;
        RECT 214.950 409.950 217.050 410.400 ;
        RECT 313.950 411.600 316.050 412.050 ;
        RECT 397.950 411.600 400.050 412.050 ;
        RECT 463.950 411.600 466.050 412.050 ;
        RECT 313.950 410.400 466.050 411.600 ;
        RECT 313.950 409.950 316.050 410.400 ;
        RECT 397.950 409.950 400.050 410.400 ;
        RECT 463.950 409.950 466.050 410.400 ;
        RECT 490.950 411.600 493.050 412.050 ;
        RECT 511.950 411.600 514.050 412.050 ;
        RECT 490.950 410.400 514.050 411.600 ;
        RECT 490.950 409.950 493.050 410.400 ;
        RECT 511.950 409.950 514.050 410.400 ;
        RECT 55.950 408.600 58.050 409.050 ;
        RECT 91.950 408.600 94.050 409.050 ;
        RECT 55.950 407.400 94.050 408.600 ;
        RECT 55.950 406.950 58.050 407.400 ;
        RECT 91.950 406.950 94.050 407.400 ;
        RECT 163.950 408.600 166.050 409.050 ;
        RECT 178.950 408.600 181.050 409.050 ;
        RECT 163.950 407.400 181.050 408.600 ;
        RECT 163.950 406.950 166.050 407.400 ;
        RECT 178.950 406.950 181.050 407.400 ;
        RECT 232.950 408.600 235.050 409.050 ;
        RECT 262.950 408.600 265.050 409.050 ;
        RECT 232.950 407.400 265.050 408.600 ;
        RECT 232.950 406.950 235.050 407.400 ;
        RECT 262.950 406.950 265.050 407.400 ;
        RECT 409.950 408.600 412.050 409.050 ;
        RECT 568.950 408.600 571.050 409.050 ;
        RECT 409.950 407.400 571.050 408.600 ;
        RECT 409.950 406.950 412.050 407.400 ;
        RECT 568.950 406.950 571.050 407.400 ;
        RECT 700.950 408.600 703.050 409.050 ;
        RECT 736.950 408.600 739.050 409.050 ;
        RECT 700.950 407.400 739.050 408.600 ;
        RECT 700.950 406.950 703.050 407.400 ;
        RECT 736.950 406.950 739.050 407.400 ;
        RECT 127.950 405.600 130.050 406.050 ;
        RECT 235.950 405.600 238.050 406.050 ;
        RECT 352.950 405.600 355.050 406.050 ;
        RECT 373.950 405.600 376.050 406.050 ;
        RECT 127.950 404.400 376.050 405.600 ;
        RECT 127.950 403.950 130.050 404.400 ;
        RECT 235.950 403.950 238.050 404.400 ;
        RECT 352.950 403.950 355.050 404.400 ;
        RECT 373.950 403.950 376.050 404.400 ;
        RECT 34.950 402.600 37.050 403.050 ;
        RECT 67.950 402.600 70.050 403.050 ;
        RECT 229.950 402.600 232.050 403.050 ;
        RECT 244.950 402.600 247.050 403.050 ;
        RECT 34.950 401.400 247.050 402.600 ;
        RECT 34.950 400.950 37.050 401.400 ;
        RECT 67.950 400.950 70.050 401.400 ;
        RECT 229.950 400.950 232.050 401.400 ;
        RECT 244.950 400.950 247.050 401.400 ;
        RECT 730.950 402.600 733.050 403.050 ;
        RECT 739.950 402.600 742.050 403.050 ;
        RECT 730.950 401.400 742.050 402.600 ;
        RECT 730.950 400.950 733.050 401.400 ;
        RECT 739.950 400.950 742.050 401.400 ;
        RECT 13.950 399.600 16.050 400.050 ;
        RECT 37.950 399.600 40.050 400.050 ;
        RECT 13.950 398.400 40.050 399.600 ;
        RECT 13.950 397.950 16.050 398.400 ;
        RECT 37.950 397.950 40.050 398.400 ;
        RECT 49.950 399.600 52.050 400.050 ;
        RECT 79.950 399.600 82.050 400.050 ;
        RECT 49.950 398.400 82.050 399.600 ;
        RECT 49.950 397.950 52.050 398.400 ;
        RECT 79.950 397.950 82.050 398.400 ;
        RECT 313.950 396.600 316.050 397.050 ;
        RECT 370.950 396.600 373.050 397.050 ;
        RECT 403.950 396.600 406.050 397.050 ;
        RECT 436.950 396.600 439.050 397.050 ;
        RECT 514.950 396.600 517.050 397.050 ;
        RECT 517.950 396.600 520.050 397.050 ;
        RECT 565.950 396.600 568.050 397.050 ;
        RECT 313.950 395.400 568.050 396.600 ;
        RECT 313.950 394.950 316.050 395.400 ;
        RECT 370.950 394.950 373.050 395.400 ;
        RECT 403.950 394.950 406.050 395.400 ;
        RECT 436.950 394.950 439.050 395.400 ;
        RECT 514.950 394.950 517.050 395.400 ;
        RECT 517.950 394.950 520.050 395.400 ;
        RECT 565.950 394.950 568.050 395.400 ;
        RECT 418.950 393.600 421.050 394.050 ;
        RECT 502.950 393.600 505.050 394.050 ;
        RECT 622.950 393.600 625.050 394.050 ;
        RECT 418.950 392.400 625.050 393.600 ;
        RECT 418.950 391.950 421.050 392.400 ;
        RECT 502.950 391.950 505.050 392.400 ;
        RECT 622.950 391.950 625.050 392.400 ;
        RECT 703.950 393.600 706.050 394.050 ;
        RECT 712.950 393.600 715.050 394.050 ;
        RECT 703.950 392.400 715.050 393.600 ;
        RECT 703.950 391.950 706.050 392.400 ;
        RECT 712.950 391.950 715.050 392.400 ;
        RECT 289.950 390.600 292.050 391.050 ;
        RECT 364.950 390.600 367.050 391.050 ;
        RECT 370.950 390.600 373.050 391.050 ;
        RECT 289.950 389.400 373.050 390.600 ;
        RECT 289.950 388.950 292.050 389.400 ;
        RECT 364.950 388.950 367.050 389.400 ;
        RECT 370.950 388.950 373.050 389.400 ;
        RECT 544.950 390.600 547.050 391.050 ;
        RECT 613.950 390.600 616.050 391.050 ;
        RECT 544.950 389.400 616.050 390.600 ;
        RECT 544.950 388.950 547.050 389.400 ;
        RECT 613.950 388.950 616.050 389.400 ;
        RECT 637.950 390.600 640.050 391.050 ;
        RECT 655.950 390.600 658.050 391.050 ;
        RECT 637.950 389.400 658.050 390.600 ;
        RECT 637.950 388.950 640.050 389.400 ;
        RECT 655.950 388.950 658.050 389.400 ;
        RECT 697.950 390.600 700.050 391.050 ;
        RECT 712.950 390.600 715.050 391.050 ;
        RECT 742.950 390.600 745.050 391.050 ;
        RECT 697.950 389.400 745.050 390.600 ;
        RECT 697.950 388.950 700.050 389.400 ;
        RECT 712.950 388.950 715.050 389.400 ;
        RECT 742.950 388.950 745.050 389.400 ;
        RECT 43.950 387.600 46.050 388.050 ;
        RECT 94.950 387.600 97.050 388.050 ;
        RECT 43.950 386.400 97.050 387.600 ;
        RECT 43.950 385.950 46.050 386.400 ;
        RECT 94.950 385.950 97.050 386.400 ;
        RECT 163.950 387.600 166.050 388.050 ;
        RECT 196.950 387.600 199.050 388.050 ;
        RECT 202.950 387.600 205.050 388.050 ;
        RECT 163.950 386.400 205.050 387.600 ;
        RECT 163.950 385.950 166.050 386.400 ;
        RECT 196.950 385.950 199.050 386.400 ;
        RECT 202.950 385.950 205.050 386.400 ;
        RECT 283.950 387.600 286.050 388.050 ;
        RECT 286.950 387.600 289.050 388.050 ;
        RECT 331.950 387.600 334.050 388.050 ;
        RECT 283.950 386.400 334.050 387.600 ;
        RECT 283.950 385.950 286.050 386.400 ;
        RECT 286.950 385.950 289.050 386.400 ;
        RECT 331.950 385.950 334.050 386.400 ;
        RECT 559.950 387.600 562.050 388.050 ;
        RECT 571.950 387.600 574.050 388.050 ;
        RECT 559.950 386.400 574.050 387.600 ;
        RECT 559.950 385.950 562.050 386.400 ;
        RECT 571.950 385.950 574.050 386.400 ;
        RECT 580.950 387.600 583.050 388.050 ;
        RECT 610.950 387.600 613.050 388.050 ;
        RECT 580.950 386.400 613.050 387.600 ;
        RECT 580.950 385.950 583.050 386.400 ;
        RECT 610.950 385.950 613.050 386.400 ;
        RECT 658.950 387.600 661.050 388.050 ;
        RECT 691.950 387.600 694.050 388.050 ;
        RECT 658.950 386.400 694.050 387.600 ;
        RECT 658.950 385.950 661.050 386.400 ;
        RECT 691.950 385.950 694.050 386.400 ;
        RECT 34.950 384.600 37.050 385.050 ;
        RECT 46.950 384.600 49.050 385.050 ;
        RECT 34.950 383.400 49.050 384.600 ;
        RECT 34.950 382.950 37.050 383.400 ;
        RECT 46.950 382.950 49.050 383.400 ;
        RECT 73.950 384.600 76.050 385.050 ;
        RECT 250.950 384.600 253.050 385.050 ;
        RECT 295.950 384.600 298.050 385.050 ;
        RECT 73.950 383.400 81.600 384.600 ;
        RECT 73.950 382.950 76.050 383.400 ;
        RECT 40.950 381.600 43.050 382.050 ;
        RECT 76.950 381.600 79.050 382.050 ;
        RECT 40.950 380.400 79.050 381.600 ;
        RECT 80.400 381.600 81.600 383.400 ;
        RECT 250.950 383.400 298.050 384.600 ;
        RECT 250.950 382.950 253.050 383.400 ;
        RECT 295.950 382.950 298.050 383.400 ;
        RECT 397.950 384.600 400.050 385.050 ;
        RECT 457.950 384.600 460.050 385.050 ;
        RECT 397.950 383.400 460.050 384.600 ;
        RECT 397.950 382.950 400.050 383.400 ;
        RECT 457.950 382.950 460.050 383.400 ;
        RECT 565.950 384.600 568.050 385.050 ;
        RECT 589.950 384.600 592.050 385.050 ;
        RECT 643.950 384.600 646.050 385.050 ;
        RECT 649.950 384.600 652.050 385.050 ;
        RECT 565.950 383.400 652.050 384.600 ;
        RECT 565.950 382.950 568.050 383.400 ;
        RECT 589.950 382.950 592.050 383.400 ;
        RECT 643.950 382.950 646.050 383.400 ;
        RECT 649.950 382.950 652.050 383.400 ;
        RECT 106.950 381.600 109.050 382.050 ;
        RECT 121.950 381.600 124.050 382.050 ;
        RECT 80.400 380.400 124.050 381.600 ;
        RECT 40.950 379.950 43.050 380.400 ;
        RECT 76.950 379.950 79.050 380.400 ;
        RECT 106.950 379.950 109.050 380.400 ;
        RECT 121.950 379.950 124.050 380.400 ;
        RECT 175.950 381.600 178.050 382.050 ;
        RECT 205.950 381.600 208.050 382.050 ;
        RECT 175.950 380.400 208.050 381.600 ;
        RECT 175.950 379.950 178.050 380.400 ;
        RECT 205.950 379.950 208.050 380.400 ;
        RECT 247.950 381.600 250.050 382.050 ;
        RECT 280.950 381.600 283.050 382.050 ;
        RECT 292.950 381.600 295.050 382.050 ;
        RECT 247.950 380.400 295.050 381.600 ;
        RECT 247.950 379.950 250.050 380.400 ;
        RECT 280.950 379.950 283.050 380.400 ;
        RECT 292.950 379.950 295.050 380.400 ;
        RECT 334.950 381.600 337.050 382.050 ;
        RECT 343.950 381.600 346.050 382.050 ;
        RECT 334.950 380.400 346.050 381.600 ;
        RECT 334.950 379.950 337.050 380.400 ;
        RECT 343.950 379.950 346.050 380.400 ;
        RECT 379.950 381.600 382.050 382.050 ;
        RECT 400.950 381.600 403.050 382.050 ;
        RECT 379.950 380.400 403.050 381.600 ;
        RECT 379.950 379.950 382.050 380.400 ;
        RECT 400.950 379.950 403.050 380.400 ;
        RECT 448.950 381.600 451.050 382.050 ;
        RECT 460.950 381.600 463.050 382.050 ;
        RECT 448.950 380.400 463.050 381.600 ;
        RECT 448.950 379.950 451.050 380.400 ;
        RECT 460.950 379.950 463.050 380.400 ;
        RECT 466.950 381.600 469.050 382.050 ;
        RECT 499.950 381.600 502.050 382.050 ;
        RECT 466.950 380.400 502.050 381.600 ;
        RECT 466.950 379.950 469.050 380.400 ;
        RECT 499.950 379.950 502.050 380.400 ;
        RECT 724.950 381.600 727.050 382.050 ;
        RECT 733.950 381.600 736.050 382.050 ;
        RECT 724.950 380.400 736.050 381.600 ;
        RECT 724.950 379.950 727.050 380.400 ;
        RECT 733.950 379.950 736.050 380.400 ;
        RECT 169.950 378.600 172.050 379.050 ;
        RECT 199.950 378.600 202.050 379.050 ;
        RECT 169.950 377.400 202.050 378.600 ;
        RECT 169.950 376.950 172.050 377.400 ;
        RECT 199.950 376.950 202.050 377.400 ;
        RECT 451.950 378.600 454.050 379.050 ;
        RECT 466.950 378.600 469.050 379.050 ;
        RECT 451.950 377.400 469.050 378.600 ;
        RECT 451.950 376.950 454.050 377.400 ;
        RECT 466.950 376.950 469.050 377.400 ;
        RECT 661.950 378.600 664.050 379.050 ;
        RECT 694.950 378.600 697.050 379.050 ;
        RECT 739.950 378.600 742.050 379.050 ;
        RECT 661.950 377.400 742.050 378.600 ;
        RECT 661.950 376.950 664.050 377.400 ;
        RECT 694.950 376.950 697.050 377.400 ;
        RECT 739.950 376.950 742.050 377.400 ;
        RECT 277.950 348.600 280.050 349.050 ;
        RECT 286.950 348.600 289.050 349.050 ;
        RECT 277.950 347.400 289.050 348.600 ;
        RECT 277.950 346.950 280.050 347.400 ;
        RECT 286.950 346.950 289.050 347.400 ;
        RECT 706.950 348.600 709.050 349.050 ;
        RECT 736.950 348.600 739.050 349.050 ;
        RECT 706.950 347.400 739.050 348.600 ;
        RECT 706.950 346.950 709.050 347.400 ;
        RECT 736.950 346.950 739.050 347.400 ;
        RECT 163.950 345.600 166.050 346.050 ;
        RECT 223.950 345.600 226.050 346.050 ;
        RECT 163.950 344.400 226.050 345.600 ;
        RECT 163.950 343.950 166.050 344.400 ;
        RECT 223.950 343.950 226.050 344.400 ;
        RECT 235.950 345.600 238.050 346.050 ;
        RECT 280.950 345.600 283.050 346.050 ;
        RECT 235.950 344.400 283.050 345.600 ;
        RECT 235.950 343.950 238.050 344.400 ;
        RECT 280.950 343.950 283.050 344.400 ;
        RECT 361.950 345.600 364.050 346.050 ;
        RECT 400.950 345.600 403.050 346.050 ;
        RECT 412.950 345.600 415.050 346.050 ;
        RECT 484.950 345.600 487.050 346.050 ;
        RECT 361.950 344.400 399.600 345.600 ;
        RECT 361.950 343.950 364.050 344.400 ;
        RECT 64.950 342.600 67.050 343.050 ;
        RECT 76.950 342.600 79.050 343.050 ;
        RECT 115.950 342.600 118.050 343.050 ;
        RECT 64.950 341.400 118.050 342.600 ;
        RECT 64.950 340.950 67.050 341.400 ;
        RECT 76.950 340.950 79.050 341.400 ;
        RECT 115.950 340.950 118.050 341.400 ;
        RECT 121.950 342.600 124.050 343.050 ;
        RECT 127.950 342.600 130.050 343.050 ;
        RECT 121.950 341.400 130.050 342.600 ;
        RECT 121.950 340.950 124.050 341.400 ;
        RECT 127.950 340.950 130.050 341.400 ;
        RECT 151.950 342.600 154.050 343.050 ;
        RECT 160.950 342.600 163.050 343.050 ;
        RECT 151.950 341.400 163.050 342.600 ;
        RECT 151.950 340.950 154.050 341.400 ;
        RECT 160.950 340.950 163.050 341.400 ;
        RECT 244.950 342.600 247.050 343.050 ;
        RECT 253.950 342.600 256.050 343.050 ;
        RECT 244.950 341.400 256.050 342.600 ;
        RECT 244.950 340.950 247.050 341.400 ;
        RECT 253.950 340.950 256.050 341.400 ;
        RECT 283.950 342.600 286.050 343.050 ;
        RECT 307.950 342.600 310.050 343.050 ;
        RECT 283.950 341.400 310.050 342.600 ;
        RECT 283.950 340.950 286.050 341.400 ;
        RECT 307.950 340.950 310.050 341.400 ;
        RECT 322.950 342.600 325.050 343.050 ;
        RECT 334.950 342.600 337.050 343.050 ;
        RECT 358.950 342.600 361.050 343.050 ;
        RECT 367.950 342.600 370.050 343.050 ;
        RECT 322.950 341.400 370.050 342.600 ;
        RECT 398.400 342.600 399.600 344.400 ;
        RECT 400.950 344.400 411.600 345.600 ;
        RECT 400.950 343.950 403.050 344.400 ;
        RECT 410.400 343.050 411.600 344.400 ;
        RECT 412.950 344.400 487.050 345.600 ;
        RECT 412.950 343.950 415.050 344.400 ;
        RECT 484.950 343.950 487.050 344.400 ;
        RECT 541.950 345.600 544.050 346.050 ;
        RECT 625.950 345.600 628.050 346.050 ;
        RECT 628.950 345.600 631.050 346.050 ;
        RECT 541.950 344.400 631.050 345.600 ;
        RECT 541.950 343.950 544.050 344.400 ;
        RECT 625.950 343.950 628.050 344.400 ;
        RECT 628.950 343.950 631.050 344.400 ;
        RECT 634.950 345.600 637.050 346.050 ;
        RECT 640.950 345.600 643.050 346.050 ;
        RECT 634.950 344.400 643.050 345.600 ;
        RECT 634.950 343.950 637.050 344.400 ;
        RECT 640.950 343.950 643.050 344.400 ;
        RECT 712.950 345.600 715.050 346.050 ;
        RECT 742.950 345.600 745.050 346.050 ;
        RECT 712.950 344.400 745.050 345.600 ;
        RECT 712.950 343.950 715.050 344.400 ;
        RECT 742.950 343.950 745.050 344.400 ;
        RECT 745.950 345.600 748.050 346.050 ;
        RECT 757.950 345.600 760.050 346.050 ;
        RECT 745.950 344.400 760.050 345.600 ;
        RECT 745.950 343.950 748.050 344.400 ;
        RECT 757.950 343.950 760.050 344.400 ;
        RECT 406.950 342.600 409.050 343.050 ;
        RECT 398.400 341.400 409.050 342.600 ;
        RECT 322.950 340.950 325.050 341.400 ;
        RECT 334.950 340.950 337.050 341.400 ;
        RECT 358.950 340.950 361.050 341.400 ;
        RECT 367.950 340.950 370.050 341.400 ;
        RECT 406.950 340.950 409.050 341.400 ;
        RECT 409.950 340.950 412.050 343.050 ;
        RECT 460.950 342.600 463.050 343.050 ;
        RECT 493.950 342.600 496.050 343.050 ;
        RECT 460.950 341.400 496.050 342.600 ;
        RECT 460.950 340.950 463.050 341.400 ;
        RECT 493.950 340.950 496.050 341.400 ;
        RECT 709.950 342.600 712.050 343.050 ;
        RECT 715.950 342.600 718.050 343.050 ;
        RECT 709.950 341.400 718.050 342.600 ;
        RECT 709.950 340.950 712.050 341.400 ;
        RECT 715.950 340.950 718.050 341.400 ;
        RECT 739.950 342.600 742.050 343.050 ;
        RECT 748.950 342.600 751.050 343.050 ;
        RECT 739.950 341.400 751.050 342.600 ;
        RECT 739.950 340.950 742.050 341.400 ;
        RECT 748.950 340.950 751.050 341.400 ;
        RECT 754.950 342.600 757.050 343.050 ;
        RECT 760.950 342.600 763.050 343.050 ;
        RECT 754.950 341.400 763.050 342.600 ;
        RECT 754.950 340.950 757.050 341.400 ;
        RECT 760.950 340.950 763.050 341.400 ;
        RECT 46.950 339.600 49.050 340.050 ;
        RECT 73.950 339.600 76.050 340.050 ;
        RECT 46.950 338.400 76.050 339.600 ;
        RECT 46.950 337.950 49.050 338.400 ;
        RECT 73.950 337.950 76.050 338.400 ;
        RECT 79.950 339.600 82.050 340.050 ;
        RECT 112.950 339.600 115.050 340.050 ;
        RECT 79.950 338.400 115.050 339.600 ;
        RECT 79.950 337.950 82.050 338.400 ;
        RECT 112.950 337.950 115.050 338.400 ;
        RECT 202.950 339.600 205.050 340.050 ;
        RECT 241.950 339.600 244.050 340.050 ;
        RECT 202.950 338.400 244.050 339.600 ;
        RECT 202.950 337.950 205.050 338.400 ;
        RECT 241.950 337.950 244.050 338.400 ;
        RECT 403.950 339.600 406.050 340.050 ;
        RECT 409.950 339.600 412.050 340.050 ;
        RECT 403.950 338.400 412.050 339.600 ;
        RECT 403.950 337.950 406.050 338.400 ;
        RECT 409.950 337.950 412.050 338.400 ;
        RECT 421.950 337.950 424.050 340.050 ;
        RECT 439.950 339.600 442.050 340.050 ;
        RECT 484.950 339.600 487.050 340.050 ;
        RECT 439.950 338.400 487.050 339.600 ;
        RECT 439.950 337.950 442.050 338.400 ;
        RECT 484.950 337.950 487.050 338.400 ;
        RECT 490.950 339.600 493.050 340.050 ;
        RECT 511.950 339.600 514.050 340.050 ;
        RECT 490.950 338.400 514.050 339.600 ;
        RECT 490.950 337.950 493.050 338.400 ;
        RECT 511.950 337.950 514.050 338.400 ;
        RECT 529.950 339.600 532.050 340.050 ;
        RECT 571.950 339.600 574.050 340.050 ;
        RECT 529.950 338.400 574.050 339.600 ;
        RECT 529.950 337.950 532.050 338.400 ;
        RECT 571.950 337.950 574.050 338.400 ;
        RECT 646.950 339.600 649.050 340.050 ;
        RECT 658.950 339.600 661.050 340.050 ;
        RECT 646.950 338.400 661.050 339.600 ;
        RECT 646.950 337.950 649.050 338.400 ;
        RECT 658.950 337.950 661.050 338.400 ;
        RECT 730.950 339.600 733.050 340.050 ;
        RECT 751.950 339.600 754.050 340.050 ;
        RECT 730.950 338.400 754.050 339.600 ;
        RECT 730.950 337.950 733.050 338.400 ;
        RECT 751.950 337.950 754.050 338.400 ;
        RECT 34.950 336.600 37.050 337.050 ;
        RECT 70.950 336.600 73.050 337.050 ;
        RECT 79.950 336.600 82.050 337.050 ;
        RECT 34.950 335.400 82.050 336.600 ;
        RECT 34.950 334.950 37.050 335.400 ;
        RECT 70.950 334.950 73.050 335.400 ;
        RECT 79.950 334.950 82.050 335.400 ;
        RECT 85.950 336.600 88.050 337.050 ;
        RECT 118.950 336.600 121.050 337.050 ;
        RECT 85.950 335.400 121.050 336.600 ;
        RECT 85.950 334.950 88.050 335.400 ;
        RECT 118.950 334.950 121.050 335.400 ;
        RECT 238.950 336.600 241.050 337.050 ;
        RECT 268.950 336.600 271.050 337.050 ;
        RECT 238.950 335.400 271.050 336.600 ;
        RECT 238.950 334.950 241.050 335.400 ;
        RECT 268.950 334.950 271.050 335.400 ;
        RECT 340.950 336.600 343.050 337.050 ;
        RECT 370.950 336.600 373.050 337.050 ;
        RECT 422.400 336.600 423.600 337.950 ;
        RECT 439.950 336.600 442.050 337.050 ;
        RECT 340.950 335.400 442.050 336.600 ;
        RECT 340.950 334.950 343.050 335.400 ;
        RECT 370.950 334.950 373.050 335.400 ;
        RECT 439.950 334.950 442.050 335.400 ;
        RECT 496.950 336.600 499.050 337.050 ;
        RECT 565.950 336.600 568.050 337.050 ;
        RECT 739.950 336.600 742.050 337.050 ;
        RECT 496.950 335.400 742.050 336.600 ;
        RECT 496.950 334.950 499.050 335.400 ;
        RECT 565.950 334.950 568.050 335.400 ;
        RECT 739.950 334.950 742.050 335.400 ;
        RECT 304.950 333.600 307.050 334.050 ;
        RECT 322.950 333.600 325.050 334.050 ;
        RECT 304.950 332.400 325.050 333.600 ;
        RECT 304.950 331.950 307.050 332.400 ;
        RECT 322.950 331.950 325.050 332.400 ;
        RECT 112.950 321.600 115.050 322.050 ;
        RECT 313.950 321.600 316.050 322.050 ;
        RECT 328.950 321.600 331.050 322.050 ;
        RECT 478.950 321.600 481.050 322.050 ;
        RECT 520.950 321.600 523.050 322.050 ;
        RECT 112.950 320.400 523.050 321.600 ;
        RECT 112.950 319.950 115.050 320.400 ;
        RECT 313.950 319.950 316.050 320.400 ;
        RECT 328.950 319.950 331.050 320.400 ;
        RECT 478.950 319.950 481.050 320.400 ;
        RECT 520.950 319.950 523.050 320.400 ;
        RECT 325.950 318.600 328.050 319.050 ;
        RECT 334.950 318.600 337.050 319.050 ;
        RECT 364.950 318.600 367.050 319.050 ;
        RECT 325.950 317.400 367.050 318.600 ;
        RECT 325.950 316.950 328.050 317.400 ;
        RECT 334.950 316.950 337.050 317.400 ;
        RECT 364.950 316.950 367.050 317.400 ;
        RECT 64.950 315.600 67.050 316.050 ;
        RECT 76.950 315.600 79.050 316.050 ;
        RECT 64.950 314.400 79.050 315.600 ;
        RECT 64.950 313.950 67.050 314.400 ;
        RECT 76.950 313.950 79.050 314.400 ;
        RECT 136.950 315.600 139.050 316.050 ;
        RECT 193.950 315.600 196.050 316.050 ;
        RECT 136.950 314.400 196.050 315.600 ;
        RECT 136.950 313.950 139.050 314.400 ;
        RECT 193.950 313.950 196.050 314.400 ;
        RECT 196.950 315.600 199.050 316.050 ;
        RECT 226.950 315.600 229.050 316.050 ;
        RECT 196.950 314.400 229.050 315.600 ;
        RECT 196.950 313.950 199.050 314.400 ;
        RECT 226.950 313.950 229.050 314.400 ;
        RECT 304.950 315.600 307.050 316.050 ;
        RECT 442.950 315.600 445.050 316.050 ;
        RECT 304.950 314.400 445.050 315.600 ;
        RECT 304.950 313.950 307.050 314.400 ;
        RECT 442.950 313.950 445.050 314.400 ;
        RECT 652.950 315.600 655.050 316.050 ;
        RECT 664.950 315.600 667.050 316.050 ;
        RECT 673.950 315.600 676.050 316.050 ;
        RECT 652.950 314.400 676.050 315.600 ;
        RECT 652.950 313.950 655.050 314.400 ;
        RECT 664.950 313.950 667.050 314.400 ;
        RECT 673.950 313.950 676.050 314.400 ;
        RECT 112.950 312.600 115.050 313.050 ;
        RECT 133.950 312.600 136.050 313.050 ;
        RECT 112.950 311.400 136.050 312.600 ;
        RECT 112.950 310.950 115.050 311.400 ;
        RECT 133.950 310.950 136.050 311.400 ;
        RECT 244.950 312.600 247.050 313.050 ;
        RECT 253.950 312.600 256.050 313.050 ;
        RECT 274.950 312.600 277.050 313.050 ;
        RECT 244.950 311.400 277.050 312.600 ;
        RECT 244.950 310.950 247.050 311.400 ;
        RECT 253.950 310.950 256.050 311.400 ;
        RECT 274.950 310.950 277.050 311.400 ;
        RECT 406.950 310.950 409.050 313.050 ;
        RECT 625.950 312.600 628.050 313.050 ;
        RECT 652.950 312.600 655.050 313.050 ;
        RECT 625.950 311.400 655.050 312.600 ;
        RECT 625.950 310.950 628.050 311.400 ;
        RECT 652.950 310.950 655.050 311.400 ;
        RECT 658.950 312.600 661.050 313.050 ;
        RECT 667.950 312.600 670.050 313.050 ;
        RECT 658.950 311.400 670.050 312.600 ;
        RECT 658.950 310.950 661.050 311.400 ;
        RECT 667.950 310.950 670.050 311.400 ;
        RECT 685.950 312.600 688.050 313.050 ;
        RECT 703.950 312.600 706.050 313.050 ;
        RECT 685.950 311.400 706.050 312.600 ;
        RECT 685.950 310.950 688.050 311.400 ;
        RECT 703.950 310.950 706.050 311.400 ;
        RECT 40.950 309.600 43.050 310.050 ;
        RECT 52.950 309.600 55.050 310.050 ;
        RECT 73.950 309.600 76.050 310.050 ;
        RECT 40.950 308.400 76.050 309.600 ;
        RECT 40.950 307.950 43.050 308.400 ;
        RECT 52.950 307.950 55.050 308.400 ;
        RECT 73.950 307.950 76.050 308.400 ;
        RECT 325.950 309.600 328.050 310.050 ;
        RECT 361.950 309.600 364.050 310.050 ;
        RECT 397.950 309.600 400.050 310.050 ;
        RECT 325.950 308.400 400.050 309.600 ;
        RECT 407.400 309.600 408.600 310.950 ;
        RECT 442.950 309.600 445.050 310.050 ;
        RECT 481.950 309.600 484.050 310.050 ;
        RECT 407.400 308.400 484.050 309.600 ;
        RECT 325.950 307.950 328.050 308.400 ;
        RECT 361.950 307.950 364.050 308.400 ;
        RECT 397.950 307.950 400.050 308.400 ;
        RECT 442.950 307.950 445.050 308.400 ;
        RECT 481.950 307.950 484.050 308.400 ;
        RECT 487.950 309.600 490.050 310.050 ;
        RECT 526.950 309.600 529.050 310.050 ;
        RECT 487.950 308.400 529.050 309.600 ;
        RECT 487.950 307.950 490.050 308.400 ;
        RECT 526.950 307.950 529.050 308.400 ;
        RECT 631.950 309.600 634.050 310.050 ;
        RECT 643.950 309.600 646.050 310.050 ;
        RECT 631.950 308.400 646.050 309.600 ;
        RECT 631.950 307.950 634.050 308.400 ;
        RECT 643.950 307.950 646.050 308.400 ;
        RECT 196.950 306.600 199.050 307.050 ;
        RECT 232.950 306.600 235.050 307.050 ;
        RECT 244.950 306.600 247.050 307.050 ;
        RECT 196.950 305.400 247.050 306.600 ;
        RECT 196.950 304.950 199.050 305.400 ;
        RECT 232.950 304.950 235.050 305.400 ;
        RECT 244.950 304.950 247.050 305.400 ;
        RECT 250.950 306.600 253.050 307.050 ;
        RECT 370.950 306.600 373.050 307.050 ;
        RECT 403.950 306.600 406.050 307.050 ;
        RECT 250.950 305.400 406.050 306.600 ;
        RECT 250.950 304.950 253.050 305.400 ;
        RECT 370.950 304.950 373.050 305.400 ;
        RECT 403.950 304.950 406.050 305.400 ;
        RECT 727.950 306.600 730.050 307.050 ;
        RECT 742.950 306.600 745.050 307.050 ;
        RECT 727.950 305.400 745.050 306.600 ;
        RECT 727.950 304.950 730.050 305.400 ;
        RECT 742.950 304.950 745.050 305.400 ;
        RECT 643.950 303.600 646.050 304.050 ;
        RECT 649.950 303.600 652.050 304.050 ;
        RECT 643.950 302.400 652.050 303.600 ;
        RECT 643.950 301.950 646.050 302.400 ;
        RECT 649.950 301.950 652.050 302.400 ;
        RECT 31.950 300.600 34.050 301.050 ;
        RECT 358.950 300.600 361.050 301.050 ;
        RECT 31.950 299.400 361.050 300.600 ;
        RECT 31.950 298.950 34.050 299.400 ;
        RECT 358.950 298.950 361.050 299.400 ;
        RECT 154.950 297.600 157.050 298.050 ;
        RECT 202.950 297.600 205.050 298.050 ;
        RECT 154.950 296.400 205.050 297.600 ;
        RECT 154.950 295.950 157.050 296.400 ;
        RECT 202.950 295.950 205.050 296.400 ;
        RECT 238.950 282.600 241.050 283.050 ;
        RECT 268.950 282.600 271.050 283.050 ;
        RECT 274.950 282.600 277.050 283.050 ;
        RECT 238.950 281.400 277.050 282.600 ;
        RECT 238.950 280.950 241.050 281.400 ;
        RECT 268.950 280.950 271.050 281.400 ;
        RECT 274.950 280.950 277.050 281.400 ;
        RECT 409.950 279.600 412.050 280.050 ;
        RECT 577.950 279.600 580.050 280.050 ;
        RECT 409.950 278.400 580.050 279.600 ;
        RECT 409.950 277.950 412.050 278.400 ;
        RECT 577.950 277.950 580.050 278.400 ;
        RECT 514.950 276.600 517.050 277.050 ;
        RECT 535.950 276.600 538.050 277.050 ;
        RECT 514.950 275.400 538.050 276.600 ;
        RECT 514.950 274.950 517.050 275.400 ;
        RECT 535.950 274.950 538.050 275.400 ;
        RECT 127.950 273.600 130.050 274.050 ;
        RECT 193.950 273.600 196.050 274.050 ;
        RECT 127.950 272.400 196.050 273.600 ;
        RECT 127.950 271.950 130.050 272.400 ;
        RECT 193.950 271.950 196.050 272.400 ;
        RECT 199.950 273.600 202.050 274.050 ;
        RECT 313.950 273.600 316.050 274.050 ;
        RECT 322.950 273.600 325.050 274.050 ;
        RECT 199.950 272.400 285.600 273.600 ;
        RECT 199.950 271.950 202.050 272.400 ;
        RECT 284.400 271.050 285.600 272.400 ;
        RECT 313.950 272.400 325.050 273.600 ;
        RECT 313.950 271.950 316.050 272.400 ;
        RECT 322.950 271.950 325.050 272.400 ;
        RECT 421.950 273.600 424.050 274.050 ;
        RECT 445.950 273.600 448.050 274.050 ;
        RECT 478.950 273.600 481.050 274.050 ;
        RECT 421.950 272.400 481.050 273.600 ;
        RECT 421.950 271.950 424.050 272.400 ;
        RECT 445.950 271.950 448.050 272.400 ;
        RECT 478.950 271.950 481.050 272.400 ;
        RECT 490.950 273.600 493.050 274.050 ;
        RECT 529.950 273.600 532.050 274.050 ;
        RECT 490.950 272.400 532.050 273.600 ;
        RECT 490.950 271.950 493.050 272.400 ;
        RECT 529.950 271.950 532.050 272.400 ;
        RECT 622.950 273.600 625.050 274.050 ;
        RECT 697.950 273.600 700.050 274.050 ;
        RECT 706.950 273.600 709.050 274.050 ;
        RECT 622.950 272.400 709.050 273.600 ;
        RECT 622.950 271.950 625.050 272.400 ;
        RECT 697.950 271.950 700.050 272.400 ;
        RECT 706.950 271.950 709.050 272.400 ;
        RECT 37.950 270.600 40.050 271.050 ;
        RECT 49.950 270.600 52.050 271.050 ;
        RECT 76.950 270.600 79.050 271.050 ;
        RECT 37.950 269.400 79.050 270.600 ;
        RECT 37.950 268.950 40.050 269.400 ;
        RECT 49.950 268.950 52.050 269.400 ;
        RECT 76.950 268.950 79.050 269.400 ;
        RECT 157.950 270.600 160.050 271.050 ;
        RECT 190.950 270.600 193.050 271.050 ;
        RECT 157.950 269.400 193.050 270.600 ;
        RECT 157.950 268.950 160.050 269.400 ;
        RECT 190.950 268.950 193.050 269.400 ;
        RECT 196.950 270.600 199.050 271.050 ;
        RECT 202.950 270.600 205.050 271.050 ;
        RECT 238.950 270.600 241.050 271.050 ;
        RECT 196.950 269.400 241.050 270.600 ;
        RECT 196.950 268.950 199.050 269.400 ;
        RECT 202.950 268.950 205.050 269.400 ;
        RECT 238.950 268.950 241.050 269.400 ;
        RECT 283.950 268.950 286.050 271.050 ;
        RECT 316.950 270.600 319.050 271.050 ;
        RECT 325.950 270.600 328.050 271.050 ;
        RECT 316.950 269.400 328.050 270.600 ;
        RECT 316.950 268.950 319.050 269.400 ;
        RECT 325.950 268.950 328.050 269.400 ;
        RECT 358.950 270.600 361.050 271.050 ;
        RECT 400.950 270.600 403.050 271.050 ;
        RECT 358.950 269.400 403.050 270.600 ;
        RECT 358.950 268.950 361.050 269.400 ;
        RECT 400.950 268.950 403.050 269.400 ;
        RECT 406.950 270.600 409.050 271.050 ;
        RECT 412.950 270.600 415.050 271.050 ;
        RECT 406.950 269.400 415.050 270.600 ;
        RECT 406.950 268.950 409.050 269.400 ;
        RECT 412.950 268.950 415.050 269.400 ;
        RECT 448.950 270.600 451.050 271.050 ;
        RECT 514.950 270.600 517.050 271.050 ;
        RECT 448.950 269.400 517.050 270.600 ;
        RECT 448.950 268.950 451.050 269.400 ;
        RECT 514.950 268.950 517.050 269.400 ;
        RECT 517.950 270.600 520.050 271.050 ;
        RECT 532.950 270.600 535.050 271.050 ;
        RECT 517.950 269.400 535.050 270.600 ;
        RECT 517.950 268.950 520.050 269.400 ;
        RECT 532.950 268.950 535.050 269.400 ;
        RECT 625.950 270.600 628.050 271.050 ;
        RECT 652.950 270.600 655.050 271.050 ;
        RECT 625.950 269.400 655.050 270.600 ;
        RECT 625.950 268.950 628.050 269.400 ;
        RECT 652.950 268.950 655.050 269.400 ;
        RECT 658.950 270.600 661.050 271.050 ;
        RECT 700.950 270.600 703.050 271.050 ;
        RECT 658.950 269.400 703.050 270.600 ;
        RECT 658.950 268.950 661.050 269.400 ;
        RECT 700.950 268.950 703.050 269.400 ;
        RECT 40.950 267.600 43.050 268.050 ;
        RECT 46.950 267.600 49.050 268.050 ;
        RECT 70.950 267.600 73.050 268.050 ;
        RECT 73.950 267.600 76.050 268.050 ;
        RECT 40.950 266.400 76.050 267.600 ;
        RECT 40.950 265.950 43.050 266.400 ;
        RECT 46.950 265.950 49.050 266.400 ;
        RECT 70.950 265.950 73.050 266.400 ;
        RECT 73.950 265.950 76.050 266.400 ;
        RECT 82.950 267.600 85.050 268.050 ;
        RECT 118.950 267.600 121.050 268.050 ;
        RECT 367.950 267.600 370.050 268.050 ;
        RECT 454.950 267.600 457.050 268.050 ;
        RECT 484.950 267.600 487.050 268.050 ;
        RECT 82.950 266.400 487.050 267.600 ;
        RECT 82.950 265.950 85.050 266.400 ;
        RECT 118.950 265.950 121.050 266.400 ;
        RECT 367.950 265.950 370.050 266.400 ;
        RECT 454.950 265.950 457.050 266.400 ;
        RECT 484.950 265.950 487.050 266.400 ;
        RECT 580.950 267.600 583.050 268.050 ;
        RECT 607.950 267.600 610.050 268.050 ;
        RECT 580.950 266.400 610.050 267.600 ;
        RECT 580.950 265.950 583.050 266.400 ;
        RECT 607.950 265.950 610.050 266.400 ;
        RECT 655.950 267.600 658.050 268.050 ;
        RECT 661.950 267.600 664.050 268.050 ;
        RECT 655.950 266.400 664.050 267.600 ;
        RECT 655.950 265.950 658.050 266.400 ;
        RECT 661.950 265.950 664.050 266.400 ;
        RECT 664.950 267.600 667.050 268.050 ;
        RECT 724.950 267.600 727.050 268.050 ;
        RECT 664.950 266.400 727.050 267.600 ;
        RECT 664.950 265.950 667.050 266.400 ;
        RECT 724.950 265.950 727.050 266.400 ;
        RECT 736.950 267.600 739.050 268.050 ;
        RECT 745.950 267.600 748.050 268.050 ;
        RECT 736.950 266.400 748.050 267.600 ;
        RECT 736.950 265.950 739.050 266.400 ;
        RECT 745.950 265.950 748.050 266.400 ;
        RECT 16.950 264.600 19.050 265.050 ;
        RECT 37.950 264.600 40.050 265.050 ;
        RECT 16.950 263.400 40.050 264.600 ;
        RECT 16.950 262.950 19.050 263.400 ;
        RECT 37.950 262.950 40.050 263.400 ;
        RECT 199.950 264.600 202.050 265.050 ;
        RECT 280.950 264.600 283.050 265.050 ;
        RECT 199.950 263.400 283.050 264.600 ;
        RECT 199.950 262.950 202.050 263.400 ;
        RECT 280.950 262.950 283.050 263.400 ;
        RECT 289.950 264.600 292.050 265.050 ;
        RECT 571.950 264.600 574.050 265.050 ;
        RECT 289.950 263.400 574.050 264.600 ;
        RECT 289.950 262.950 292.050 263.400 ;
        RECT 571.950 262.950 574.050 263.400 ;
        RECT 574.950 264.600 577.050 265.050 ;
        RECT 595.950 264.600 598.050 265.050 ;
        RECT 574.950 263.400 598.050 264.600 ;
        RECT 574.950 262.950 577.050 263.400 ;
        RECT 595.950 262.950 598.050 263.400 ;
        RECT 601.950 264.600 604.050 265.050 ;
        RECT 664.950 264.600 667.050 265.050 ;
        RECT 601.950 263.400 667.050 264.600 ;
        RECT 601.950 262.950 604.050 263.400 ;
        RECT 664.950 262.950 667.050 263.400 ;
        RECT 82.950 261.600 85.050 262.050 ;
        RECT 100.950 261.600 103.050 262.050 ;
        RECT 82.950 260.400 103.050 261.600 ;
        RECT 82.950 259.950 85.050 260.400 ;
        RECT 100.950 259.950 103.050 260.400 ;
        RECT 712.950 255.600 715.050 256.050 ;
        RECT 718.950 255.600 721.050 256.050 ;
        RECT 712.950 254.400 721.050 255.600 ;
        RECT 712.950 253.950 715.050 254.400 ;
        RECT 718.950 253.950 721.050 254.400 ;
        RECT 154.950 249.600 157.050 250.050 ;
        RECT 208.950 249.600 211.050 250.050 ;
        RECT 154.950 248.400 211.050 249.600 ;
        RECT 154.950 247.950 157.050 248.400 ;
        RECT 208.950 247.950 211.050 248.400 ;
        RECT 121.950 246.600 124.050 247.050 ;
        RECT 220.950 246.600 223.050 247.050 ;
        RECT 286.950 246.600 289.050 247.050 ;
        RECT 367.950 246.600 370.050 247.050 ;
        RECT 121.950 245.400 370.050 246.600 ;
        RECT 121.950 244.950 124.050 245.400 ;
        RECT 220.950 244.950 223.050 245.400 ;
        RECT 286.950 244.950 289.050 245.400 ;
        RECT 367.950 244.950 370.050 245.400 ;
        RECT 160.950 243.600 163.050 244.050 ;
        RECT 253.950 243.600 256.050 244.050 ;
        RECT 160.950 242.400 256.050 243.600 ;
        RECT 160.950 241.950 163.050 242.400 ;
        RECT 253.950 241.950 256.050 242.400 ;
        RECT 370.950 243.600 373.050 244.050 ;
        RECT 427.950 243.600 430.050 244.050 ;
        RECT 445.950 243.600 448.050 244.050 ;
        RECT 370.950 242.400 448.050 243.600 ;
        RECT 370.950 241.950 373.050 242.400 ;
        RECT 427.950 241.950 430.050 242.400 ;
        RECT 445.950 241.950 448.050 242.400 ;
        RECT 547.950 243.600 550.050 244.050 ;
        RECT 568.950 243.600 571.050 244.050 ;
        RECT 547.950 242.400 571.050 243.600 ;
        RECT 547.950 241.950 550.050 242.400 ;
        RECT 568.950 241.950 571.050 242.400 ;
        RECT 586.950 243.600 589.050 244.050 ;
        RECT 625.950 243.600 628.050 244.050 ;
        RECT 586.950 242.400 628.050 243.600 ;
        RECT 586.950 241.950 589.050 242.400 ;
        RECT 625.950 241.950 628.050 242.400 ;
        RECT 43.950 240.600 46.050 241.050 ;
        RECT 67.950 240.600 70.050 241.050 ;
        RECT 43.950 239.400 70.050 240.600 ;
        RECT 43.950 238.950 46.050 239.400 ;
        RECT 67.950 238.950 70.050 239.400 ;
        RECT 88.950 240.600 91.050 241.050 ;
        RECT 103.950 240.600 106.050 241.050 ;
        RECT 88.950 239.400 106.050 240.600 ;
        RECT 88.950 238.950 91.050 239.400 ;
        RECT 103.950 238.950 106.050 239.400 ;
        RECT 133.950 240.600 136.050 241.050 ;
        RECT 211.950 240.600 214.050 241.050 ;
        RECT 229.950 240.600 232.050 241.050 ;
        RECT 133.950 239.400 232.050 240.600 ;
        RECT 133.950 238.950 136.050 239.400 ;
        RECT 211.950 238.950 214.050 239.400 ;
        RECT 229.950 238.950 232.050 239.400 ;
        RECT 292.950 240.600 295.050 241.050 ;
        RECT 322.950 240.600 325.050 241.050 ;
        RECT 334.950 240.600 337.050 241.050 ;
        RECT 292.950 239.400 337.050 240.600 ;
        RECT 292.950 238.950 295.050 239.400 ;
        RECT 322.950 238.950 325.050 239.400 ;
        RECT 334.950 238.950 337.050 239.400 ;
        RECT 337.950 240.600 340.050 241.050 ;
        RECT 343.950 240.600 346.050 241.050 ;
        RECT 337.950 239.400 346.050 240.600 ;
        RECT 337.950 238.950 340.050 239.400 ;
        RECT 343.950 238.950 346.050 239.400 ;
        RECT 376.950 240.600 379.050 241.050 ;
        RECT 412.950 240.600 415.050 241.050 ;
        RECT 463.950 240.600 466.050 241.050 ;
        RECT 517.950 240.600 520.050 241.050 ;
        RECT 376.950 239.400 411.600 240.600 ;
        RECT 376.950 238.950 379.050 239.400 ;
        RECT 40.950 237.600 43.050 238.050 ;
        RECT 52.950 237.600 55.050 238.050 ;
        RECT 85.950 237.600 88.050 238.050 ;
        RECT 40.950 236.400 88.050 237.600 ;
        RECT 40.950 235.950 43.050 236.400 ;
        RECT 52.950 235.950 55.050 236.400 ;
        RECT 85.950 235.950 88.050 236.400 ;
        RECT 205.950 235.950 208.050 238.050 ;
        RECT 247.950 237.600 250.050 238.050 ;
        RECT 265.950 237.600 268.050 238.050 ;
        RECT 289.950 237.600 292.050 238.050 ;
        RECT 325.950 237.600 328.050 238.050 ;
        RECT 247.950 236.400 328.050 237.600 ;
        RECT 410.400 237.600 411.600 239.400 ;
        RECT 412.950 239.400 466.050 240.600 ;
        RECT 412.950 238.950 415.050 239.400 ;
        RECT 463.950 238.950 466.050 239.400 ;
        RECT 509.400 239.400 520.050 240.600 ;
        RECT 509.400 237.600 510.600 239.400 ;
        RECT 517.950 238.950 520.050 239.400 ;
        RECT 592.950 240.600 595.050 241.050 ;
        RECT 652.950 240.600 655.050 241.050 ;
        RECT 592.950 239.400 655.050 240.600 ;
        RECT 592.950 238.950 595.050 239.400 ;
        RECT 652.950 238.950 655.050 239.400 ;
        RECT 658.950 240.600 661.050 241.050 ;
        RECT 664.950 240.600 667.050 241.050 ;
        RECT 658.950 239.400 667.050 240.600 ;
        RECT 658.950 238.950 661.050 239.400 ;
        RECT 664.950 238.950 667.050 239.400 ;
        RECT 670.950 240.600 673.050 241.050 ;
        RECT 721.950 240.600 724.050 241.050 ;
        RECT 670.950 239.400 724.050 240.600 ;
        RECT 670.950 238.950 673.050 239.400 ;
        RECT 721.950 238.950 724.050 239.400 ;
        RECT 410.400 236.400 510.600 237.600 ;
        RECT 511.950 237.600 514.050 238.050 ;
        RECT 589.950 237.600 592.050 238.050 ;
        RECT 511.950 236.400 592.050 237.600 ;
        RECT 247.950 235.950 250.050 236.400 ;
        RECT 265.950 235.950 268.050 236.400 ;
        RECT 289.950 235.950 292.050 236.400 ;
        RECT 325.950 235.950 328.050 236.400 ;
        RECT 511.950 235.950 514.050 236.400 ;
        RECT 589.950 235.950 592.050 236.400 ;
        RECT 595.950 237.600 598.050 238.050 ;
        RECT 634.950 237.600 637.050 238.050 ;
        RECT 595.950 236.400 637.050 237.600 ;
        RECT 595.950 235.950 598.050 236.400 ;
        RECT 634.950 235.950 637.050 236.400 ;
        RECT 715.950 237.600 718.050 238.050 ;
        RECT 751.950 237.600 754.050 238.050 ;
        RECT 715.950 236.400 754.050 237.600 ;
        RECT 715.950 235.950 718.050 236.400 ;
        RECT 751.950 235.950 754.050 236.400 ;
        RECT 124.950 234.600 127.050 235.050 ;
        RECT 169.950 234.600 172.050 235.050 ;
        RECT 124.950 233.400 172.050 234.600 ;
        RECT 206.400 234.600 207.600 235.950 ;
        RECT 244.950 234.600 247.050 235.050 ;
        RECT 206.400 233.400 247.050 234.600 ;
        RECT 124.950 232.950 127.050 233.400 ;
        RECT 169.950 232.950 172.050 233.400 ;
        RECT 244.950 232.950 247.050 233.400 ;
        RECT 250.950 234.600 253.050 235.050 ;
        RECT 259.950 234.600 262.050 235.050 ;
        RECT 250.950 233.400 262.050 234.600 ;
        RECT 250.950 232.950 253.050 233.400 ;
        RECT 259.950 232.950 262.050 233.400 ;
        RECT 331.950 234.600 334.050 235.050 ;
        RECT 349.950 234.600 352.050 235.050 ;
        RECT 364.950 234.600 367.050 235.050 ;
        RECT 331.950 233.400 367.050 234.600 ;
        RECT 331.950 232.950 334.050 233.400 ;
        RECT 349.950 232.950 352.050 233.400 ;
        RECT 364.950 232.950 367.050 233.400 ;
        RECT 412.950 234.600 415.050 235.050 ;
        RECT 424.950 234.600 427.050 235.050 ;
        RECT 412.950 233.400 427.050 234.600 ;
        RECT 412.950 232.950 415.050 233.400 ;
        RECT 424.950 232.950 427.050 233.400 ;
        RECT 469.950 234.600 472.050 235.050 ;
        RECT 508.950 234.600 511.050 235.050 ;
        RECT 469.950 233.400 511.050 234.600 ;
        RECT 469.950 232.950 472.050 233.400 ;
        RECT 508.950 232.950 511.050 233.400 ;
        RECT 625.950 234.600 628.050 235.050 ;
        RECT 631.950 234.600 634.050 235.050 ;
        RECT 625.950 233.400 634.050 234.600 ;
        RECT 625.950 232.950 628.050 233.400 ;
        RECT 631.950 232.950 634.050 233.400 ;
        RECT 637.950 234.600 640.050 235.050 ;
        RECT 670.950 234.600 673.050 235.050 ;
        RECT 637.950 233.400 673.050 234.600 ;
        RECT 637.950 232.950 640.050 233.400 ;
        RECT 670.950 232.950 673.050 233.400 ;
        RECT 703.950 234.600 706.050 235.050 ;
        RECT 754.950 234.600 757.050 235.050 ;
        RECT 703.950 233.400 757.050 234.600 ;
        RECT 703.950 232.950 706.050 233.400 ;
        RECT 754.950 232.950 757.050 233.400 ;
        RECT 415.950 231.600 418.050 232.050 ;
        RECT 457.950 231.600 460.050 232.050 ;
        RECT 415.950 230.400 460.050 231.600 ;
        RECT 415.950 229.950 418.050 230.400 ;
        RECT 457.950 229.950 460.050 230.400 ;
        RECT 550.950 231.600 553.050 232.050 ;
        RECT 574.950 231.600 577.050 232.050 ;
        RECT 649.950 231.600 652.050 232.050 ;
        RECT 550.950 230.400 652.050 231.600 ;
        RECT 550.950 229.950 553.050 230.400 ;
        RECT 574.950 229.950 577.050 230.400 ;
        RECT 649.950 229.950 652.050 230.400 ;
        RECT 547.950 228.600 550.050 229.050 ;
        RECT 709.950 228.600 712.050 229.050 ;
        RECT 547.950 227.400 712.050 228.600 ;
        RECT 547.950 226.950 550.050 227.400 ;
        RECT 709.950 226.950 712.050 227.400 ;
        RECT 451.950 204.600 454.050 205.050 ;
        RECT 511.950 204.600 514.050 205.050 ;
        RECT 451.950 203.400 514.050 204.600 ;
        RECT 451.950 202.950 454.050 203.400 ;
        RECT 511.950 202.950 514.050 203.400 ;
        RECT 625.950 204.600 628.050 205.050 ;
        RECT 637.950 204.600 640.050 205.050 ;
        RECT 625.950 203.400 640.050 204.600 ;
        RECT 625.950 202.950 628.050 203.400 ;
        RECT 637.950 202.950 640.050 203.400 ;
        RECT 61.950 201.600 64.050 202.050 ;
        RECT 85.950 201.600 88.050 202.050 ;
        RECT 94.950 201.600 97.050 202.050 ;
        RECT 61.950 200.400 97.050 201.600 ;
        RECT 61.950 199.950 64.050 200.400 ;
        RECT 85.950 199.950 88.050 200.400 ;
        RECT 94.950 199.950 97.050 200.400 ;
        RECT 100.950 201.600 103.050 202.050 ;
        RECT 124.950 201.600 127.050 202.050 ;
        RECT 100.950 200.400 127.050 201.600 ;
        RECT 100.950 199.950 103.050 200.400 ;
        RECT 124.950 199.950 127.050 200.400 ;
        RECT 127.950 201.600 130.050 202.050 ;
        RECT 154.950 201.600 157.050 202.050 ;
        RECT 127.950 200.400 157.050 201.600 ;
        RECT 127.950 199.950 130.050 200.400 ;
        RECT 154.950 199.950 157.050 200.400 ;
        RECT 166.950 201.600 169.050 202.050 ;
        RECT 178.950 201.600 181.050 202.050 ;
        RECT 166.950 200.400 181.050 201.600 ;
        RECT 166.950 199.950 169.050 200.400 ;
        RECT 178.950 199.950 181.050 200.400 ;
        RECT 259.950 201.600 262.050 202.050 ;
        RECT 280.950 201.600 283.050 202.050 ;
        RECT 259.950 200.400 283.050 201.600 ;
        RECT 259.950 199.950 262.050 200.400 ;
        RECT 280.950 199.950 283.050 200.400 ;
        RECT 343.950 201.600 346.050 202.050 ;
        RECT 373.950 201.600 376.050 202.050 ;
        RECT 343.950 200.400 376.050 201.600 ;
        RECT 343.950 199.950 346.050 200.400 ;
        RECT 373.950 199.950 376.050 200.400 ;
        RECT 433.950 201.600 436.050 202.050 ;
        RECT 478.950 201.600 481.050 202.050 ;
        RECT 433.950 200.400 481.050 201.600 ;
        RECT 433.950 199.950 436.050 200.400 ;
        RECT 478.950 199.950 481.050 200.400 ;
        RECT 502.950 201.600 505.050 202.050 ;
        RECT 517.950 201.600 520.050 202.050 ;
        RECT 502.950 200.400 520.050 201.600 ;
        RECT 502.950 199.950 505.050 200.400 ;
        RECT 517.950 199.950 520.050 200.400 ;
        RECT 559.950 201.600 562.050 202.050 ;
        RECT 631.950 201.600 634.050 202.050 ;
        RECT 559.950 200.400 634.050 201.600 ;
        RECT 559.950 199.950 562.050 200.400 ;
        RECT 631.950 199.950 634.050 200.400 ;
        RECT 22.950 198.600 25.050 199.050 ;
        RECT 34.950 198.600 37.050 199.050 ;
        RECT 118.950 198.600 121.050 199.050 ;
        RECT 154.950 198.600 157.050 199.050 ;
        RECT 172.950 198.600 175.050 199.050 ;
        RECT 22.950 197.400 54.600 198.600 ;
        RECT 22.950 196.950 25.050 197.400 ;
        RECT 34.950 196.950 37.050 197.400 ;
        RECT 53.400 195.600 54.600 197.400 ;
        RECT 118.950 197.400 126.600 198.600 ;
        RECT 118.950 196.950 121.050 197.400 ;
        RECT 100.950 195.600 103.050 196.050 ;
        RECT 106.950 195.600 109.050 196.050 ;
        RECT 121.950 195.600 124.050 196.050 ;
        RECT 53.400 194.400 124.050 195.600 ;
        RECT 125.400 195.600 126.600 197.400 ;
        RECT 154.950 197.400 175.050 198.600 ;
        RECT 154.950 196.950 157.050 197.400 ;
        RECT 172.950 196.950 175.050 197.400 ;
        RECT 220.950 198.600 223.050 199.050 ;
        RECT 241.950 198.600 244.050 199.050 ;
        RECT 262.950 198.600 265.050 199.050 ;
        RECT 472.950 198.600 475.050 199.050 ;
        RECT 487.950 198.600 490.050 199.050 ;
        RECT 220.950 197.400 265.050 198.600 ;
        RECT 220.950 196.950 223.050 197.400 ;
        RECT 241.950 196.950 244.050 197.400 ;
        RECT 262.950 196.950 265.050 197.400 ;
        RECT 425.400 197.400 490.050 198.600 ;
        RECT 425.400 196.050 426.600 197.400 ;
        RECT 472.950 196.950 475.050 197.400 ;
        RECT 487.950 196.950 490.050 197.400 ;
        RECT 514.950 198.600 517.050 199.050 ;
        RECT 547.950 198.600 550.050 199.050 ;
        RECT 514.950 197.400 550.050 198.600 ;
        RECT 514.950 196.950 517.050 197.400 ;
        RECT 547.950 196.950 550.050 197.400 ;
        RECT 553.950 198.600 556.050 199.050 ;
        RECT 568.950 198.600 571.050 199.050 ;
        RECT 553.950 197.400 571.050 198.600 ;
        RECT 553.950 196.950 556.050 197.400 ;
        RECT 568.950 196.950 571.050 197.400 ;
        RECT 634.950 198.600 637.050 199.050 ;
        RECT 709.950 198.600 712.050 199.050 ;
        RECT 634.950 197.400 712.050 198.600 ;
        RECT 634.950 196.950 637.050 197.400 ;
        RECT 709.950 196.950 712.050 197.400 ;
        RECT 175.950 195.600 178.050 196.050 ;
        RECT 125.400 194.400 178.050 195.600 ;
        RECT 100.950 193.950 103.050 194.400 ;
        RECT 106.950 193.950 109.050 194.400 ;
        RECT 121.950 193.950 124.050 194.400 ;
        RECT 175.950 193.950 178.050 194.400 ;
        RECT 214.950 195.600 217.050 196.050 ;
        RECT 229.950 195.600 232.050 196.050 ;
        RECT 214.950 194.400 232.050 195.600 ;
        RECT 214.950 193.950 217.050 194.400 ;
        RECT 229.950 193.950 232.050 194.400 ;
        RECT 277.950 195.600 280.050 196.050 ;
        RECT 307.950 195.600 310.050 196.050 ;
        RECT 277.950 194.400 310.050 195.600 ;
        RECT 277.950 193.950 280.050 194.400 ;
        RECT 307.950 193.950 310.050 194.400 ;
        RECT 367.950 195.600 370.050 196.050 ;
        RECT 382.950 195.600 385.050 196.050 ;
        RECT 367.950 194.400 385.050 195.600 ;
        RECT 367.950 193.950 370.050 194.400 ;
        RECT 382.950 193.950 385.050 194.400 ;
        RECT 424.950 193.950 427.050 196.050 ;
        RECT 457.950 195.600 460.050 196.050 ;
        RECT 469.950 195.600 472.050 196.050 ;
        RECT 457.950 194.400 472.050 195.600 ;
        RECT 457.950 193.950 460.050 194.400 ;
        RECT 469.950 193.950 472.050 194.400 ;
        RECT 475.950 195.600 478.050 196.050 ;
        RECT 478.950 195.600 481.050 196.050 ;
        RECT 553.950 195.600 556.050 196.050 ;
        RECT 475.950 194.400 556.050 195.600 ;
        RECT 475.950 193.950 478.050 194.400 ;
        RECT 478.950 193.950 481.050 194.400 ;
        RECT 553.950 193.950 556.050 194.400 ;
        RECT 580.950 195.600 583.050 196.050 ;
        RECT 661.950 195.600 664.050 196.050 ;
        RECT 580.950 194.400 664.050 195.600 ;
        RECT 580.950 193.950 583.050 194.400 ;
        RECT 661.950 193.950 664.050 194.400 ;
        RECT 712.950 195.600 715.050 196.050 ;
        RECT 733.950 195.600 736.050 196.050 ;
        RECT 712.950 194.400 736.050 195.600 ;
        RECT 712.950 193.950 715.050 194.400 ;
        RECT 733.950 193.950 736.050 194.400 ;
        RECT 751.950 195.600 754.050 196.050 ;
        RECT 757.950 195.600 760.050 196.050 ;
        RECT 751.950 194.400 760.050 195.600 ;
        RECT 751.950 193.950 754.050 194.400 ;
        RECT 757.950 193.950 760.050 194.400 ;
        RECT 34.950 192.600 37.050 193.050 ;
        RECT 49.950 192.600 52.050 193.050 ;
        RECT 34.950 191.400 52.050 192.600 ;
        RECT 34.950 190.950 37.050 191.400 ;
        RECT 49.950 190.950 52.050 191.400 ;
        RECT 373.950 192.600 376.050 193.050 ;
        RECT 427.950 192.600 430.050 193.050 ;
        RECT 373.950 191.400 430.050 192.600 ;
        RECT 373.950 190.950 376.050 191.400 ;
        RECT 427.950 190.950 430.050 191.400 ;
        RECT 580.950 192.600 583.050 193.050 ;
        RECT 586.950 192.600 589.050 193.050 ;
        RECT 580.950 191.400 589.050 192.600 ;
        RECT 580.950 190.950 583.050 191.400 ;
        RECT 586.950 190.950 589.050 191.400 ;
        RECT 655.950 192.600 658.050 193.050 ;
        RECT 667.950 192.600 670.050 193.050 ;
        RECT 655.950 191.400 670.050 192.600 ;
        RECT 655.950 190.950 658.050 191.400 ;
        RECT 667.950 190.950 670.050 191.400 ;
        RECT 724.950 192.600 727.050 193.050 ;
        RECT 739.950 192.600 742.050 193.050 ;
        RECT 724.950 191.400 742.050 192.600 ;
        RECT 724.950 190.950 727.050 191.400 ;
        RECT 739.950 190.950 742.050 191.400 ;
        RECT 388.950 189.600 391.050 190.050 ;
        RECT 418.950 189.600 421.050 190.050 ;
        RECT 466.950 189.600 469.050 190.050 ;
        RECT 490.950 189.600 493.050 190.050 ;
        RECT 520.950 189.600 523.050 190.050 ;
        RECT 550.950 189.600 553.050 190.050 ;
        RECT 388.950 188.400 553.050 189.600 ;
        RECT 388.950 187.950 391.050 188.400 ;
        RECT 418.950 187.950 421.050 188.400 ;
        RECT 466.950 187.950 469.050 188.400 ;
        RECT 490.950 187.950 493.050 188.400 ;
        RECT 520.950 187.950 523.050 188.400 ;
        RECT 550.950 187.950 553.050 188.400 ;
        RECT 715.950 186.600 718.050 187.050 ;
        RECT 751.950 186.600 754.050 187.050 ;
        RECT 715.950 185.400 754.050 186.600 ;
        RECT 715.950 184.950 718.050 185.400 ;
        RECT 751.950 184.950 754.050 185.400 ;
        RECT 76.950 174.600 79.050 175.050 ;
        RECT 97.950 174.600 100.050 175.050 ;
        RECT 76.950 173.400 100.050 174.600 ;
        RECT 76.950 172.950 79.050 173.400 ;
        RECT 97.950 172.950 100.050 173.400 ;
        RECT 307.950 174.600 310.050 175.050 ;
        RECT 400.950 174.600 403.050 175.050 ;
        RECT 409.950 174.600 412.050 175.050 ;
        RECT 478.950 174.600 481.050 175.050 ;
        RECT 307.950 173.400 481.050 174.600 ;
        RECT 307.950 172.950 310.050 173.400 ;
        RECT 400.950 172.950 403.050 173.400 ;
        RECT 409.950 172.950 412.050 173.400 ;
        RECT 478.950 172.950 481.050 173.400 ;
        RECT 67.950 171.600 70.050 172.050 ;
        RECT 181.950 171.600 184.050 172.050 ;
        RECT 67.950 170.400 184.050 171.600 ;
        RECT 67.950 169.950 70.050 170.400 ;
        RECT 181.950 169.950 184.050 170.400 ;
        RECT 313.950 171.600 316.050 172.050 ;
        RECT 346.950 171.600 349.050 172.050 ;
        RECT 313.950 170.400 349.050 171.600 ;
        RECT 313.950 169.950 316.050 170.400 ;
        RECT 346.950 169.950 349.050 170.400 ;
        RECT 445.950 171.600 448.050 172.050 ;
        RECT 619.950 171.600 622.050 172.050 ;
        RECT 445.950 170.400 622.050 171.600 ;
        RECT 445.950 169.950 448.050 170.400 ;
        RECT 619.950 169.950 622.050 170.400 ;
        RECT 73.950 168.600 76.050 169.050 ;
        RECT 94.950 168.600 97.050 169.050 ;
        RECT 73.950 167.400 97.050 168.600 ;
        RECT 73.950 166.950 76.050 167.400 ;
        RECT 94.950 166.950 97.050 167.400 ;
        RECT 112.950 168.600 115.050 169.050 ;
        RECT 124.950 168.600 127.050 169.050 ;
        RECT 217.950 168.600 220.050 169.050 ;
        RECT 112.950 167.400 220.050 168.600 ;
        RECT 112.950 166.950 115.050 167.400 ;
        RECT 124.950 166.950 127.050 167.400 ;
        RECT 217.950 166.950 220.050 167.400 ;
        RECT 232.950 168.600 235.050 169.050 ;
        RECT 268.950 168.600 271.050 169.050 ;
        RECT 232.950 167.400 271.050 168.600 ;
        RECT 232.950 166.950 235.050 167.400 ;
        RECT 268.950 166.950 271.050 167.400 ;
        RECT 274.950 168.600 277.050 169.050 ;
        RECT 319.950 168.600 322.050 169.050 ;
        RECT 274.950 167.400 322.050 168.600 ;
        RECT 274.950 166.950 277.050 167.400 ;
        RECT 319.950 166.950 322.050 167.400 ;
        RECT 346.950 168.600 349.050 169.050 ;
        RECT 496.950 168.600 499.050 169.050 ;
        RECT 511.950 168.600 514.050 169.050 ;
        RECT 346.950 167.400 514.050 168.600 ;
        RECT 346.950 166.950 349.050 167.400 ;
        RECT 496.950 166.950 499.050 167.400 ;
        RECT 511.950 166.950 514.050 167.400 ;
        RECT 538.950 168.600 541.050 169.050 ;
        RECT 577.950 168.600 580.050 169.050 ;
        RECT 538.950 167.400 580.050 168.600 ;
        RECT 538.950 166.950 541.050 167.400 ;
        RECT 577.950 166.950 580.050 167.400 ;
        RECT 706.950 168.600 709.050 169.050 ;
        RECT 712.950 168.600 715.050 169.050 ;
        RECT 706.950 167.400 715.050 168.600 ;
        RECT 706.950 166.950 709.050 167.400 ;
        RECT 712.950 166.950 715.050 167.400 ;
        RECT 70.950 165.600 73.050 166.050 ;
        RECT 85.950 165.600 88.050 166.050 ;
        RECT 70.950 164.400 88.050 165.600 ;
        RECT 70.950 163.950 73.050 164.400 ;
        RECT 85.950 163.950 88.050 164.400 ;
        RECT 181.950 165.600 184.050 166.050 ;
        RECT 190.950 165.600 193.050 166.050 ;
        RECT 181.950 164.400 193.050 165.600 ;
        RECT 181.950 163.950 184.050 164.400 ;
        RECT 190.950 163.950 193.050 164.400 ;
        RECT 208.950 165.600 211.050 166.050 ;
        RECT 226.950 165.600 229.050 166.050 ;
        RECT 235.950 165.600 238.050 166.050 ;
        RECT 208.950 164.400 238.050 165.600 ;
        RECT 208.950 163.950 211.050 164.400 ;
        RECT 226.950 163.950 229.050 164.400 ;
        RECT 235.950 163.950 238.050 164.400 ;
        RECT 322.950 165.600 325.050 166.050 ;
        RECT 337.950 165.600 340.050 166.050 ;
        RECT 322.950 164.400 340.050 165.600 ;
        RECT 322.950 163.950 325.050 164.400 ;
        RECT 337.950 163.950 340.050 164.400 ;
        RECT 364.950 165.600 367.050 166.050 ;
        RECT 403.950 165.600 406.050 166.050 ;
        RECT 364.950 164.400 406.050 165.600 ;
        RECT 364.950 163.950 367.050 164.400 ;
        RECT 403.950 163.950 406.050 164.400 ;
        RECT 406.950 163.950 409.050 166.050 ;
        RECT 436.950 165.600 439.050 166.050 ;
        RECT 448.950 165.600 451.050 166.050 ;
        RECT 436.950 164.400 451.050 165.600 ;
        RECT 436.950 163.950 439.050 164.400 ;
        RECT 448.950 163.950 451.050 164.400 ;
        RECT 454.950 163.950 457.050 166.050 ;
        RECT 574.950 165.600 577.050 166.050 ;
        RECT 583.950 165.600 586.050 166.050 ;
        RECT 622.950 165.600 625.050 166.050 ;
        RECT 574.950 164.400 625.050 165.600 ;
        RECT 574.950 163.950 577.050 164.400 ;
        RECT 583.950 163.950 586.050 164.400 ;
        RECT 622.950 163.950 625.050 164.400 ;
        RECT 673.950 165.600 676.050 166.050 ;
        RECT 706.950 165.600 709.050 166.050 ;
        RECT 673.950 164.400 709.050 165.600 ;
        RECT 673.950 163.950 676.050 164.400 ;
        RECT 706.950 163.950 709.050 164.400 ;
        RECT 136.950 162.600 139.050 163.050 ;
        RECT 157.950 162.600 160.050 163.050 ;
        RECT 241.950 162.600 244.050 163.050 ;
        RECT 136.950 161.400 244.050 162.600 ;
        RECT 136.950 160.950 139.050 161.400 ;
        RECT 157.950 160.950 160.050 161.400 ;
        RECT 241.950 160.950 244.050 161.400 ;
        RECT 271.950 160.950 274.050 163.050 ;
        RECT 277.950 162.600 280.050 163.050 ;
        RECT 361.950 162.600 364.050 163.050 ;
        RECT 277.950 161.400 364.050 162.600 ;
        RECT 277.950 160.950 280.050 161.400 ;
        RECT 361.950 160.950 364.050 161.400 ;
        RECT 272.400 159.600 273.600 160.950 ;
        RECT 274.950 159.600 277.050 160.050 ;
        RECT 272.400 158.400 277.050 159.600 ;
        RECT 407.400 159.600 408.600 163.950 ;
        RECT 448.950 162.600 451.050 163.050 ;
        RECT 455.400 162.600 456.600 163.950 ;
        RECT 448.950 161.400 456.600 162.600 ;
        RECT 493.950 162.600 496.050 163.050 ;
        RECT 505.950 162.600 508.050 163.050 ;
        RECT 493.950 161.400 508.050 162.600 ;
        RECT 448.950 160.950 451.050 161.400 ;
        RECT 493.950 160.950 496.050 161.400 ;
        RECT 505.950 160.950 508.050 161.400 ;
        RECT 523.950 162.600 526.050 163.050 ;
        RECT 541.950 162.600 544.050 163.050 ;
        RECT 589.950 162.600 592.050 163.050 ;
        RECT 610.950 162.600 613.050 163.050 ;
        RECT 523.950 161.400 613.050 162.600 ;
        RECT 523.950 160.950 526.050 161.400 ;
        RECT 541.950 160.950 544.050 161.400 ;
        RECT 589.950 160.950 592.050 161.400 ;
        RECT 610.950 160.950 613.050 161.400 ;
        RECT 676.950 162.600 679.050 163.050 ;
        RECT 703.950 162.600 706.050 163.050 ;
        RECT 676.950 161.400 706.050 162.600 ;
        RECT 676.950 160.950 679.050 161.400 ;
        RECT 703.950 160.950 706.050 161.400 ;
        RECT 712.950 162.600 715.050 163.050 ;
        RECT 748.950 162.600 751.050 163.050 ;
        RECT 712.950 161.400 751.050 162.600 ;
        RECT 712.950 160.950 715.050 161.400 ;
        RECT 748.950 160.950 751.050 161.400 ;
        RECT 409.950 159.600 412.050 160.050 ;
        RECT 407.400 158.400 412.050 159.600 ;
        RECT 274.950 157.950 277.050 158.400 ;
        RECT 409.950 157.950 412.050 158.400 ;
        RECT 559.950 159.600 562.050 160.050 ;
        RECT 631.950 159.600 634.050 160.050 ;
        RECT 559.950 158.400 634.050 159.600 ;
        RECT 559.950 157.950 562.050 158.400 ;
        RECT 631.950 157.950 634.050 158.400 ;
        RECT 412.950 156.600 415.050 157.050 ;
        RECT 664.950 156.600 667.050 157.050 ;
        RECT 412.950 155.400 667.050 156.600 ;
        RECT 412.950 154.950 415.050 155.400 ;
        RECT 664.950 154.950 667.050 155.400 ;
        RECT 367.950 153.600 370.050 154.050 ;
        RECT 376.950 153.600 379.050 154.050 ;
        RECT 367.950 152.400 379.050 153.600 ;
        RECT 367.950 151.950 370.050 152.400 ;
        RECT 376.950 151.950 379.050 152.400 ;
        RECT 289.950 150.600 292.050 151.050 ;
        RECT 436.950 150.600 439.050 151.050 ;
        RECT 289.950 149.400 439.050 150.600 ;
        RECT 289.950 148.950 292.050 149.400 ;
        RECT 436.950 148.950 439.050 149.400 ;
        RECT 184.950 132.600 187.050 133.050 ;
        RECT 301.950 132.600 304.050 133.050 ;
        RECT 184.950 131.400 304.050 132.600 ;
        RECT 184.950 130.950 187.050 131.400 ;
        RECT 301.950 130.950 304.050 131.400 ;
        RECT 337.950 132.600 340.050 133.050 ;
        RECT 379.950 132.600 382.050 133.050 ;
        RECT 337.950 131.400 382.050 132.600 ;
        RECT 337.950 130.950 340.050 131.400 ;
        RECT 379.950 130.950 382.050 131.400 ;
        RECT 4.950 129.600 7.050 130.050 ;
        RECT 10.950 129.600 13.050 130.050 ;
        RECT 34.950 129.600 37.050 130.050 ;
        RECT 4.950 128.400 37.050 129.600 ;
        RECT 4.950 127.950 7.050 128.400 ;
        RECT 10.950 127.950 13.050 128.400 ;
        RECT 34.950 127.950 37.050 128.400 ;
        RECT 151.950 129.600 154.050 130.050 ;
        RECT 166.950 129.600 169.050 130.050 ;
        RECT 178.950 129.600 181.050 130.050 ;
        RECT 214.950 129.600 217.050 130.050 ;
        RECT 151.950 128.400 217.050 129.600 ;
        RECT 151.950 127.950 154.050 128.400 ;
        RECT 166.950 127.950 169.050 128.400 ;
        RECT 178.950 127.950 181.050 128.400 ;
        RECT 214.950 127.950 217.050 128.400 ;
        RECT 289.950 129.600 292.050 130.050 ;
        RECT 295.950 129.600 298.050 130.050 ;
        RECT 289.950 128.400 298.050 129.600 ;
        RECT 289.950 127.950 292.050 128.400 ;
        RECT 295.950 127.950 298.050 128.400 ;
        RECT 328.950 129.600 331.050 130.050 ;
        RECT 343.950 129.600 346.050 130.050 ;
        RECT 424.950 129.600 427.050 130.050 ;
        RECT 328.950 128.400 427.050 129.600 ;
        RECT 328.950 127.950 331.050 128.400 ;
        RECT 343.950 127.950 346.050 128.400 ;
        RECT 424.950 127.950 427.050 128.400 ;
        RECT 430.950 129.600 433.050 130.050 ;
        RECT 472.950 129.600 475.050 130.050 ;
        RECT 430.950 128.400 475.050 129.600 ;
        RECT 430.950 127.950 433.050 128.400 ;
        RECT 472.950 127.950 475.050 128.400 ;
        RECT 637.950 129.600 640.050 130.050 ;
        RECT 679.950 129.600 682.050 130.050 ;
        RECT 637.950 128.400 682.050 129.600 ;
        RECT 637.950 127.950 640.050 128.400 ;
        RECT 679.950 127.950 682.050 128.400 ;
        RECT 724.950 129.600 727.050 130.050 ;
        RECT 745.950 129.600 748.050 130.050 ;
        RECT 724.950 128.400 748.050 129.600 ;
        RECT 724.950 127.950 727.050 128.400 ;
        RECT 745.950 127.950 748.050 128.400 ;
        RECT 19.950 126.600 22.050 127.050 ;
        RECT 70.950 126.600 73.050 127.050 ;
        RECT 112.950 126.600 115.050 127.050 ;
        RECT 148.950 126.600 151.050 127.050 ;
        RECT 19.950 125.400 151.050 126.600 ;
        RECT 19.950 124.950 22.050 125.400 ;
        RECT 70.950 124.950 73.050 125.400 ;
        RECT 112.950 124.950 115.050 125.400 ;
        RECT 148.950 124.950 151.050 125.400 ;
        RECT 172.950 126.600 175.050 127.050 ;
        RECT 211.950 126.600 214.050 127.050 ;
        RECT 172.950 125.400 214.050 126.600 ;
        RECT 172.950 124.950 175.050 125.400 ;
        RECT 211.950 124.950 214.050 125.400 ;
        RECT 274.950 126.600 277.050 127.050 ;
        RECT 340.950 126.600 343.050 127.050 ;
        RECT 274.950 125.400 343.050 126.600 ;
        RECT 274.950 124.950 277.050 125.400 ;
        RECT 340.950 124.950 343.050 125.400 ;
        RECT 358.950 126.600 361.050 127.050 ;
        RECT 469.950 126.600 472.050 127.050 ;
        RECT 358.950 125.400 472.050 126.600 ;
        RECT 358.950 124.950 361.050 125.400 ;
        RECT 469.950 124.950 472.050 125.400 ;
        RECT 553.950 126.600 556.050 127.050 ;
        RECT 559.950 126.600 562.050 127.050 ;
        RECT 553.950 125.400 562.050 126.600 ;
        RECT 553.950 124.950 556.050 125.400 ;
        RECT 559.950 124.950 562.050 125.400 ;
        RECT 592.950 126.600 595.050 127.050 ;
        RECT 670.950 126.600 673.050 127.050 ;
        RECT 592.950 125.400 673.050 126.600 ;
        RECT 592.950 124.950 595.050 125.400 ;
        RECT 670.950 124.950 673.050 125.400 ;
        RECT 688.950 126.600 691.050 127.050 ;
        RECT 721.950 126.600 724.050 127.050 ;
        RECT 688.950 125.400 724.050 126.600 ;
        RECT 688.950 124.950 691.050 125.400 ;
        RECT 721.950 124.950 724.050 125.400 ;
        RECT 22.950 123.600 25.050 124.050 ;
        RECT 40.950 123.600 43.050 124.050 ;
        RECT 46.950 123.600 49.050 124.050 ;
        RECT 22.950 122.400 49.050 123.600 ;
        RECT 22.950 121.950 25.050 122.400 ;
        RECT 40.950 121.950 43.050 122.400 ;
        RECT 46.950 121.950 49.050 122.400 ;
        RECT 85.950 123.600 88.050 124.050 ;
        RECT 127.950 123.600 130.050 124.050 ;
        RECT 235.950 123.600 238.050 124.050 ;
        RECT 85.950 122.400 238.050 123.600 ;
        RECT 85.950 121.950 88.050 122.400 ;
        RECT 127.950 121.950 130.050 122.400 ;
        RECT 235.950 121.950 238.050 122.400 ;
        RECT 241.950 123.600 244.050 124.050 ;
        RECT 250.950 123.600 253.050 124.050 ;
        RECT 241.950 122.400 253.050 123.600 ;
        RECT 241.950 121.950 244.050 122.400 ;
        RECT 250.950 121.950 253.050 122.400 ;
        RECT 304.950 123.600 307.050 124.050 ;
        RECT 388.950 123.600 391.050 124.050 ;
        RECT 427.950 123.600 430.050 124.050 ;
        RECT 304.950 122.400 430.050 123.600 ;
        RECT 304.950 121.950 307.050 122.400 ;
        RECT 388.950 121.950 391.050 122.400 ;
        RECT 427.950 121.950 430.050 122.400 ;
        RECT 586.950 123.600 589.050 124.050 ;
        RECT 631.950 123.600 634.050 124.050 ;
        RECT 586.950 122.400 634.050 123.600 ;
        RECT 586.950 121.950 589.050 122.400 ;
        RECT 631.950 121.950 634.050 122.400 ;
        RECT 643.950 123.600 646.050 124.050 ;
        RECT 676.950 123.600 679.050 124.050 ;
        RECT 643.950 122.400 679.050 123.600 ;
        RECT 643.950 121.950 646.050 122.400 ;
        RECT 676.950 121.950 679.050 122.400 ;
        RECT 109.950 120.600 112.050 121.050 ;
        RECT 121.950 120.600 124.050 121.050 ;
        RECT 109.950 119.400 124.050 120.600 ;
        RECT 109.950 118.950 112.050 119.400 ;
        RECT 121.950 118.950 124.050 119.400 ;
        RECT 253.950 120.600 256.050 121.050 ;
        RECT 292.950 120.600 295.050 121.050 ;
        RECT 253.950 119.400 295.050 120.600 ;
        RECT 253.950 118.950 256.050 119.400 ;
        RECT 292.950 118.950 295.050 119.400 ;
        RECT 514.950 120.600 517.050 121.050 ;
        RECT 598.950 120.600 601.050 121.050 ;
        RECT 628.950 120.600 631.050 121.050 ;
        RECT 514.950 119.400 631.050 120.600 ;
        RECT 514.950 118.950 517.050 119.400 ;
        RECT 598.950 118.950 601.050 119.400 ;
        RECT 628.950 118.950 631.050 119.400 ;
        RECT 226.950 117.600 229.050 118.050 ;
        RECT 256.950 117.600 259.050 118.050 ;
        RECT 226.950 116.400 259.050 117.600 ;
        RECT 226.950 115.950 229.050 116.400 ;
        RECT 256.950 115.950 259.050 116.400 ;
        RECT 487.950 117.600 490.050 118.050 ;
        RECT 550.950 117.600 553.050 118.050 ;
        RECT 556.950 117.600 559.050 118.050 ;
        RECT 487.950 116.400 559.050 117.600 ;
        RECT 487.950 115.950 490.050 116.400 ;
        RECT 550.950 115.950 553.050 116.400 ;
        RECT 556.950 115.950 559.050 116.400 ;
        RECT 271.950 114.600 274.050 115.050 ;
        RECT 298.950 114.600 301.050 115.050 ;
        RECT 271.950 113.400 301.050 114.600 ;
        RECT 271.950 112.950 274.050 113.400 ;
        RECT 298.950 112.950 301.050 113.400 ;
        RECT 106.950 111.600 109.050 112.050 ;
        RECT 115.950 111.600 118.050 112.050 ;
        RECT 163.950 111.600 166.050 112.050 ;
        RECT 484.950 111.600 487.050 112.050 ;
        RECT 106.950 110.400 487.050 111.600 ;
        RECT 106.950 109.950 109.050 110.400 ;
        RECT 115.950 109.950 118.050 110.400 ;
        RECT 163.950 109.950 166.050 110.400 ;
        RECT 484.950 109.950 487.050 110.400 ;
        RECT 142.950 102.600 145.050 103.050 ;
        RECT 169.950 102.600 172.050 103.050 ;
        RECT 142.950 101.400 172.050 102.600 ;
        RECT 142.950 100.950 145.050 101.400 ;
        RECT 169.950 100.950 172.050 101.400 ;
        RECT 187.950 102.600 190.050 103.050 ;
        RECT 190.950 102.600 193.050 103.050 ;
        RECT 238.950 102.600 241.050 103.050 ;
        RECT 187.950 101.400 241.050 102.600 ;
        RECT 187.950 100.950 190.050 101.400 ;
        RECT 190.950 100.950 193.050 101.400 ;
        RECT 238.950 100.950 241.050 101.400 ;
        RECT 460.950 102.600 463.050 103.050 ;
        RECT 502.950 102.600 505.050 103.050 ;
        RECT 661.950 102.600 664.050 103.050 ;
        RECT 460.950 101.400 664.050 102.600 ;
        RECT 460.950 100.950 463.050 101.400 ;
        RECT 502.950 100.950 505.050 101.400 ;
        RECT 661.950 100.950 664.050 101.400 ;
        RECT 37.950 99.600 40.050 100.050 ;
        RECT 67.950 99.600 70.050 100.050 ;
        RECT 37.950 98.400 70.050 99.600 ;
        RECT 37.950 97.950 40.050 98.400 ;
        RECT 67.950 97.950 70.050 98.400 ;
        RECT 148.950 99.600 151.050 100.050 ;
        RECT 175.950 99.600 178.050 100.050 ;
        RECT 181.950 99.600 184.050 100.050 ;
        RECT 148.950 98.400 184.050 99.600 ;
        RECT 148.950 97.950 151.050 98.400 ;
        RECT 175.950 97.950 178.050 98.400 ;
        RECT 181.950 97.950 184.050 98.400 ;
        RECT 232.950 99.600 235.050 100.050 ;
        RECT 277.950 99.600 280.050 100.050 ;
        RECT 322.950 99.600 325.050 100.050 ;
        RECT 232.950 98.400 325.050 99.600 ;
        RECT 232.950 97.950 235.050 98.400 ;
        RECT 277.950 97.950 280.050 98.400 ;
        RECT 322.950 97.950 325.050 98.400 ;
        RECT 436.950 99.600 439.050 100.050 ;
        RECT 442.950 99.600 445.050 100.050 ;
        RECT 505.950 99.600 508.050 100.050 ;
        RECT 559.950 99.600 562.050 100.050 ;
        RECT 436.950 98.400 508.050 99.600 ;
        RECT 436.950 97.950 439.050 98.400 ;
        RECT 442.950 97.950 445.050 98.400 ;
        RECT 505.950 97.950 508.050 98.400 ;
        RECT 557.400 98.400 562.050 99.600 ;
        RECT 160.950 96.600 163.050 97.050 ;
        RECT 226.950 96.600 229.050 97.050 ;
        RECT 160.950 95.400 229.050 96.600 ;
        RECT 160.950 94.950 163.050 95.400 ;
        RECT 226.950 94.950 229.050 95.400 ;
        RECT 340.950 96.600 343.050 97.050 ;
        RECT 400.950 96.600 403.050 97.050 ;
        RECT 340.950 95.400 403.050 96.600 ;
        RECT 340.950 94.950 343.050 95.400 ;
        RECT 400.950 94.950 403.050 95.400 ;
        RECT 541.950 96.600 544.050 97.050 ;
        RECT 553.950 96.600 556.050 97.050 ;
        RECT 541.950 95.400 556.050 96.600 ;
        RECT 541.950 94.950 544.050 95.400 ;
        RECT 553.950 94.950 556.050 95.400 ;
        RECT 557.400 94.050 558.600 98.400 ;
        RECT 559.950 97.950 562.050 98.400 ;
        RECT 700.950 99.600 703.050 100.050 ;
        RECT 709.950 99.600 712.050 100.050 ;
        RECT 700.950 98.400 712.050 99.600 ;
        RECT 700.950 97.950 703.050 98.400 ;
        RECT 709.950 97.950 712.050 98.400 ;
        RECT 559.950 96.600 562.050 97.050 ;
        RECT 565.950 96.600 568.050 97.050 ;
        RECT 559.950 95.400 568.050 96.600 ;
        RECT 559.950 94.950 562.050 95.400 ;
        RECT 565.950 94.950 568.050 95.400 ;
        RECT 79.950 93.600 82.050 94.050 ;
        RECT 124.950 93.600 127.050 94.050 ;
        RECT 79.950 92.400 127.050 93.600 ;
        RECT 79.950 91.950 82.050 92.400 ;
        RECT 124.950 91.950 127.050 92.400 ;
        RECT 169.950 93.600 172.050 94.050 ;
        RECT 184.950 93.600 187.050 94.050 ;
        RECT 169.950 92.400 187.050 93.600 ;
        RECT 169.950 91.950 172.050 92.400 ;
        RECT 184.950 91.950 187.050 92.400 ;
        RECT 382.950 93.600 385.050 94.050 ;
        RECT 403.950 93.600 406.050 94.050 ;
        RECT 382.950 92.400 406.050 93.600 ;
        RECT 382.950 91.950 385.050 92.400 ;
        RECT 403.950 91.950 406.050 92.400 ;
        RECT 556.950 91.950 559.050 94.050 ;
        RECT 562.950 93.600 565.050 94.050 ;
        RECT 604.950 93.600 607.050 94.050 ;
        RECT 562.950 92.400 607.050 93.600 ;
        RECT 562.950 91.950 565.050 92.400 ;
        RECT 604.950 91.950 607.050 92.400 ;
        RECT 70.950 90.600 73.050 91.050 ;
        RECT 73.950 90.600 76.050 91.050 ;
        RECT 76.950 90.600 79.050 91.050 ;
        RECT 118.950 90.600 121.050 91.050 ;
        RECT 70.950 89.400 121.050 90.600 ;
        RECT 70.950 88.950 73.050 89.400 ;
        RECT 73.950 88.950 76.050 89.400 ;
        RECT 76.950 88.950 79.050 89.400 ;
        RECT 118.950 88.950 121.050 89.400 ;
        RECT 283.950 90.600 286.050 91.050 ;
        RECT 313.950 90.600 316.050 91.050 ;
        RECT 283.950 89.400 316.050 90.600 ;
        RECT 283.950 88.950 286.050 89.400 ;
        RECT 313.950 88.950 316.050 89.400 ;
        RECT 361.950 90.600 364.050 91.050 ;
        RECT 382.950 90.600 385.050 91.050 ;
        RECT 361.950 89.400 385.050 90.600 ;
        RECT 361.950 88.950 364.050 89.400 ;
        RECT 382.950 88.950 385.050 89.400 ;
        RECT 511.950 90.600 514.050 91.050 ;
        RECT 565.950 90.600 568.050 91.050 ;
        RECT 511.950 89.400 568.050 90.600 ;
        RECT 511.950 88.950 514.050 89.400 ;
        RECT 565.950 88.950 568.050 89.400 ;
        RECT 613.950 90.600 616.050 91.050 ;
        RECT 703.950 90.600 706.050 91.050 ;
        RECT 742.950 90.600 745.050 91.050 ;
        RECT 613.950 89.400 745.050 90.600 ;
        RECT 613.950 88.950 616.050 89.400 ;
        RECT 703.950 88.950 706.050 89.400 ;
        RECT 742.950 88.950 745.050 89.400 ;
        RECT 394.950 84.600 397.050 85.050 ;
        RECT 400.950 84.600 403.050 85.050 ;
        RECT 394.950 83.400 403.050 84.600 ;
        RECT 394.950 82.950 397.050 83.400 ;
        RECT 400.950 82.950 403.050 83.400 ;
        RECT 514.950 78.600 517.050 79.050 ;
        RECT 586.950 78.600 589.050 79.050 ;
        RECT 514.950 77.400 589.050 78.600 ;
        RECT 514.950 76.950 517.050 77.400 ;
        RECT 586.950 76.950 589.050 77.400 ;
        RECT 427.950 63.600 430.050 64.050 ;
        RECT 445.950 63.600 448.050 64.050 ;
        RECT 427.950 62.400 448.050 63.600 ;
        RECT 427.950 61.950 430.050 62.400 ;
        RECT 445.950 61.950 448.050 62.400 ;
        RECT 634.950 60.600 637.050 61.050 ;
        RECT 709.950 60.600 712.050 61.050 ;
        RECT 634.950 59.400 712.050 60.600 ;
        RECT 634.950 58.950 637.050 59.400 ;
        RECT 709.950 58.950 712.050 59.400 ;
        RECT 196.950 57.600 199.050 58.050 ;
        RECT 211.950 57.600 214.050 58.050 ;
        RECT 196.950 56.400 214.050 57.600 ;
        RECT 196.950 55.950 199.050 56.400 ;
        RECT 211.950 55.950 214.050 56.400 ;
        RECT 373.950 57.600 376.050 58.050 ;
        RECT 439.950 57.600 442.050 58.050 ;
        RECT 547.950 57.600 550.050 58.050 ;
        RECT 550.950 57.600 553.050 58.050 ;
        RECT 598.950 57.600 601.050 58.050 ;
        RECT 373.950 56.400 601.050 57.600 ;
        RECT 373.950 55.950 376.050 56.400 ;
        RECT 439.950 55.950 442.050 56.400 ;
        RECT 547.950 55.950 550.050 56.400 ;
        RECT 550.950 55.950 553.050 56.400 ;
        RECT 598.950 55.950 601.050 56.400 ;
        RECT 676.950 57.600 679.050 58.050 ;
        RECT 715.950 57.600 718.050 58.050 ;
        RECT 754.950 57.600 757.050 58.050 ;
        RECT 676.950 56.400 757.050 57.600 ;
        RECT 676.950 55.950 679.050 56.400 ;
        RECT 715.950 55.950 718.050 56.400 ;
        RECT 754.950 55.950 757.050 56.400 ;
        RECT 67.950 54.600 70.050 55.050 ;
        RECT 73.950 54.600 76.050 55.050 ;
        RECT 67.950 53.400 76.050 54.600 ;
        RECT 67.950 52.950 70.050 53.400 ;
        RECT 73.950 52.950 76.050 53.400 ;
        RECT 178.950 54.600 181.050 55.050 ;
        RECT 199.950 54.600 202.050 55.050 ;
        RECT 178.950 53.400 202.050 54.600 ;
        RECT 178.950 52.950 181.050 53.400 ;
        RECT 199.950 52.950 202.050 53.400 ;
        RECT 307.950 54.600 310.050 55.050 ;
        RECT 322.950 54.600 325.050 55.050 ;
        RECT 355.950 54.600 358.050 55.050 ;
        RECT 307.950 53.400 358.050 54.600 ;
        RECT 307.950 52.950 310.050 53.400 ;
        RECT 322.950 52.950 325.050 53.400 ;
        RECT 355.950 52.950 358.050 53.400 ;
        RECT 370.950 54.600 373.050 55.050 ;
        RECT 436.950 54.600 439.050 55.050 ;
        RECT 370.950 53.400 439.050 54.600 ;
        RECT 370.950 52.950 373.050 53.400 ;
        RECT 436.950 52.950 439.050 53.400 ;
        RECT 553.950 54.600 556.050 55.050 ;
        RECT 592.950 54.600 595.050 55.050 ;
        RECT 553.950 53.400 595.050 54.600 ;
        RECT 553.950 52.950 556.050 53.400 ;
        RECT 592.950 52.950 595.050 53.400 ;
        RECT 712.950 54.600 715.050 55.050 ;
        RECT 718.950 54.600 721.050 55.050 ;
        RECT 712.950 53.400 721.050 54.600 ;
        RECT 712.950 52.950 715.050 53.400 ;
        RECT 718.950 52.950 721.050 53.400 ;
        RECT 73.950 51.600 76.050 52.050 ;
        RECT 151.950 51.600 154.050 52.050 ;
        RECT 73.950 50.400 154.050 51.600 ;
        RECT 73.950 49.950 76.050 50.400 ;
        RECT 151.950 49.950 154.050 50.400 ;
        RECT 160.950 51.600 163.050 52.050 ;
        RECT 205.950 51.600 208.050 52.050 ;
        RECT 247.950 51.600 250.050 52.050 ;
        RECT 160.950 50.400 250.050 51.600 ;
        RECT 160.950 49.950 163.050 50.400 ;
        RECT 205.950 49.950 208.050 50.400 ;
        RECT 247.950 49.950 250.050 50.400 ;
        RECT 361.950 51.600 364.050 52.050 ;
        RECT 445.950 51.600 448.050 52.050 ;
        RECT 361.950 50.400 448.050 51.600 ;
        RECT 361.950 49.950 364.050 50.400 ;
        RECT 445.950 49.950 448.050 50.400 ;
        RECT 601.950 51.600 604.050 52.050 ;
        RECT 613.950 51.600 616.050 52.050 ;
        RECT 601.950 50.400 616.050 51.600 ;
        RECT 601.950 49.950 604.050 50.400 ;
        RECT 613.950 49.950 616.050 50.400 ;
        RECT 622.950 51.600 625.050 52.050 ;
        RECT 664.950 51.600 667.050 52.050 ;
        RECT 622.950 50.400 667.050 51.600 ;
        RECT 622.950 49.950 625.050 50.400 ;
        RECT 664.950 49.950 667.050 50.400 ;
        RECT 115.950 48.600 118.050 49.050 ;
        RECT 154.950 48.600 157.050 49.050 ;
        RECT 115.950 47.400 157.050 48.600 ;
        RECT 115.950 46.950 118.050 47.400 ;
        RECT 154.950 46.950 157.050 47.400 ;
        RECT 241.950 48.600 244.050 49.050 ;
        RECT 286.950 48.600 289.050 49.050 ;
        RECT 241.950 47.400 289.050 48.600 ;
        RECT 241.950 46.950 244.050 47.400 ;
        RECT 286.950 46.950 289.050 47.400 ;
        RECT 313.950 48.600 316.050 49.050 ;
        RECT 364.950 48.600 367.050 49.050 ;
        RECT 313.950 47.400 367.050 48.600 ;
        RECT 446.400 48.600 447.600 49.950 ;
        RECT 508.950 48.600 511.050 49.050 ;
        RECT 446.400 47.400 511.050 48.600 ;
        RECT 313.950 46.950 316.050 47.400 ;
        RECT 364.950 46.950 367.050 47.400 ;
        RECT 508.950 46.950 511.050 47.400 ;
        RECT 595.950 48.600 598.050 49.050 ;
        RECT 616.950 48.600 619.050 49.050 ;
        RECT 595.950 47.400 619.050 48.600 ;
        RECT 595.950 46.950 598.050 47.400 ;
        RECT 616.950 46.950 619.050 47.400 ;
        RECT 76.950 45.600 79.050 46.050 ;
        RECT 118.950 45.600 121.050 46.050 ;
        RECT 166.950 45.600 169.050 46.050 ;
        RECT 76.950 44.400 169.050 45.600 ;
        RECT 76.950 43.950 79.050 44.400 ;
        RECT 118.950 43.950 121.050 44.400 ;
        RECT 166.950 43.950 169.050 44.400 ;
        RECT 328.950 45.600 331.050 46.050 ;
        RECT 424.950 45.600 427.050 46.050 ;
        RECT 457.950 45.600 460.050 46.050 ;
        RECT 328.950 44.400 460.050 45.600 ;
        RECT 328.950 43.950 331.050 44.400 ;
        RECT 424.950 43.950 427.050 44.400 ;
        RECT 457.950 43.950 460.050 44.400 ;
        RECT 463.950 45.600 466.050 46.050 ;
        RECT 508.950 45.600 511.050 46.050 ;
        RECT 463.950 44.400 511.050 45.600 ;
        RECT 463.950 43.950 466.050 44.400 ;
        RECT 508.950 43.950 511.050 44.400 ;
        RECT 376.950 39.600 379.050 40.050 ;
        RECT 403.950 39.600 406.050 40.050 ;
        RECT 715.950 39.600 718.050 40.050 ;
        RECT 376.950 38.400 718.050 39.600 ;
        RECT 376.950 37.950 379.050 38.400 ;
        RECT 403.950 37.950 406.050 38.400 ;
        RECT 715.950 37.950 718.050 38.400 ;
        RECT 106.950 30.600 109.050 31.050 ;
        RECT 259.950 30.600 262.050 31.050 ;
        RECT 376.950 30.600 379.050 31.050 ;
        RECT 106.950 29.400 379.050 30.600 ;
        RECT 106.950 28.950 109.050 29.400 ;
        RECT 259.950 28.950 262.050 29.400 ;
        RECT 376.950 28.950 379.050 29.400 ;
        RECT 34.950 27.600 37.050 28.050 ;
        RECT 49.950 27.600 52.050 28.050 ;
        RECT 112.950 27.600 115.050 28.050 ;
        RECT 34.950 26.400 115.050 27.600 ;
        RECT 34.950 25.950 37.050 26.400 ;
        RECT 49.950 25.950 52.050 26.400 ;
        RECT 112.950 25.950 115.050 26.400 ;
        RECT 19.950 24.600 22.050 25.050 ;
        RECT 55.950 24.600 58.050 25.050 ;
        RECT 19.950 23.400 58.050 24.600 ;
        RECT 19.950 22.950 22.050 23.400 ;
        RECT 55.950 22.950 58.050 23.400 ;
        RECT 67.950 24.600 70.050 25.050 ;
        RECT 76.950 24.600 79.050 25.050 ;
        RECT 67.950 23.400 79.050 24.600 ;
        RECT 67.950 22.950 70.050 23.400 ;
        RECT 76.950 22.950 79.050 23.400 ;
        RECT 79.950 24.600 82.050 25.050 ;
        RECT 103.950 24.600 106.050 25.050 ;
        RECT 79.950 23.400 106.050 24.600 ;
        RECT 79.950 22.950 82.050 23.400 ;
        RECT 103.950 22.950 106.050 23.400 ;
        RECT 175.950 24.600 178.050 25.050 ;
        RECT 205.950 24.600 208.050 25.050 ;
        RECT 211.950 24.600 214.050 25.050 ;
        RECT 280.950 24.600 283.050 25.050 ;
        RECT 175.950 23.400 208.050 24.600 ;
        RECT 175.950 22.950 178.050 23.400 ;
        RECT 205.950 22.950 208.050 23.400 ;
        RECT 209.400 23.400 283.050 24.600 ;
        RECT 31.950 21.600 34.050 22.050 ;
        RECT 79.950 21.600 82.050 22.050 ;
        RECT 31.950 20.400 82.050 21.600 ;
        RECT 31.950 19.950 34.050 20.400 ;
        RECT 79.950 19.950 82.050 20.400 ;
        RECT 112.950 21.600 115.050 22.050 ;
        RECT 148.950 21.600 151.050 22.050 ;
        RECT 112.950 20.400 151.050 21.600 ;
        RECT 112.950 19.950 115.050 20.400 ;
        RECT 148.950 19.950 151.050 20.400 ;
        RECT 184.950 21.600 187.050 22.050 ;
        RECT 209.400 21.600 210.600 23.400 ;
        RECT 211.950 22.950 214.050 23.400 ;
        RECT 280.950 22.950 283.050 23.400 ;
        RECT 301.950 24.600 304.050 25.050 ;
        RECT 322.950 24.600 325.050 25.050 ;
        RECT 301.950 23.400 325.050 24.600 ;
        RECT 301.950 22.950 304.050 23.400 ;
        RECT 322.950 22.950 325.050 23.400 ;
        RECT 325.950 24.600 328.050 25.050 ;
        RECT 340.950 24.600 343.050 25.050 ;
        RECT 325.950 23.400 343.050 24.600 ;
        RECT 325.950 22.950 328.050 23.400 ;
        RECT 340.950 22.950 343.050 23.400 ;
        RECT 595.950 24.600 598.050 25.050 ;
        RECT 616.950 24.600 619.050 25.050 ;
        RECT 595.950 23.400 619.050 24.600 ;
        RECT 595.950 22.950 598.050 23.400 ;
        RECT 616.950 22.950 619.050 23.400 ;
        RECT 634.950 24.600 637.050 25.050 ;
        RECT 667.950 24.600 670.050 25.050 ;
        RECT 634.950 23.400 670.050 24.600 ;
        RECT 634.950 22.950 637.050 23.400 ;
        RECT 667.950 22.950 670.050 23.400 ;
        RECT 184.950 20.400 210.600 21.600 ;
        RECT 262.950 21.600 265.050 22.050 ;
        RECT 298.950 21.600 301.050 22.050 ;
        RECT 262.950 20.400 301.050 21.600 ;
        RECT 184.950 19.950 187.050 20.400 ;
        RECT 262.950 19.950 265.050 20.400 ;
        RECT 298.950 19.950 301.050 20.400 ;
        RECT 382.950 21.600 385.050 22.050 ;
        RECT 418.950 21.600 421.050 22.050 ;
        RECT 382.950 20.400 421.050 21.600 ;
        RECT 382.950 19.950 385.050 20.400 ;
        RECT 418.950 19.950 421.050 20.400 ;
        RECT 466.950 21.600 469.050 22.050 ;
        RECT 505.950 21.600 508.050 22.050 ;
        RECT 466.950 20.400 508.050 21.600 ;
        RECT 466.950 19.950 469.050 20.400 ;
        RECT 505.950 19.950 508.050 20.400 ;
        RECT 553.950 21.600 556.050 22.050 ;
        RECT 592.950 21.600 595.050 22.050 ;
        RECT 553.950 20.400 595.050 21.600 ;
        RECT 553.950 19.950 556.050 20.400 ;
        RECT 592.950 19.950 595.050 20.400 ;
        RECT 604.950 21.600 607.050 22.050 ;
        RECT 673.950 21.600 676.050 22.050 ;
        RECT 721.950 21.600 724.050 22.050 ;
        RECT 751.950 21.600 754.050 22.050 ;
        RECT 604.950 20.400 720.600 21.600 ;
        RECT 604.950 19.950 607.050 20.400 ;
        RECT 673.950 19.950 676.050 20.400 ;
        RECT 259.950 18.600 262.050 19.050 ;
        RECT 283.950 18.600 286.050 19.050 ;
        RECT 304.950 18.600 307.050 19.050 ;
        RECT 373.950 18.600 376.050 19.050 ;
        RECT 259.950 17.400 376.050 18.600 ;
        RECT 259.950 16.950 262.050 17.400 ;
        RECT 283.950 16.950 286.050 17.400 ;
        RECT 304.950 16.950 307.050 17.400 ;
        RECT 373.950 16.950 376.050 17.400 ;
        RECT 379.950 18.600 382.050 19.050 ;
        RECT 424.950 18.600 427.050 19.050 ;
        RECT 463.950 18.600 466.050 19.050 ;
        RECT 511.950 18.600 514.050 19.050 ;
        RECT 379.950 17.400 514.050 18.600 ;
        RECT 379.950 16.950 382.050 17.400 ;
        RECT 424.950 16.950 427.050 17.400 ;
        RECT 463.950 16.950 466.050 17.400 ;
        RECT 511.950 16.950 514.050 17.400 ;
        RECT 550.950 18.600 553.050 19.050 ;
        RECT 598.950 18.600 601.050 19.050 ;
        RECT 550.950 17.400 601.050 18.600 ;
        RECT 550.950 16.950 553.050 17.400 ;
        RECT 598.950 16.950 601.050 17.400 ;
        RECT 676.950 18.600 679.050 19.050 ;
        RECT 712.950 18.600 715.050 19.050 ;
        RECT 676.950 17.400 715.050 18.600 ;
        RECT 719.400 18.600 720.600 20.400 ;
        RECT 721.950 20.400 754.050 21.600 ;
        RECT 721.950 19.950 724.050 20.400 ;
        RECT 751.950 19.950 754.050 20.400 ;
        RECT 754.950 18.600 757.050 19.050 ;
        RECT 719.400 17.400 757.050 18.600 ;
        RECT 676.950 16.950 679.050 17.400 ;
        RECT 712.950 16.950 715.050 17.400 ;
        RECT 754.950 16.950 757.050 17.400 ;
  END
END output_terminal
END LIBRARY

