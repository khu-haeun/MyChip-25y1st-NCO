magic
tech scmos
magscale 1 2
timestamp 1764070200
<< metal1 >>
rect -62 16818 -2 17058
rect 17170 17042 17262 17058
rect -62 16802 30 16818
rect -62 16338 -2 16802
rect 17202 16578 17262 17042
rect 17170 16562 17262 16578
rect -62 16322 30 16338
rect -62 15858 -2 16322
rect 17202 16098 17262 16562
rect 17170 16082 17262 16098
rect -62 15842 30 15858
rect -62 15378 -2 15842
rect 17202 15618 17262 16082
rect 17170 15602 17262 15618
rect -62 15362 30 15378
rect -62 14898 -2 15362
rect 17202 15138 17262 15602
rect 17170 15122 17262 15138
rect -62 14882 30 14898
rect -62 14418 -2 14882
rect 17202 14658 17262 15122
rect 17170 14642 17262 14658
rect -62 14402 30 14418
rect -62 13938 -2 14402
rect 17202 14178 17262 14642
rect 17170 14162 17262 14178
rect -62 13922 30 13938
rect -62 13458 -2 13922
rect 17202 13698 17262 14162
rect 17170 13682 17262 13698
rect -62 13442 30 13458
rect -62 12978 -2 13442
rect 17202 13218 17262 13682
rect 17170 13202 17262 13218
rect -62 12962 30 12978
rect -62 12498 -2 12962
rect 17202 12738 17262 13202
rect 17170 12722 17262 12738
rect -62 12482 30 12498
rect -62 12018 -2 12482
rect 17202 12258 17262 12722
rect 17170 12242 17262 12258
rect -62 12002 30 12018
rect -62 11538 -2 12002
rect 17202 11778 17262 12242
rect 17170 11762 17262 11778
rect -62 11522 30 11538
rect -62 11058 -2 11522
rect 17202 11298 17262 11762
rect 17170 11282 17262 11298
rect -62 11042 30 11058
rect -62 10578 -2 11042
rect 17202 10818 17262 11282
rect 17170 10802 17262 10818
rect -62 10562 30 10578
rect -62 10098 -2 10562
rect 17202 10338 17262 10802
rect 17170 10322 17262 10338
rect -62 10082 30 10098
rect -62 9618 -2 10082
rect 17202 9858 17262 10322
rect 17170 9842 17262 9858
rect -62 9602 30 9618
rect -62 9138 -2 9602
rect 17202 9378 17262 9842
rect 17170 9362 17262 9378
rect -62 9122 30 9138
rect -62 8658 -2 9122
rect 17202 8898 17262 9362
rect 17170 8882 17262 8898
rect -62 8642 30 8658
rect -62 8178 -2 8642
rect 17202 8418 17262 8882
rect 17170 8402 17262 8418
rect -62 8162 30 8178
rect -62 7698 -2 8162
rect 17202 7938 17262 8402
rect 17170 7922 17262 7938
rect -62 7682 30 7698
rect -62 7218 -2 7682
rect 17202 7458 17262 7922
rect 17170 7442 17262 7458
rect -62 7202 30 7218
rect -62 6738 -2 7202
rect 17202 6978 17262 7442
rect 17170 6962 17262 6978
rect -62 6722 30 6738
rect -62 6258 -2 6722
rect 17202 6498 17262 6962
rect 17170 6482 17262 6498
rect -62 6242 30 6258
rect -62 5778 -2 6242
rect 17202 6018 17262 6482
rect 17170 6002 17262 6018
rect -62 5762 30 5778
rect -62 5298 -2 5762
rect 17202 5538 17262 6002
rect 17170 5522 17262 5538
rect -62 5282 30 5298
rect -62 4818 -2 5282
rect 17202 5058 17262 5522
rect 17170 5042 17262 5058
rect -62 4802 30 4818
rect -62 4338 -2 4802
rect 17202 4578 17262 5042
rect 17170 4562 17262 4578
rect -62 4322 30 4338
rect -62 3858 -2 4322
rect 17202 4098 17262 4562
rect 17170 4082 17262 4098
rect -62 3842 30 3858
rect -62 3378 -2 3842
rect 17202 3618 17262 4082
rect 17170 3602 17262 3618
rect -62 3362 30 3378
rect -62 2898 -2 3362
rect 17202 3138 17262 3602
rect 17170 3122 17262 3138
rect -62 2882 30 2898
rect -62 2418 -2 2882
rect 17202 2658 17262 3122
rect 17170 2642 17262 2658
rect -62 2402 30 2418
rect -62 1938 -2 2402
rect 17202 2178 17262 2642
rect 17170 2162 17262 2178
rect -62 1922 30 1938
rect -62 1458 -2 1922
rect 17202 1698 17262 2162
rect 17170 1682 17262 1698
rect -62 1442 30 1458
rect -62 978 -2 1442
rect 17202 1218 17262 1682
rect 17170 1202 17262 1218
rect -62 962 30 978
rect -62 498 -2 962
rect 17202 738 17262 1202
rect 17170 722 17262 738
rect -62 482 30 498
rect -62 18 -2 482
rect 17202 258 17262 722
rect 17170 242 17262 258
rect -62 2 30 18
rect 17202 2 17262 242
<< metal2 >>
rect 8317 17097 8323 17103
rect 8957 17097 8963 17103
rect 7637 -23 7643 -17
rect 7997 -23 8003 -17
rect 8117 -23 8123 -17
rect 8157 -23 8163 -17
rect 8297 -23 8303 -17
rect 8497 -23 8503 -17
rect 8537 -23 8543 -17
rect 9037 -23 9043 -17
rect 9177 -23 9183 -17
rect 9817 -23 9823 -17
rect 10317 -23 10323 -17
rect 10717 -23 10723 -17
rect 11137 -23 11143 -17
rect 11317 -23 11323 -17
rect 12097 -23 12103 -17
rect 12177 -23 12183 -17
rect 12357 -23 12363 -17
rect 13657 -23 13663 -17
rect 13897 -23 13903 -17
rect 14417 -23 14423 -17
rect 14637 -23 14643 -17
rect 14677 -23 14683 -17
rect 14717 -23 14723 -17
rect 15017 -23 15023 -17
rect 15457 -23 15463 -17
rect 15677 -23 15683 -17
rect 15837 -23 15843 -17
rect 16137 -23 16143 -17
rect 16977 -23 16983 -17
<< metal3 >>
rect -24 8036 -16 8044
rect -24 7556 -16 7564
rect -24 7096 -16 7104
rect -24 7056 -16 7064
rect 17236 1796 17244 1804
rect 17236 116 17244 124
use INVX1  _7072_
timestamp 0
transform 1 0 6190 0 1 6490
box -6 -8 66 248
use INVX2  _7073_
timestamp 0
transform 1 0 8830 0 1 4570
box -6 -8 66 248
use NOR2X1  _7074_
timestamp 0
transform 1 0 6730 0 -1 4570
box -6 -8 86 248
use INVX2  _7075_
timestamp 0
transform 1 0 7670 0 1 4090
box -6 -8 66 248
use NOR2X1  _7076_
timestamp 0
transform -1 0 5930 0 -1 5050
box -6 -8 86 248
use INVX4  _7077_
timestamp 0
transform -1 0 8690 0 -1 5050
box -6 -8 86 248
use NOR2X1  _7078_
timestamp 0
transform -1 0 5550 0 1 4570
box -6 -8 86 248
use OAI21X1  _7079_
timestamp 0
transform -1 0 6910 0 -1 5050
box -6 -8 106 248
use INVX2  _7080_
timestamp 0
transform -1 0 8670 0 -1 4570
box -6 -8 66 248
use AND2X2  _7081_
timestamp 0
transform -1 0 5530 0 1 5050
box -6 -8 106 248
use AOI22X1  _7082_
timestamp 0
transform -1 0 6510 0 1 5050
box -6 -8 126 248
use OAI21X1  _7083_
timestamp 0
transform 1 0 5970 0 -1 5050
box -6 -8 106 248
use NOR2X1  _7084_
timestamp 0
transform 1 0 8710 0 1 4570
box -6 -8 86 248
use AOI22X1  _7085_
timestamp 0
transform 1 0 5850 0 1 5050
box -6 -8 126 248
use OAI21X1  _7086_
timestamp 0
transform -1 0 5730 0 -1 6010
box -6 -8 106 248
use INVX1  _7087_
timestamp 0
transform -1 0 5550 0 -1 5050
box -6 -8 66 248
use OAI21X1  _7088_
timestamp 0
transform -1 0 5310 0 -1 5050
box -6 -8 106 248
use AOI21X1  _7089_
timestamp 0
transform -1 0 5450 0 -1 5050
box -6 -8 106 248
use INVX1  _7090_
timestamp 0
transform -1 0 7930 0 1 5050
box -6 -8 66 248
use NAND2X1  _7091_
timestamp 0
transform -1 0 5530 0 -1 5530
box -6 -8 86 248
use OAI21X1  _7092_
timestamp 0
transform -1 0 5670 0 1 5050
box -6 -8 106 248
use OAI21X1  _7093_
timestamp 0
transform -1 0 5370 0 1 5050
box -6 -8 106 248
use AOI22X1  _7094_
timestamp 0
transform 1 0 5330 0 -1 6010
box -6 -8 126 248
use NAND2X1  _7095_
timestamp 0
transform -1 0 5290 0 -1 6010
box -6 -8 86 248
use INVX1  _7096_
timestamp 0
transform -1 0 5770 0 -1 3610
box -6 -8 66 248
use OAI21X1  _7097_
timestamp 0
transform -1 0 5910 0 -1 3610
box -6 -8 106 248
use AOI21X1  _7098_
timestamp 0
transform -1 0 5930 0 1 3610
box -6 -8 106 248
use INVX1  _7099_
timestamp 0
transform 1 0 5650 0 1 3130
box -6 -8 66 248
use NAND2X1  _7100_
timestamp 0
transform 1 0 5490 0 -1 4090
box -6 -8 86 248
use OAI21X1  _7101_
timestamp 0
transform 1 0 5390 0 1 4090
box -6 -8 106 248
use OAI21X1  _7102_
timestamp 0
transform -1 0 5350 0 1 4090
box -6 -8 106 248
use AOI22X1  _7103_
timestamp 0
transform 1 0 6430 0 -1 4090
box -6 -8 126 248
use NAND2X1  _7104_
timestamp 0
transform 1 0 5130 0 1 4090
box -6 -8 86 248
use INVX1  _7105_
timestamp 0
transform 1 0 5370 0 1 4570
box -6 -8 66 248
use OAI21X1  _7106_
timestamp 0
transform 1 0 4990 0 1 4090
box -6 -8 106 248
use AOI21X1  _7107_
timestamp 0
transform 1 0 4930 0 -1 4570
box -6 -8 106 248
use INVX1  _7108_
timestamp 0
transform 1 0 5970 0 -1 4090
box -6 -8 66 248
use NAND2X1  _7109_
timestamp 0
transform 1 0 5230 0 -1 4570
box -6 -8 86 248
use OAI21X1  _7110_
timestamp 0
transform -1 0 5470 0 -1 4570
box -6 -8 106 248
use OAI21X1  _7111_
timestamp 0
transform 1 0 5510 0 -1 4570
box -6 -8 106 248
use AOI22X1  _7112_
timestamp 0
transform -1 0 6370 0 -1 4090
box -6 -8 126 248
use NAND2X1  _7113_
timestamp 0
transform -1 0 5670 0 1 4570
box -6 -8 86 248
use INVX1  _7114_
timestamp 0
transform -1 0 10430 0 1 3610
box -6 -8 66 248
use OAI21X1  _7115_
timestamp 0
transform -1 0 9090 0 1 4090
box -6 -8 106 248
use AOI21X1  _7116_
timestamp 0
transform -1 0 8930 0 1 4090
box -6 -8 106 248
use INVX1  _7117_
timestamp 0
transform -1 0 10870 0 1 3130
box -6 -8 66 248
use NAND2X1  _7118_
timestamp 0
transform -1 0 9090 0 -1 4570
box -6 -8 86 248
use OAI21X1  _7119_
timestamp 0
transform 1 0 8690 0 1 4090
box -6 -8 106 248
use OAI21X1  _7120_
timestamp 0
transform -1 0 8130 0 1 4090
box -6 -8 106 248
use AOI22X1  _7121_
timestamp 0
transform -1 0 8210 0 -1 4090
box -6 -8 126 248
use NAND2X1  _7122_
timestamp 0
transform -1 0 7990 0 1 4090
box -6 -8 86 248
use INVX1  _7123_
timestamp 0
transform -1 0 9510 0 -1 3610
box -6 -8 66 248
use NOR2X1  _7124_
timestamp 0
transform 1 0 9150 0 1 4090
box -6 -8 86 248
use OAI21X1  _7125_
timestamp 0
transform -1 0 9350 0 1 3610
box -6 -8 106 248
use AOI22X1  _7126_
timestamp 0
transform 1 0 9270 0 -1 4090
box -6 -8 126 248
use OAI21X1  _7127_
timestamp 0
transform 1 0 9130 0 -1 4090
box -6 -8 106 248
use AOI22X1  _7128_
timestamp 0
transform 1 0 8790 0 -1 4090
box -6 -8 126 248
use OAI21X1  _7129_
timestamp 0
transform -1 0 9070 0 -1 4090
box -6 -8 106 248
use INVX1  _7130_
timestamp 0
transform 1 0 7470 0 -1 4090
box -6 -8 66 248
use INVX1  _7131_
timestamp 0
transform 1 0 8510 0 -1 3130
box -6 -8 66 248
use INVX8  _7132_
timestamp 0
transform 1 0 8470 0 -1 1210
box -6 -8 126 248
use INVX8  _7133_
timestamp 0
transform 1 0 7410 0 -1 250
box -6 -8 126 248
use INVX1  _7134_
timestamp 0
transform 1 0 13090 0 -1 2170
box -6 -8 66 248
use NAND2X1  _7135_
timestamp 0
transform 1 0 13290 0 1 2170
box -6 -8 86 248
use OAI21X1  _7136_
timestamp 0
transform 1 0 13150 0 1 2170
box -6 -8 106 248
use INVX1  _7137_
timestamp 0
transform 1 0 12030 0 -1 2170
box -6 -8 66 248
use NAND2X1  _7138_
timestamp 0
transform -1 0 10570 0 -1 2170
box -6 -8 86 248
use OAI21X1  _7139_
timestamp 0
transform -1 0 10950 0 -1 2170
box -6 -8 106 248
use MUX2X1  _7140_
timestamp 0
transform 1 0 10790 0 1 2170
box -6 -8 126 248
use INVX1  _7141_
timestamp 0
transform -1 0 9370 0 -1 2650
box -6 -8 66 248
use NAND2X1  _7142_
timestamp 0
transform -1 0 9090 0 -1 2650
box -6 -8 86 248
use OAI21X1  _7143_
timestamp 0
transform -1 0 9250 0 -1 2650
box -6 -8 106 248
use INVX1  _7144_
timestamp 0
transform -1 0 9330 0 -1 3130
box -6 -8 66 248
use NAND2X1  _7145_
timestamp 0
transform 1 0 9730 0 1 2650
box -6 -8 86 248
use OAI21X1  _7146_
timestamp 0
transform 1 0 9590 0 1 2650
box -6 -8 106 248
use MUX2X1  _7147_
timestamp 0
transform 1 0 9550 0 -1 2650
box -6 -8 126 248
use MUX2X1  _7148_
timestamp 0
transform -1 0 10130 0 1 2170
box -6 -8 126 248
use NOR2X1  _7149_
timestamp 0
transform 1 0 8370 0 -1 3130
box -6 -8 86 248
use NAND2X1  _7150_
timestamp 0
transform 1 0 8930 0 1 2650
box -6 -8 86 248
use INVX1  _7151_
timestamp 0
transform -1 0 7930 0 1 3130
box -6 -8 66 248
use NAND2X1  _7152_
timestamp 0
transform -1 0 9830 0 1 2170
box -6 -8 86 248
use OAI21X1  _7153_
timestamp 0
transform 1 0 9770 0 1 3610
box -6 -8 106 248
use INVX2  _7154_
timestamp 0
transform 1 0 11030 0 1 3610
box -6 -8 66 248
use OAI21X1  _7155_
timestamp 0
transform 1 0 7990 0 1 3130
box -6 -8 106 248
use OAI21X1  _7156_
timestamp 0
transform 1 0 7570 0 -1 4090
box -6 -8 106 248
use INVX8  _7157_
timestamp 0
transform -1 0 6610 0 1 4570
box -6 -8 126 248
use NAND2X1  _7158_
timestamp 0
transform -1 0 6570 0 1 3610
box -6 -8 86 248
use NOR2X1  _7159_
timestamp 0
transform 1 0 9350 0 1 2650
box -6 -8 86 248
use MUX2X1  _7160_
timestamp 0
transform -1 0 10310 0 -1 2170
box -6 -8 126 248
use MUX2X1  _7161_
timestamp 0
transform -1 0 10130 0 -1 2170
box -6 -8 126 248
use MUX2X1  _7162_
timestamp 0
transform 1 0 9230 0 -1 2170
box -6 -8 126 248
use INVX2  _7163_
timestamp 0
transform 1 0 7990 0 -1 4090
box -6 -8 66 248
use NAND2X1  _7164_
timestamp 0
transform -1 0 8690 0 -1 3130
box -6 -8 86 248
use AOI21X1  _7165_
timestamp 0
transform 1 0 8690 0 -1 2650
box -6 -8 106 248
use NAND3X1  _7166_
timestamp 0
transform 1 0 8850 0 -1 3130
box -6 -8 106 248
use NAND3X1  _7167_
timestamp 0
transform -1 0 9310 0 1 2650
box -6 -8 106 248
use NAND3X1  _7168_
timestamp 0
transform -1 0 9150 0 1 2650
box -6 -8 106 248
use OAI22X1  _7169_
timestamp 0
transform 1 0 8850 0 -1 2650
box -6 -8 126 248
use INVX1  _7170_
timestamp 0
transform -1 0 7670 0 -1 3610
box -6 -8 66 248
use INVX8  _7171_
timestamp 0
transform -1 0 8750 0 -1 1210
box -6 -8 126 248
use INVX1  _7172_
timestamp 0
transform 1 0 11170 0 1 1690
box -6 -8 66 248
use NAND2X1  _7173_
timestamp 0
transform -1 0 9830 0 1 1690
box -6 -8 86 248
use OAI21X1  _7174_
timestamp 0
transform -1 0 9990 0 1 1690
box -6 -8 106 248
use INVX1  _7175_
timestamp 0
transform 1 0 8330 0 -1 1690
box -6 -8 66 248
use NAND2X1  _7176_
timestamp 0
transform 1 0 8510 0 1 1210
box -6 -8 86 248
use OAI21X1  _7177_
timestamp 0
transform 1 0 8370 0 1 1210
box -6 -8 106 248
use MUX2X1  _7178_
timestamp 0
transform -1 0 8490 0 1 1690
box -6 -8 126 248
use INVX1  _7179_
timestamp 0
transform 1 0 10370 0 -1 2170
box -6 -8 66 248
use NAND2X1  _7180_
timestamp 0
transform 1 0 9310 0 1 1690
box -6 -8 86 248
use OAI21X1  _7181_
timestamp 0
transform 1 0 9170 0 1 1690
box -6 -8 106 248
use INVX1  _7182_
timestamp 0
transform 1 0 9470 0 1 2650
box -6 -8 66 248
use NAND2X1  _7183_
timestamp 0
transform 1 0 8870 0 1 1690
box -6 -8 86 248
use OAI21X1  _7184_
timestamp 0
transform -1 0 9110 0 1 1690
box -6 -8 106 248
use MUX2X1  _7185_
timestamp 0
transform 1 0 8710 0 1 1690
box -6 -8 126 248
use MUX2X1  _7186_
timestamp 0
transform 1 0 8550 0 1 1690
box -6 -8 126 248
use NAND3X1  _7187_
timestamp 0
transform -1 0 8490 0 -1 2650
box -6 -8 106 248
use MUX2X1  _7188_
timestamp 0
transform -1 0 8130 0 -1 1690
box -6 -8 126 248
use MUX2X1  _7189_
timestamp 0
transform -1 0 8290 0 -1 1690
box -6 -8 126 248
use MUX2X1  _7190_
timestamp 0
transform 1 0 7830 0 -1 1690
box -6 -8 126 248
use MUX2X1  _7191_
timestamp 0
transform 1 0 10370 0 1 2170
box -6 -8 126 248
use MUX2X1  _7192_
timestamp 0
transform 1 0 9830 0 -1 2650
box -6 -8 126 248
use MUX2X1  _7193_
timestamp 0
transform -1 0 10310 0 1 2170
box -6 -8 126 248
use MUX2X1  _7194_
timestamp 0
transform 1 0 9590 0 1 2170
box -6 -8 126 248
use OAI21X1  _7195_
timestamp 0
transform 1 0 8530 0 -1 2650
box -6 -8 106 248
use AOI21X1  _7196_
timestamp 0
transform -1 0 8070 0 -1 2650
box -6 -8 106 248
use INVX1  _7197_
timestamp 0
transform 1 0 8110 0 1 2650
box -6 -8 66 248
use NAND3X1  _7198_
timestamp 0
transform 1 0 8130 0 -1 2650
box -6 -8 106 248
use AND2X2  _7199_
timestamp 0
transform 1 0 8210 0 1 2650
box -6 -8 106 248
use OAI21X1  _7200_
timestamp 0
transform 1 0 8490 0 1 2650
box -6 -8 106 248
use OR2X2  _7201_
timestamp 0
transform 1 0 8770 0 1 2650
box -6 -8 106 248
use AOI21X1  _7202_
timestamp 0
transform -1 0 8730 0 1 2650
box -6 -8 106 248
use OAI21X1  _7203_
timestamp 0
transform -1 0 6730 0 1 3610
box -6 -8 106 248
use INVX1  _7204_
timestamp 0
transform 1 0 7770 0 -1 6490
box -6 -8 66 248
use NAND2X1  _7205_
timestamp 0
transform 1 0 9430 0 -1 4570
box -6 -8 86 248
use OAI21X1  _7206_
timestamp 0
transform 1 0 7970 0 1 6010
box -6 -8 106 248
use NAND2X1  _7207_
timestamp 0
transform -1 0 6430 0 1 3610
box -6 -8 86 248
use AOI21X1  _7208_
timestamp 0
transform -1 0 7910 0 -1 2650
box -6 -8 106 248
use MUX2X1  _7209_
timestamp 0
transform -1 0 9970 0 -1 2170
box -6 -8 126 248
use MUX2X1  _7210_
timestamp 0
transform -1 0 9030 0 -1 2170
box -6 -8 126 248
use MUX2X1  _7211_
timestamp 0
transform -1 0 9810 0 -1 2170
box -6 -8 126 248
use NAND2X1  _7212_
timestamp 0
transform -1 0 9490 0 -1 2170
box -6 -8 86 248
use OAI22X1  _7213_
timestamp 0
transform 1 0 9530 0 -1 2170
box -6 -8 126 248
use AOI21X1  _7214_
timestamp 0
transform 1 0 9070 0 -1 2170
box -6 -8 106 248
use AOI21X1  _7215_
timestamp 0
transform 1 0 8930 0 1 2170
box -6 -8 106 248
use NAND2X1  _7216_
timestamp 0
transform 1 0 9070 0 1 2170
box -6 -8 86 248
use INVX1  _7217_
timestamp 0
transform 1 0 9210 0 1 2170
box -6 -8 66 248
use OAI21X1  _7218_
timestamp 0
transform 1 0 9450 0 1 2170
box -6 -8 106 248
use NAND2X1  _7219_
timestamp 0
transform 1 0 9330 0 1 2170
box -6 -8 86 248
use AOI21X1  _7220_
timestamp 0
transform -1 0 8730 0 1 2170
box -6 -8 106 248
use NAND3X1  _7221_
timestamp 0
transform 1 0 8770 0 1 2170
box -6 -8 106 248
use INVX1  _7222_
timestamp 0
transform -1 0 8430 0 1 2650
box -6 -8 66 248
use OR2X2  _7223_
timestamp 0
transform -1 0 7930 0 1 2650
box -6 -8 106 248
use NOR2X1  _7224_
timestamp 0
transform -1 0 7790 0 1 2650
box -6 -8 86 248
use INVX1  _7225_
timestamp 0
transform -1 0 7650 0 1 2650
box -6 -8 66 248
use OAI21X1  _7226_
timestamp 0
transform 1 0 7970 0 1 2650
box -6 -8 106 248
use AOI21X1  _7227_
timestamp 0
transform -1 0 7550 0 1 2650
box -6 -8 106 248
use INVX2  _7228_
timestamp 0
transform -1 0 7790 0 -1 1690
box -6 -8 66 248
use OAI21X1  _7229_
timestamp 0
transform -1 0 6250 0 -1 3610
box -6 -8 106 248
use OAI21X1  _7230_
timestamp 0
transform 1 0 6390 0 -1 3610
box -6 -8 106 248
use INVX1  _7231_
timestamp 0
transform -1 0 5990 0 1 3130
box -6 -8 66 248
use INVX2  _7232_
timestamp 0
transform 1 0 6290 0 -1 3610
box -6 -8 66 248
use OAI21X1  _7233_
timestamp 0
transform 1 0 8490 0 1 2170
box -6 -8 106 248
use INVX1  _7234_
timestamp 0
transform 1 0 8390 0 1 2170
box -6 -8 66 248
use INVX1  _7235_
timestamp 0
transform -1 0 7010 0 -1 1210
box -6 -8 66 248
use NAND3X1  _7236_
timestamp 0
transform -1 0 8850 0 -1 2170
box -6 -8 106 248
use INVX1  _7237_
timestamp 0
transform 1 0 11270 0 -1 2170
box -6 -8 66 248
use NAND2X1  _7238_
timestamp 0
transform -1 0 9410 0 -1 1690
box -6 -8 86 248
use OAI21X1  _7239_
timestamp 0
transform -1 0 9570 0 -1 1690
box -6 -8 106 248
use NAND2X1  _7240_
timestamp 0
transform 1 0 7810 0 1 1210
box -6 -8 86 248
use OAI21X1  _7241_
timestamp 0
transform 1 0 7670 0 1 1210
box -6 -8 106 248
use NOR2X1  _7242_
timestamp 0
transform 1 0 7990 0 -1 730
box -6 -8 86 248
use NOR2X1  _7243_
timestamp 0
transform -1 0 8190 0 1 3610
box -6 -8 86 248
use AOI22X1  _7244_
timestamp 0
transform -1 0 8310 0 1 1210
box -6 -8 126 248
use OAI21X1  _7245_
timestamp 0
transform 1 0 7330 0 -1 1210
box -6 -8 106 248
use NAND3X1  _7246_
timestamp 0
transform -1 0 6590 0 -1 1210
box -6 -8 106 248
use INVX1  _7247_
timestamp 0
transform 1 0 6390 0 -1 730
box -6 -8 66 248
use INVX1  _7248_
timestamp 0
transform 1 0 6550 0 1 730
box -6 -8 66 248
use OAI21X1  _7249_
timestamp 0
transform 1 0 6390 0 1 730
box -6 -8 106 248
use NAND3X1  _7250_
timestamp 0
transform -1 0 6290 0 -1 1210
box -6 -8 106 248
use AOI21X1  _7251_
timestamp 0
transform -1 0 6430 0 -1 1210
box -6 -8 106 248
use INVX1  _7252_
timestamp 0
transform 1 0 6430 0 1 1210
box -6 -8 66 248
use NAND2X1  _7253_
timestamp 0
transform 1 0 6450 0 -1 1690
box -6 -8 86 248
use AOI21X1  _7254_
timestamp 0
transform 1 0 8230 0 1 2170
box -6 -8 106 248
use OAI21X1  _7255_
timestamp 0
transform -1 0 8190 0 1 2170
box -6 -8 106 248
use AOI22X1  _7256_
timestamp 0
transform 1 0 6290 0 -1 3130
box -6 -8 126 248
use AOI21X1  _7257_
timestamp 0
transform -1 0 6390 0 1 1210
box -6 -8 106 248
use INVX1  _7258_
timestamp 0
transform -1 0 5850 0 -1 250
box -6 -8 66 248
use INVX1  _7259_
timestamp 0
transform -1 0 9890 0 1 1210
box -6 -8 66 248
use NAND2X1  _7260_
timestamp 0
transform -1 0 8030 0 1 730
box -6 -8 86 248
use OAI21X1  _7261_
timestamp 0
transform -1 0 8150 0 1 1210
box -6 -8 106 248
use NAND2X1  _7262_
timestamp 0
transform -1 0 8330 0 1 1690
box -6 -8 86 248
use OAI21X1  _7263_
timestamp 0
transform 1 0 7590 0 -1 1690
box -6 -8 106 248
use NAND2X1  _7264_
timestamp 0
transform -1 0 8050 0 1 1690
box -6 -8 86 248
use OAI21X1  _7265_
timestamp 0
transform -1 0 6790 0 1 1210
box -6 -8 106 248
use INVX2  _7266_
timestamp 0
transform -1 0 6550 0 -1 730
box -6 -8 66 248
use OAI21X1  _7267_
timestamp 0
transform -1 0 5790 0 1 250
box -6 -8 106 248
use OR2X2  _7268_
timestamp 0
transform -1 0 5130 0 -1 250
box -6 -8 106 248
use NOR2X1  _7269_
timestamp 0
transform 1 0 5830 0 1 250
box -6 -8 86 248
use OAI21X1  _7270_
timestamp 0
transform -1 0 5290 0 -1 250
box -6 -8 106 248
use NAND3X1  _7271_
timestamp 0
transform 1 0 4890 0 -1 250
box -6 -8 106 248
use NOR2X1  _7272_
timestamp 0
transform -1 0 5570 0 -1 250
box -6 -8 86 248
use AND2X2  _7273_
timestamp 0
transform 1 0 5330 0 -1 250
box -6 -8 106 248
use OAI21X1  _7274_
timestamp 0
transform 1 0 5630 0 -1 250
box -6 -8 106 248
use NAND2X1  _7275_
timestamp 0
transform -1 0 5710 0 -1 1210
box -6 -8 86 248
use AOI21X1  _7276_
timestamp 0
transform -1 0 6090 0 1 1210
box -6 -8 106 248
use OAI21X1  _7277_
timestamp 0
transform 1 0 5850 0 1 1210
box -6 -8 106 248
use AOI22X1  _7278_
timestamp 0
transform 1 0 5750 0 1 3130
box -6 -8 126 248
use OAI21X1  _7279_
timestamp 0
transform 1 0 6150 0 1 1210
box -6 -8 106 248
use INVX1  _7280_
timestamp 0
transform 1 0 6590 0 1 250
box -6 -8 66 248
use NAND3X1  _7281_
timestamp 0
transform -1 0 6350 0 -1 730
box -6 -8 106 248
use NAND2X1  _7282_
timestamp 0
transform -1 0 7490 0 1 730
box -6 -8 86 248
use INVX1  _7283_
timestamp 0
transform 1 0 7470 0 -1 1210
box -6 -8 66 248
use AOI21X1  _7284_
timestamp 0
transform -1 0 7470 0 1 1210
box -6 -8 106 248
use NAND2X1  _7285_
timestamp 0
transform 1 0 6830 0 1 1210
box -6 -8 86 248
use OAI21X1  _7286_
timestamp 0
transform 1 0 6810 0 -1 1210
box -6 -8 106 248
use NAND3X1  _7287_
timestamp 0
transform -1 0 6190 0 -1 730
box -6 -8 106 248
use NOR3X1  _7288_
timestamp 0
transform -1 0 6770 0 -1 730
box -6 -8 186 248
use INVX1  _7289_
timestamp 0
transform -1 0 5630 0 1 250
box -6 -8 66 248
use OAI21X1  _7290_
timestamp 0
transform -1 0 5750 0 -1 730
box -6 -8 106 248
use NAND3X1  _7291_
timestamp 0
transform -1 0 5910 0 -1 730
box -6 -8 106 248
use AOI21X1  _7292_
timestamp 0
transform 1 0 5950 0 -1 730
box -6 -8 106 248
use INVX1  _7293_
timestamp 0
transform 1 0 5990 0 1 730
box -6 -8 66 248
use NAND2X1  _7294_
timestamp 0
transform 1 0 6050 0 -1 1210
box -6 -8 86 248
use AND2X2  _7295_
timestamp 0
transform -1 0 7910 0 -1 2170
box -6 -8 106 248
use OAI21X1  _7296_
timestamp 0
transform 1 0 7930 0 1 2170
box -6 -8 106 248
use OAI21X1  _7297_
timestamp 0
transform -1 0 7390 0 1 2650
box -6 -8 106 248
use OAI21X1  _7298_
timestamp 0
transform 1 0 6090 0 -1 4090
box -6 -8 106 248
use INVX1  _7299_
timestamp 0
transform 1 0 5410 0 -1 3610
box -6 -8 66 248
use INVX1  _7300_
timestamp 0
transform -1 0 4350 0 -1 250
box -6 -8 66 248
use NAND3X1  _7301_
timestamp 0
transform -1 0 5230 0 1 250
box -6 -8 106 248
use AOI21X1  _7302_
timestamp 0
transform -1 0 7610 0 1 1210
box -6 -8 106 248
use NAND2X1  _7303_
timestamp 0
transform 1 0 7110 0 1 1210
box -6 -8 86 248
use OAI21X1  _7304_
timestamp 0
transform 1 0 6950 0 1 1210
box -6 -8 106 248
use NAND3X1  _7305_
timestamp 0
transform -1 0 4930 0 1 250
box -6 -8 106 248
use INVX1  _7306_
timestamp 0
transform -1 0 4450 0 -1 250
box -6 -8 66 248
use OAI21X1  _7307_
timestamp 0
transform -1 0 5510 0 1 250
box -6 -8 106 248
use NAND2X1  _7308_
timestamp 0
transform -1 0 4230 0 -1 250
box -6 -8 86 248
use NAND3X1  _7309_
timestamp 0
transform 1 0 3990 0 -1 250
box -6 -8 106 248
use NAND3X1  _7310_
timestamp 0
transform -1 0 4770 0 1 250
box -6 -8 106 248
use NAND2X1  _7311_
timestamp 0
transform -1 0 4570 0 -1 250
box -6 -8 86 248
use NAND3X1  _7312_
timestamp 0
transform -1 0 4610 0 1 250
box -6 -8 106 248
use NAND2X1  _7313_
timestamp 0
transform -1 0 4710 0 -1 1210
box -6 -8 86 248
use AOI21X1  _7314_
timestamp 0
transform -1 0 4850 0 -1 250
box -6 -8 106 248
use NOR2X1  _7315_
timestamp 0
transform 1 0 5530 0 -1 730
box -6 -8 86 248
use OAI21X1  _7316_
timestamp 0
transform -1 0 5590 0 -1 1210
box -6 -8 106 248
use NAND2X1  _7317_
timestamp 0
transform -1 0 5450 0 -1 1210
box -6 -8 86 248
use AOI21X1  _7318_
timestamp 0
transform 1 0 5690 0 1 1210
box -6 -8 106 248
use OAI21X1  _7319_
timestamp 0
transform 1 0 5550 0 1 1210
box -6 -8 106 248
use AOI22X1  _7320_
timestamp 0
transform 1 0 5530 0 -1 3610
box -6 -8 126 248
use INVX1  _7321_
timestamp 0
transform 1 0 5230 0 -1 4090
box -6 -8 66 248
use AOI21X1  _7322_
timestamp 0
transform -1 0 3950 0 -1 250
box -6 -8 106 248
use AND2X2  _7323_
timestamp 0
transform 1 0 5830 0 1 730
box -6 -8 106 248
use NAND3X1  _7324_
timestamp 0
transform -1 0 6010 0 -1 1210
box -6 -8 106 248
use AOI21X1  _7325_
timestamp 0
transform 1 0 5690 0 1 730
box -6 -8 106 248
use OAI21X1  _7326_
timestamp 0
transform -1 0 5850 0 -1 1210
box -6 -8 106 248
use AOI21X1  _7327_
timestamp 0
transform -1 0 4870 0 -1 1210
box -6 -8 106 248
use INVX1  _7328_
timestamp 0
transform -1 0 6710 0 1 730
box -6 -8 66 248
use NAND3X1  _7329_
timestamp 0
transform 1 0 5210 0 -1 730
box -6 -8 106 248
use INVX1  _7330_
timestamp 0
transform -1 0 7410 0 -1 730
box -6 -8 66 248
use NOR2X1  _7331_
timestamp 0
transform -1 0 7370 0 1 730
box -6 -8 86 248
use INVX1  _7332_
timestamp 0
transform -1 0 7230 0 1 730
box -6 -8 66 248
use OAI21X1  _7333_
timestamp 0
transform -1 0 7150 0 -1 1210
box -6 -8 106 248
use NAND3X1  _7334_
timestamp 0
transform -1 0 6350 0 1 730
box -6 -8 106 248
use INVX1  _7335_
timestamp 0
transform -1 0 5150 0 -1 730
box -6 -8 66 248
use OAI21X1  _7336_
timestamp 0
transform -1 0 5090 0 1 250
box -6 -8 106 248
use NAND2X1  _7337_
timestamp 0
transform -1 0 5050 0 -1 730
box -6 -8 86 248
use NAND3X1  _7338_
timestamp 0
transform -1 0 6190 0 1 730
box -6 -8 106 248
use NAND3X1  _7339_
timestamp 0
transform 1 0 5370 0 -1 730
box -6 -8 106 248
use NAND2X1  _7340_
timestamp 0
transform 1 0 5570 0 1 730
box -6 -8 86 248
use NAND3X1  _7341_
timestamp 0
transform 1 0 5430 0 1 730
box -6 -8 106 248
use NAND2X1  _7342_
timestamp 0
transform 1 0 5290 0 1 730
box -6 -8 86 248
use INVX1  _7343_
timestamp 0
transform -1 0 5090 0 1 1210
box -6 -8 66 248
use NOR2X1  _7344_
timestamp 0
transform -1 0 4970 0 1 1210
box -6 -8 86 248
use OAI21X1  _7345_
timestamp 0
transform -1 0 5170 0 -1 1210
box -6 -8 106 248
use OAI21X1  _7346_
timestamp 0
transform 1 0 5170 0 -1 1690
box -6 -8 106 248
use OAI21X1  _7347_
timestamp 0
transform -1 0 5370 0 -1 3610
box -6 -8 106 248
use INVX1  _7348_
timestamp 0
transform 1 0 5350 0 -1 3130
box -6 -8 66 248
use OAI21X1  _7349_
timestamp 0
transform 1 0 5290 0 1 1690
box -6 -8 106 248
use OAI21X1  _7350_
timestamp 0
transform 1 0 5330 0 -1 4090
box -6 -8 106 248
use INVX1  _7351_
timestamp 0
transform 1 0 6190 0 -1 3130
box -6 -8 66 248
use OAI21X1  _7352_
timestamp 0
transform 1 0 5210 0 -1 1210
box -6 -8 106 248
use NOR2X1  _7353_
timestamp 0
transform -1 0 5370 0 1 1210
box -6 -8 86 248
use AOI21X1  _7354_
timestamp 0
transform 1 0 5410 0 1 1210
box -6 -8 106 248
use INVX1  _7355_
timestamp 0
transform -1 0 5510 0 1 1690
box -6 -8 66 248
use OR2X2  _7356_
timestamp 0
transform 1 0 5950 0 -1 1690
box -6 -8 106 248
use OAI21X1  _7357_
timestamp 0
transform -1 0 6770 0 -1 1690
box -6 -8 106 248
use NAND3X1  _7358_
timestamp 0
transform -1 0 5950 0 1 1690
box -6 -8 106 248
use NOR2X1  _7359_
timestamp 0
transform -1 0 5630 0 -1 1690
box -6 -8 86 248
use INVX1  _7360_
timestamp 0
transform -1 0 5790 0 1 1690
box -6 -8 66 248
use OAI21X1  _7361_
timestamp 0
transform -1 0 5770 0 -1 1690
box -6 -8 106 248
use NAND3X1  _7362_
timestamp 0
transform 1 0 5570 0 1 1690
box -6 -8 106 248
use NAND3X1  _7363_
timestamp 0
transform 1 0 5990 0 1 1690
box -6 -8 106 248
use OAI21X1  _7364_
timestamp 0
transform 1 0 5810 0 -1 1690
box -6 -8 106 248
use NAND3X1  _7365_
timestamp 0
transform 1 0 6150 0 1 1690
box -6 -8 106 248
use AND2X2  _7366_
timestamp 0
transform 1 0 6830 0 -1 2170
box -6 -8 106 248
use INVX1  _7367_
timestamp 0
transform -1 0 6910 0 1 2170
box -6 -8 66 248
use AOI21X1  _7368_
timestamp 0
transform -1 0 6410 0 -1 2650
box -6 -8 106 248
use OAI21X1  _7369_
timestamp 0
transform -1 0 6270 0 -1 2650
box -6 -8 106 248
use AOI22X1  _7370_
timestamp 0
transform -1 0 6130 0 -1 3130
box -6 -8 126 248
use NAND2X1  _7371_
timestamp 0
transform 1 0 5010 0 1 730
box -6 -8 86 248
use AND2X2  _7372_
timestamp 0
transform -1 0 5030 0 -1 1210
box -6 -8 106 248
use AND2X2  _7373_
timestamp 0
transform 1 0 4830 0 -1 730
box -6 -8 106 248
use NAND3X1  _7374_
timestamp 0
transform 1 0 5150 0 1 730
box -6 -8 106 248
use OAI21X1  _7375_
timestamp 0
transform -1 0 5230 0 1 1210
box -6 -8 106 248
use INVX1  _7376_
timestamp 0
transform 1 0 6970 0 -1 2170
box -6 -8 66 248
use AOI21X1  _7377_
timestamp 0
transform -1 0 6790 0 -1 2170
box -6 -8 106 248
use INVX1  _7378_
timestamp 0
transform 1 0 7950 0 -1 2170
box -6 -8 66 248
use NOR3X1  _7379_
timestamp 0
transform 1 0 6110 0 -1 1690
box -6 -8 186 248
use INVX1  _7380_
timestamp 0
transform -1 0 6390 0 -1 1690
box -6 -8 66 248
use OAI21X1  _7381_
timestamp 0
transform 1 0 6530 0 1 1210
box -6 -8 106 248
use NAND3X1  _7382_
timestamp 0
transform 1 0 6470 0 1 1690
box -6 -8 106 248
use INVX1  _7383_
timestamp 0
transform 1 0 6570 0 -1 1690
box -6 -8 66 248
use OAI21X1  _7384_
timestamp 0
transform 1 0 6630 0 1 1690
box -6 -8 106 248
use NAND3X1  _7385_
timestamp 0
transform -1 0 7610 0 -1 2170
box -6 -8 106 248
use NAND3X1  _7386_
timestamp 0
transform 1 0 6310 0 1 1690
box -6 -8 106 248
use OAI21X1  _7387_
timestamp 0
transform -1 0 6910 0 -1 1690
box -6 -8 106 248
use NAND3X1  _7388_
timestamp 0
transform -1 0 7170 0 -1 2170
box -6 -8 106 248
use AND2X2  _7389_
timestamp 0
transform -1 0 7330 0 -1 2170
box -6 -8 106 248
use AND2X2  _7390_
timestamp 0
transform -1 0 6550 0 -1 2650
box -6 -8 106 248
use OAI21X1  _7391_
timestamp 0
transform -1 0 6610 0 1 2650
box -6 -8 106 248
use OAI21X1  _7392_
timestamp 0
transform -1 0 6450 0 1 2650
box -6 -8 106 248
use OAI21X1  _7393_
timestamp 0
transform -1 0 5190 0 -1 4570
box -6 -8 106 248
use INVX1  _7394_
timestamp 0
transform 1 0 7310 0 1 250
box -6 -8 66 248
use OAI21X1  _7395_
timestamp 0
transform -1 0 7170 0 -1 1690
box -6 -8 106 248
use INVX1  _7396_
timestamp 0
transform -1 0 7150 0 1 1690
box -6 -8 66 248
use AOI21X1  _7397_
timestamp 0
transform 1 0 6930 0 1 1690
box -6 -8 106 248
use NAND3X1  _7398_
timestamp 0
transform 1 0 6790 0 1 1690
box -6 -8 106 248
use NAND2X1  _7399_
timestamp 0
transform 1 0 8330 0 -1 2170
box -6 -8 86 248
use NAND2X1  _7400_
timestamp 0
transform -1 0 7270 0 1 1690
box -6 -8 86 248
use OAI21X1  _7401_
timestamp 0
transform -1 0 7430 0 1 1690
box -6 -8 106 248
use NAND2X1  _7402_
timestamp 0
transform 1 0 7230 0 1 1210
box -6 -8 86 248
use INVX1  _7403_
timestamp 0
transform 1 0 7610 0 1 1690
box -6 -8 66 248
use AND2X2  _7404_
timestamp 0
transform 1 0 8450 0 -1 2170
box -6 -8 106 248
use NAND2X1  _7405_
timestamp 0
transform 1 0 8210 0 -1 2170
box -6 -8 86 248
use NAND3X1  _7406_
timestamp 0
transform 1 0 8050 0 -1 2170
box -6 -8 106 248
use NAND2X1  _7407_
timestamp 0
transform 1 0 7790 0 1 2170
box -6 -8 86 248
use AOI21X1  _7408_
timestamp 0
transform 1 0 7670 0 -1 2170
box -6 -8 106 248
use AOI21X1  _7409_
timestamp 0
transform 1 0 7370 0 -1 2170
box -6 -8 106 248
use NAND3X1  _7410_
timestamp 0
transform 1 0 7230 0 1 2170
box -6 -8 106 248
use AOI21X1  _7411_
timestamp 0
transform 1 0 7650 0 1 2170
box -6 -8 106 248
use AND2X2  _7412_
timestamp 0
transform 1 0 6990 0 -1 2650
box -6 -8 106 248
use NAND3X1  _7413_
timestamp 0
transform 1 0 7370 0 1 2170
box -6 -8 106 248
use OAI21X1  _7414_
timestamp 0
transform 1 0 7510 0 1 2170
box -6 -8 106 248
use OAI21X1  _7415_
timestamp 0
transform 1 0 7150 0 -1 2650
box -6 -8 106 248
use OR2X2  _7416_
timestamp 0
transform -1 0 7250 0 1 2650
box -6 -8 106 248
use AOI22X1  _7417_
timestamp 0
transform 1 0 5970 0 -1 3610
box -6 -8 126 248
use NAND2X1  _7418_
timestamp 0
transform -1 0 5530 0 1 3610
box -6 -8 86 248
use INVX1  _7419_
timestamp 0
transform -1 0 6930 0 -1 2650
box -6 -8 66 248
use NAND2X1  _7420_
timestamp 0
transform 1 0 7470 0 -1 730
box -6 -8 86 248
use INVX1  _7421_
timestamp 0
transform 1 0 7050 0 -1 250
box -6 -8 66 248
use NAND2X1  _7422_
timestamp 0
transform 1 0 7690 0 1 250
box -6 -8 86 248
use NAND2X1  _7423_
timestamp 0
transform 1 0 7590 0 -1 730
box -6 -8 86 248
use INVX1  _7424_
timestamp 0
transform -1 0 7750 0 -1 2650
box -6 -8 66 248
use NAND2X1  _7425_
timestamp 0
transform 1 0 7430 0 -1 2650
box -6 -8 86 248
use NAND2X1  _7426_
timestamp 0
transform -1 0 7630 0 -1 2650
box -6 -8 86 248
use NAND2X1  _7427_
timestamp 0
transform -1 0 7390 0 -1 2650
box -6 -8 86 248
use INVX1  _7428_
timestamp 0
transform 1 0 7050 0 1 2650
box -6 -8 66 248
use NOR3X1  _7429_
timestamp 0
transform -1 0 7010 0 1 2650
box -6 -8 186 248
use AOI21X1  _7430_
timestamp 0
transform -1 0 6830 0 -1 2650
box -6 -8 106 248
use OAI21X1  _7431_
timestamp 0
transform -1 0 6690 0 -1 2650
box -6 -8 106 248
use OAI21X1  _7432_
timestamp 0
transform -1 0 6770 0 1 2650
box -6 -8 106 248
use NAND2X1  _7433_
timestamp 0
transform 1 0 5610 0 -1 4090
box -6 -8 86 248
use NAND2X1  _7434_
timestamp 0
transform 1 0 8250 0 1 3610
box -6 -8 86 248
use INVX1  _7435_
timestamp 0
transform 1 0 7490 0 -1 1690
box -6 -8 66 248
use NAND2X1  _7436_
timestamp 0
transform -1 0 7310 0 -1 1690
box -6 -8 86 248
use OAI21X1  _7437_
timestamp 0
transform -1 0 7450 0 -1 1690
box -6 -8 106 248
use NAND2X1  _7438_
timestamp 0
transform -1 0 7650 0 -1 1210
box -6 -8 86 248
use NOR2X1  _7439_
timestamp 0
transform 1 0 8070 0 -1 3610
box -6 -8 86 248
use NOR2X1  _7440_
timestamp 0
transform 1 0 7190 0 1 3610
box -6 -8 86 248
use AOI22X1  _7441_
timestamp 0
transform -1 0 7850 0 -1 3610
box -6 -8 126 248
use NAND3X1  _7442_
timestamp 0
transform 1 0 7690 0 -1 1210
box -6 -8 106 248
use NAND2X1  _7443_
timestamp 0
transform 1 0 5290 0 1 250
box -6 -8 86 248
use OAI21X1  _7444_
timestamp 0
transform -1 0 4710 0 -1 250
box -6 -8 106 248
use NAND2X1  _7445_
timestamp 0
transform 1 0 6550 0 -1 250
box -6 -8 86 248
use OAI21X1  _7446_
timestamp 0
transform 1 0 6410 0 -1 250
box -6 -8 106 248
use MUX2X1  _7447_
timestamp 0
transform -1 0 7810 0 -1 250
box -6 -8 126 248
use NAND2X1  _7448_
timestamp 0
transform 1 0 8270 0 -1 250
box -6 -8 86 248
use AND2X2  _7449_
timestamp 0
transform 1 0 8790 0 -1 1210
box -6 -8 106 248
use NOR2X1  _7450_
timestamp 0
transform -1 0 8810 0 -1 3130
box -6 -8 86 248
use NAND2X1  _7451_
timestamp 0
transform -1 0 8170 0 1 250
box -6 -8 86 248
use NAND2X1  _7452_
timestamp 0
transform -1 0 7650 0 -1 250
box -6 -8 86 248
use NAND2X1  _7453_
timestamp 0
transform 1 0 8230 0 1 250
box -6 -8 86 248
use OAI21X1  _7454_
timestamp 0
transform 1 0 8330 0 -1 1210
box -6 -8 106 248
use OAI21X1  _7455_
timestamp 0
transform -1 0 10170 0 -1 3130
box -6 -8 106 248
use OAI21X1  _7456_
timestamp 0
transform -1 0 8710 0 1 3610
box -6 -8 106 248
use NAND2X1  _7457_
timestamp 0
transform -1 0 8590 0 -1 4090
box -6 -8 86 248
use NOR2X1  _7458_
timestamp 0
transform 1 0 10390 0 1 2650
box -6 -8 86 248
use NAND2X1  _7459_
timestamp 0
transform -1 0 6030 0 1 250
box -6 -8 86 248
use OAI21X1  _7460_
timestamp 0
transform -1 0 6750 0 -1 1210
box -6 -8 106 248
use NAND2X1  _7461_
timestamp 0
transform -1 0 7790 0 1 1690
box -6 -8 86 248
use OAI21X1  _7462_
timestamp 0
transform -1 0 7930 0 1 1690
box -6 -8 106 248
use MUX2X1  _7463_
timestamp 0
transform 1 0 8090 0 1 730
box -6 -8 126 248
use NAND2X1  _7464_
timestamp 0
transform 1 0 8430 0 1 730
box -6 -8 86 248
use NAND2X1  _7465_
timestamp 0
transform 1 0 6910 0 1 730
box -6 -8 86 248
use OAI21X1  _7466_
timestamp 0
transform 1 0 6750 0 1 730
box -6 -8 106 248
use INVX1  _7467_
timestamp 0
transform 1 0 8530 0 -1 730
box -6 -8 66 248
use NAND2X1  _7468_
timestamp 0
transform -1 0 6890 0 -1 730
box -6 -8 86 248
use OAI21X1  _7469_
timestamp 0
transform -1 0 7030 0 -1 730
box -6 -8 106 248
use NAND2X1  _7470_
timestamp 0
transform -1 0 8330 0 -1 730
box -6 -8 86 248
use OAI21X1  _7471_
timestamp 0
transform 1 0 8370 0 -1 730
box -6 -8 106 248
use OAI21X1  _7472_
timestamp 0
transform -1 0 8830 0 1 730
box -6 -8 106 248
use NAND3X1  _7473_
timestamp 0
transform -1 0 9290 0 -1 1690
box -6 -8 106 248
use MUX2X1  _7474_
timestamp 0
transform -1 0 8390 0 1 730
box -6 -8 126 248
use MUX2X1  _7475_
timestamp 0
transform 1 0 8550 0 1 730
box -6 -8 126 248
use OAI21X1  _7476_
timestamp 0
transform -1 0 9150 0 -1 1690
box -6 -8 106 248
use AOI21X1  _7477_
timestamp 0
transform 1 0 9610 0 1 1690
box -6 -8 106 248
use INVX1  _7478_
timestamp 0
transform -1 0 11150 0 1 2170
box -6 -8 66 248
use NAND3X1  _7479_
timestamp 0
transform 1 0 9450 0 1 1690
box -6 -8 106 248
use AND2X2  _7480_
timestamp 0
transform -1 0 11050 0 1 2170
box -6 -8 106 248
use NAND2X1  _7481_
timestamp 0
transform -1 0 10230 0 -1 2650
box -6 -8 86 248
use OR2X2  _7482_
timestamp 0
transform -1 0 10110 0 -1 2650
box -6 -8 106 248
use AOI21X1  _7483_
timestamp 0
transform -1 0 9510 0 -1 2650
box -6 -8 106 248
use OAI21X1  _7484_
timestamp 0
transform -1 0 8750 0 -1 4090
box -6 -8 106 248
use NAND2X1  _7485_
timestamp 0
transform -1 0 8830 0 1 3610
box -6 -8 86 248
use AOI21X1  _7486_
timestamp 0
transform 1 0 11210 0 1 2170
box -6 -8 106 248
use NAND2X1  _7487_
timestamp 0
transform -1 0 9350 0 1 1210
box -6 -8 86 248
use NAND2X1  _7488_
timestamp 0
transform -1 0 7730 0 1 730
box -6 -8 86 248
use OAI21X1  _7489_
timestamp 0
transform -1 0 7890 0 1 730
box -6 -8 106 248
use NAND2X1  _7490_
timestamp 0
transform -1 0 7930 0 -1 250
box -6 -8 86 248
use OAI21X1  _7491_
timestamp 0
transform 1 0 8370 0 1 250
box -6 -8 106 248
use NAND2X1  _7492_
timestamp 0
transform 1 0 7830 0 -1 1210
box -6 -8 86 248
use NAND2X1  _7493_
timestamp 0
transform 1 0 7950 0 1 250
box -6 -8 86 248
use NAND2X1  _7494_
timestamp 0
transform -1 0 7910 0 1 250
box -6 -8 86 248
use AOI21X1  _7495_
timestamp 0
transform 1 0 8650 0 1 250
box -6 -8 106 248
use INVX1  _7496_
timestamp 0
transform -1 0 9150 0 -1 1210
box -6 -8 66 248
use NAND3X1  _7497_
timestamp 0
transform 1 0 9530 0 1 1210
box -6 -8 106 248
use AOI21X1  _7498_
timestamp 0
transform 1 0 8890 0 1 730
box -6 -8 106 248
use OAI21X1  _7499_
timestamp 0
transform -1 0 9030 0 -1 1210
box -6 -8 106 248
use NAND3X1  _7500_
timestamp 0
transform 1 0 10170 0 1 1690
box -6 -8 106 248
use INVX1  _7501_
timestamp 0
transform -1 0 11730 0 -1 2170
box -6 -8 66 248
use AOI21X1  _7502_
timestamp 0
transform 1 0 10030 0 1 1690
box -6 -8 106 248
use NOR2X1  _7503_
timestamp 0
transform 1 0 11650 0 1 2170
box -6 -8 86 248
use AND2X2  _7504_
timestamp 0
transform -1 0 11450 0 1 2170
box -6 -8 106 248
use NOR2X1  _7505_
timestamp 0
transform 1 0 11510 0 1 2170
box -6 -8 86 248
use OAI21X1  _7506_
timestamp 0
transform -1 0 11030 0 -1 2650
box -6 -8 106 248
use OAI21X1  _7507_
timestamp 0
transform -1 0 8970 0 1 3610
box -6 -8 106 248
use OAI21X1  _7508_
timestamp 0
transform 1 0 11790 0 1 2170
box -6 -8 106 248
use INVX1  _7509_
timestamp 0
transform 1 0 12230 0 1 2170
box -6 -8 66 248
use NAND2X1  _7510_
timestamp 0
transform -1 0 7810 0 -1 730
box -6 -8 86 248
use OAI21X1  _7511_
timestamp 0
transform -1 0 7950 0 -1 730
box -6 -8 106 248
use MUX2X1  _7512_
timestamp 0
transform 1 0 8630 0 -1 730
box -6 -8 126 248
use NOR2X1  _7513_
timestamp 0
transform 1 0 9070 0 -1 730
box -6 -8 86 248
use NAND2X1  _7514_
timestamp 0
transform -1 0 8170 0 -1 1210
box -6 -8 86 248
use NAND2X1  _7515_
timestamp 0
transform -1 0 8050 0 -1 1210
box -6 -8 86 248
use NAND2X1  _7516_
timestamp 0
transform -1 0 8290 0 -1 1210
box -6 -8 86 248
use OR2X2  _7517_
timestamp 0
transform 1 0 9210 0 -1 1210
box -6 -8 106 248
use OAI21X1  _7518_
timestamp 0
transform -1 0 9490 0 1 1210
box -6 -8 106 248
use OR2X2  _7519_
timestamp 0
transform 1 0 10170 0 1 1210
box -6 -8 106 248
use OAI21X1  _7520_
timestamp 0
transform 1 0 9370 0 -1 1210
box -6 -8 106 248
use AOI21X1  _7521_
timestamp 0
transform 1 0 11370 0 -1 2170
box -6 -8 106 248
use INVX1  _7522_
timestamp 0
transform 1 0 12150 0 -1 2170
box -6 -8 66 248
use NAND3X1  _7523_
timestamp 0
transform 1 0 11510 0 -1 2170
box -6 -8 106 248
use NAND2X1  _7524_
timestamp 0
transform 1 0 12270 0 -1 2170
box -6 -8 86 248
use OR2X2  _7525_
timestamp 0
transform 1 0 12450 0 1 2170
box -6 -8 106 248
use NAND2X1  _7526_
timestamp 0
transform -1 0 12410 0 1 2170
box -6 -8 86 248
use NAND2X1  _7527_
timestamp 0
transform 1 0 12610 0 1 2170
box -6 -8 86 248
use AOI22X1  _7528_
timestamp 0
transform 1 0 9790 0 -1 3610
box -6 -8 126 248
use AOI21X1  _7529_
timestamp 0
transform -1 0 12050 0 1 2170
box -6 -8 106 248
use NAND2X1  _7530_
timestamp 0
transform -1 0 7490 0 1 250
box -6 -8 86 248
use OAI21X1  _7531_
timestamp 0
transform -1 0 7630 0 1 250
box -6 -8 106 248
use NAND2X1  _7532_
timestamp 0
transform -1 0 8070 0 -1 250
box -6 -8 86 248
use OAI21X1  _7533_
timestamp 0
transform -1 0 8210 0 -1 250
box -6 -8 106 248
use NAND2X1  _7534_
timestamp 0
transform 1 0 8790 0 -1 250
box -6 -8 86 248
use OAI21X1  _7535_
timestamp 0
transform 1 0 8630 0 -1 250
box -6 -8 106 248
use INVX1  _7536_
timestamp 0
transform -1 0 10870 0 -1 1210
box -6 -8 66 248
use NAND3X1  _7537_
timestamp 0
transform 1 0 9130 0 1 1210
box -6 -8 106 248
use OAI21X1  _7538_
timestamp 0
transform 1 0 10830 0 1 1210
box -6 -8 106 248
use OR2X2  _7539_
timestamp 0
transform 1 0 11710 0 1 1690
box -6 -8 106 248
use NOR2X1  _7540_
timestamp 0
transform -1 0 10790 0 1 1210
box -6 -8 86 248
use OAI21X1  _7541_
timestamp 0
transform -1 0 11270 0 -1 1690
box -6 -8 106 248
use NAND3X1  _7542_
timestamp 0
transform 1 0 11850 0 1 1690
box -6 -8 106 248
use OR2X2  _7543_
timestamp 0
transform 1 0 11470 0 -1 1690
box -6 -8 106 248
use OAI21X1  _7544_
timestamp 0
transform 1 0 11330 0 -1 1690
box -6 -8 106 248
use NAND3X1  _7545_
timestamp 0
transform 1 0 12930 0 -1 2170
box -6 -8 106 248
use NAND2X1  _7546_
timestamp 0
transform 1 0 12670 0 -1 2650
box -6 -8 86 248
use OR2X2  _7547_
timestamp 0
transform -1 0 12610 0 1 2650
box -6 -8 106 248
use NAND2X1  _7548_
timestamp 0
transform 1 0 12670 0 1 2650
box -6 -8 86 248
use NAND2X1  _7549_
timestamp 0
transform -1 0 12550 0 -1 3130
box -6 -8 86 248
use AOI22X1  _7550_
timestamp 0
transform 1 0 11150 0 1 3130
box -6 -8 126 248
use INVX1  _7551_
timestamp 0
transform -1 0 9770 0 -1 4090
box -6 -8 66 248
use OAI21X1  _7552_
timestamp 0
transform -1 0 11970 0 -1 2650
box -6 -8 106 248
use NAND2X1  _7553_
timestamp 0
transform 1 0 11130 0 1 1210
box -6 -8 86 248
use NOR2X1  _7554_
timestamp 0
transform -1 0 8470 0 -1 250
box -6 -8 86 248
use AOI21X1  _7555_
timestamp 0
transform 1 0 8810 0 1 250
box -6 -8 106 248
use NAND2X1  _7556_
timestamp 0
transform -1 0 8870 0 -1 730
box -6 -8 86 248
use OAI21X1  _7557_
timestamp 0
transform -1 0 9010 0 -1 730
box -6 -8 106 248
use INVX1  _7558_
timestamp 0
transform 1 0 10450 0 1 730
box -6 -8 66 248
use NAND3X1  _7559_
timestamp 0
transform 1 0 10970 0 1 1210
box -6 -8 106 248
use NOR2X1  _7560_
timestamp 0
transform 1 0 9310 0 1 730
box -6 -8 86 248
use NAND3X1  _7561_
timestamp 0
transform 1 0 9150 0 1 730
box -6 -8 106 248
use OAI21X1  _7562_
timestamp 0
transform 1 0 10150 0 1 730
box -6 -8 106 248
use NAND2X1  _7563_
timestamp 0
transform -1 0 10390 0 1 730
box -6 -8 86 248
use AOI21X1  _7564_
timestamp 0
transform 1 0 11010 0 -1 1690
box -6 -8 106 248
use INVX1  _7565_
timestamp 0
transform 1 0 13730 0 1 2170
box -6 -8 66 248
use NAND3X1  _7566_
timestamp 0
transform 1 0 10870 0 -1 1690
box -6 -8 106 248
use NAND2X1  _7567_
timestamp 0
transform 1 0 13590 0 1 2170
box -6 -8 86 248
use NOR2X1  _7568_
timestamp 0
transform -1 0 11810 0 1 3130
box -6 -8 86 248
use AND2X2  _7569_
timestamp 0
transform -1 0 11850 0 -1 3130
box -6 -8 106 248
use OAI21X1  _7570_
timestamp 0
transform -1 0 11690 0 1 3130
box -6 -8 106 248
use OAI21X1  _7571_
timestamp 0
transform 1 0 10050 0 -1 4090
box -6 -8 106 248
use INVX1  _7572_
timestamp 0
transform 1 0 9150 0 -1 4570
box -6 -8 66 248
use NAND3X1  _7573_
timestamp 0
transform -1 0 10630 0 -1 1210
box -6 -8 106 248
use AOI21X1  _7574_
timestamp 0
transform 1 0 8950 0 1 250
box -6 -8 106 248
use NAND2X1  _7575_
timestamp 0
transform 1 0 9510 0 1 250
box -6 -8 86 248
use OAI21X1  _7576_
timestamp 0
transform 1 0 9630 0 1 250
box -6 -8 106 248
use NAND3X1  _7577_
timestamp 0
transform 1 0 10390 0 -1 1210
box -6 -8 106 248
use NOR3X1  _7578_
timestamp 0
transform 1 0 9530 0 1 730
box -6 -8 186 248
use INVX1  _7579_
timestamp 0
transform -1 0 9710 0 -1 730
box -6 -8 66 248
use OAI21X1  _7580_
timestamp 0
transform 1 0 9790 0 -1 1210
box -6 -8 106 248
use NAND2X1  _7581_
timestamp 0
transform 1 0 12530 0 -1 2170
box -6 -8 86 248
use NAND2X1  _7582_
timestamp 0
transform -1 0 13090 0 1 2170
box -6 -8 86 248
use NAND3X1  _7583_
timestamp 0
transform -1 0 12490 0 -1 2170
box -6 -8 106 248
use NAND2X1  _7584_
timestamp 0
transform -1 0 12110 0 -1 2650
box -6 -8 86 248
use AOI21X1  _7585_
timestamp 0
transform -1 0 12890 0 -1 2170
box -6 -8 106 248
use NOR2X1  _7586_
timestamp 0
transform -1 0 12750 0 -1 2170
box -6 -8 86 248
use OAI21X1  _7587_
timestamp 0
transform 1 0 12270 0 -1 2650
box -6 -8 106 248
use NAND2X1  _7588_
timestamp 0
transform -1 0 12230 0 -1 2650
box -6 -8 86 248
use NOR2X1  _7589_
timestamp 0
transform 1 0 12110 0 1 2650
box -6 -8 86 248
use AND2X2  _7590_
timestamp 0
transform -1 0 11830 0 -1 2650
box -6 -8 106 248
use AND2X2  _7591_
timestamp 0
transform 1 0 13990 0 1 2170
box -6 -8 106 248
use NAND3X1  _7592_
timestamp 0
transform 1 0 13830 0 1 2170
box -6 -8 106 248
use AOI21X1  _7593_
timestamp 0
transform 1 0 13430 0 -1 2170
box -6 -8 106 248
use OAI21X1  _7594_
timestamp 0
transform 1 0 13430 0 1 2170
box -6 -8 106 248
use NOR2X1  _7595_
timestamp 0
transform -1 0 11690 0 -1 2650
box -6 -8 86 248
use OAI21X1  _7596_
timestamp 0
transform -1 0 10870 0 -1 3610
box -6 -8 106 248
use NAND2X1  _7597_
timestamp 0
transform 1 0 10250 0 1 3610
box -6 -8 86 248
use OAI21X1  _7598_
timestamp 0
transform 1 0 9270 0 -1 4570
box -6 -8 106 248
use INVX1  _7599_
timestamp 0
transform 1 0 10190 0 -1 4090
box -6 -8 66 248
use INVX1  _7600_
timestamp 0
transform 1 0 11890 0 -1 3130
box -6 -8 66 248
use NAND2X1  _7601_
timestamp 0
transform -1 0 9750 0 -1 1210
box -6 -8 86 248
use NOR2X1  _7602_
timestamp 0
transform 1 0 9090 0 1 250
box -6 -8 86 248
use INVX1  _7603_
timestamp 0
transform 1 0 9230 0 1 250
box -6 -8 66 248
use OAI21X1  _7604_
timestamp 0
transform 1 0 9330 0 -1 730
box -6 -8 106 248
use NAND3X1  _7605_
timestamp 0
transform 1 0 10430 0 1 1210
box -6 -8 106 248
use INVX1  _7606_
timestamp 0
transform 1 0 10050 0 1 730
box -6 -8 66 248
use OAI21X1  _7607_
timestamp 0
transform 1 0 10230 0 -1 1210
box -6 -8 106 248
use NAND2X1  _7608_
timestamp 0
transform 1 0 10110 0 -1 1210
box -6 -8 86 248
use NAND3X1  _7609_
timestamp 0
transform 1 0 10490 0 -1 1690
box -6 -8 106 248
use NAND3X1  _7610_
timestamp 0
transform 1 0 9950 0 -1 1210
box -6 -8 106 248
use NAND2X1  _7611_
timestamp 0
transform -1 0 10390 0 1 1210
box -6 -8 86 248
use NAND3X1  _7612_
timestamp 0
transform 1 0 10730 0 1 1690
box -6 -8 106 248
use NAND2X1  _7613_
timestamp 0
transform 1 0 11430 0 1 1690
box -6 -8 86 248
use OAI21X1  _7614_
timestamp 0
transform -1 0 11110 0 -1 3610
box -6 -8 106 248
use NOR2X1  _7615_
timestamp 0
transform 1 0 11170 0 -1 3610
box -6 -8 86 248
use INVX1  _7616_
timestamp 0
transform -1 0 10970 0 -1 3610
box -6 -8 66 248
use AOI21X1  _7617_
timestamp 0
transform -1 0 10990 0 1 3610
box -6 -8 106 248
use AOI22X1  _7618_
timestamp 0
transform 1 0 10710 0 1 3610
box -6 -8 126 248
use OAI21X1  _7619_
timestamp 0
transform -1 0 12190 0 1 2170
box -6 -8 106 248
use NOR2X1  _7620_
timestamp 0
transform 1 0 12250 0 1 2650
box -6 -8 86 248
use AOI21X1  _7621_
timestamp 0
transform 1 0 12370 0 1 2650
box -6 -8 106 248
use INVX1  _7622_
timestamp 0
transform 1 0 11930 0 -1 2170
box -6 -8 66 248
use NAND3X1  _7623_
timestamp 0
transform -1 0 9850 0 1 730
box -6 -8 106 248
use INVX1  _7624_
timestamp 0
transform 1 0 8910 0 -1 250
box -6 -8 66 248
use OAI21X1  _7625_
timestamp 0
transform 1 0 9350 0 1 250
box -6 -8 106 248
use INVX1  _7626_
timestamp 0
transform -1 0 10690 0 -1 1690
box -6 -8 66 248
use NAND3X1  _7627_
timestamp 0
transform 1 0 10350 0 -1 1690
box -6 -8 106 248
use OAI21X1  _7628_
timestamp 0
transform 1 0 10570 0 1 1210
box -6 -8 106 248
use NAND2X1  _7629_
timestamp 0
transform 1 0 11570 0 1 1690
box -6 -8 86 248
use AOI21X1  _7630_
timestamp 0
transform 1 0 11770 0 -1 2170
box -6 -8 106 248
use NAND3X1  _7631_
timestamp 0
transform 1 0 10190 0 -1 1690
box -6 -8 106 248
use NAND2X1  _7632_
timestamp 0
transform 1 0 10750 0 -1 1690
box -6 -8 86 248
use AOI21X1  _7633_
timestamp 0
transform 1 0 11270 0 1 1690
box -6 -8 106 248
use OAI21X1  _7634_
timestamp 0
transform 1 0 11950 0 1 2650
box -6 -8 106 248
use INVX1  _7635_
timestamp 0
transform -1 0 10750 0 1 3130
box -6 -8 66 248
use OR2X2  _7636_
timestamp 0
transform -1 0 11890 0 1 2650
box -6 -8 106 248
use OAI21X1  _7637_
timestamp 0
transform -1 0 11450 0 -1 3130
box -6 -8 106 248
use OAI22X1  _7638_
timestamp 0
transform 1 0 10590 0 -1 3610
box -6 -8 126 248
use NAND2X1  _7639_
timestamp 0
transform -1 0 10370 0 1 3130
box -6 -8 86 248
use NOR2X1  _7640_
timestamp 0
transform 1 0 11630 0 -1 3130
box -6 -8 86 248
use NOR2X1  _7641_
timestamp 0
transform 1 0 11510 0 -1 3130
box -6 -8 86 248
use OAI21X1  _7642_
timestamp 0
transform 1 0 9190 0 -1 730
box -6 -8 106 248
use INVX1  _7643_
timestamp 0
transform 1 0 10070 0 1 1210
box -6 -8 66 248
use OAI21X1  _7644_
timestamp 0
transform -1 0 10150 0 -1 1690
box -6 -8 106 248
use NAND2X1  _7645_
timestamp 0
transform -1 0 10950 0 1 1690
box -6 -8 86 248
use OR2X2  _7646_
timestamp 0
transform 1 0 11010 0 1 1690
box -6 -8 106 248
use NAND3X1  _7647_
timestamp 0
transform 1 0 11070 0 -1 2650
box -6 -8 106 248
use NAND2X1  _7648_
timestamp 0
transform 1 0 12870 0 1 2170
box -6 -8 86 248
use NAND2X1  _7649_
timestamp 0
transform -1 0 12810 0 1 2170
box -6 -8 86 248
use NAND2X1  _7650_
timestamp 0
transform 1 0 11210 0 -1 2650
box -6 -8 86 248
use AND2X2  _7651_
timestamp 0
transform -1 0 11150 0 -1 3130
box -6 -8 106 248
use OAI21X1  _7652_
timestamp 0
transform 1 0 11190 0 -1 3130
box -6 -8 106 248
use OAI21X1  _7653_
timestamp 0
transform -1 0 10530 0 1 3130
box -6 -8 106 248
use INVX1  _7654_
timestamp 0
transform 1 0 10150 0 1 3610
box -6 -8 66 248
use INVX1  _7655_
timestamp 0
transform 1 0 11530 0 1 2650
box -6 -8 66 248
use AOI21X1  _7656_
timestamp 0
transform -1 0 11750 0 1 2650
box -6 -8 106 248
use NOR2X1  _7657_
timestamp 0
transform 1 0 11490 0 -1 2650
box -6 -8 86 248
use NAND3X1  _7658_
timestamp 0
transform 1 0 11350 0 -1 2650
box -6 -8 106 248
use OAI21X1  _7659_
timestamp 0
transform 1 0 11390 0 1 2650
box -6 -8 106 248
use OAI21X1  _7660_
timestamp 0
transform 1 0 9490 0 -1 730
box -6 -8 106 248
use INVX1  _7661_
timestamp 0
transform -1 0 9490 0 1 730
box -6 -8 66 248
use OR2X2  _7662_
timestamp 0
transform -1 0 9610 0 -1 1210
box -6 -8 106 248
use OAI21X1  _7663_
timestamp 0
transform 1 0 9690 0 1 1210
box -6 -8 106 248
use NAND2X1  _7664_
timestamp 0
transform -1 0 10390 0 1 1690
box -6 -8 86 248
use OR2X2  _7665_
timestamp 0
transform 1 0 10450 0 1 1690
box -6 -8 106 248
use NAND3X1  _7666_
timestamp 0
transform 1 0 10590 0 1 1690
box -6 -8 106 248
use AND2X2  _7667_
timestamp 0
transform -1 0 9730 0 -1 1690
box -6 -8 106 248
use NOR2X1  _7668_
timestamp 0
transform 1 0 9910 0 -1 1690
box -6 -8 86 248
use OAI21X1  _7669_
timestamp 0
transform -1 0 9870 0 -1 1690
box -6 -8 106 248
use NAND2X1  _7670_
timestamp 0
transform 1 0 10810 0 -1 2650
box -6 -8 86 248
use AND2X2  _7671_
timestamp 0
transform -1 0 10850 0 -1 3130
box -6 -8 106 248
use NOR2X1  _7672_
timestamp 0
transform 1 0 10910 0 -1 3130
box -6 -8 86 248
use NOR2X1  _7673_
timestamp 0
transform -1 0 10650 0 1 3130
box -6 -8 86 248
use AOI22X1  _7674_
timestamp 0
transform 1 0 10190 0 -1 3610
box -6 -8 126 248
use NAND2X1  _7675_
timestamp 0
transform 1 0 9990 0 1 3130
box -6 -8 86 248
use INVX1  _7676_
timestamp 0
transform 1 0 11290 0 1 2650
box -6 -8 66 248
use AOI21X1  _7677_
timestamp 0
transform 1 0 11150 0 1 2650
box -6 -8 106 248
use NAND2X1  _7678_
timestamp 0
transform 1 0 10410 0 -1 2650
box -6 -8 86 248
use NOR2X1  _7679_
timestamp 0
transform 1 0 10290 0 -1 2650
box -6 -8 86 248
use AOI21X1  _7680_
timestamp 0
transform 1 0 10530 0 -1 2650
box -6 -8 106 248
use NOR2X1  _7681_
timestamp 0
transform 1 0 10670 0 -1 2650
box -6 -8 86 248
use AND2X2  _7682_
timestamp 0
transform -1 0 10710 0 -1 3130
box -6 -8 106 248
use OAI21X1  _7683_
timestamp 0
transform -1 0 10550 0 -1 3130
box -6 -8 106 248
use OAI21X1  _7684_
timestamp 0
transform -1 0 10230 0 1 3130
box -6 -8 106 248
use OAI21X1  _7685_
timestamp 0
transform 1 0 6850 0 -1 4570
box -6 -8 106 248
use OAI21X1  _7686_
timestamp 0
transform 1 0 6230 0 -1 5530
box -6 -8 106 248
use INVX1  _7687_
timestamp 0
transform -1 0 6350 0 1 5050
box -6 -8 66 248
use NOR2X1  _7688_
timestamp 0
transform -1 0 6190 0 -1 5050
box -6 -8 86 248
use NAND2X1  _7689_
timestamp 0
transform -1 0 6230 0 1 5050
box -6 -8 86 248
use NAND2X1  _7690_
timestamp 0
transform 1 0 5950 0 -1 5530
box -6 -8 86 248
use NAND2X1  _7691_
timestamp 0
transform -1 0 5810 0 1 5050
box -6 -8 86 248
use OAI21X1  _7692_
timestamp 0
transform -1 0 5910 0 -1 5530
box -6 -8 106 248
use NAND2X1  _7693_
timestamp 0
transform 1 0 5170 0 1 6010
box -6 -8 86 248
use INVX1  _7694_
timestamp 0
transform -1 0 5570 0 -1 6010
box -6 -8 66 248
use NOR2X1  _7695_
timestamp 0
transform 1 0 5090 0 1 5530
box -6 -8 86 248
use AOI21X1  _7696_
timestamp 0
transform -1 0 6190 0 -1 5530
box -6 -8 106 248
use NOR2X1  _7697_
timestamp 0
transform -1 0 6450 0 1 5530
box -6 -8 86 248
use OAI21X1  _7698_
timestamp 0
transform -1 0 6490 0 -1 5530
box -6 -8 106 248
use AND2X2  _7699_
timestamp 0
transform -1 0 6330 0 1 5530
box -6 -8 106 248
use OR2X2  _7700_
timestamp 0
transform -1 0 6010 0 -1 6010
box -6 -8 106 248
use OR2X2  _7701_
timestamp 0
transform -1 0 5930 0 1 6010
box -6 -8 106 248
use OAI21X1  _7702_
timestamp 0
transform -1 0 5870 0 -1 6010
box -6 -8 106 248
use NAND2X1  _7703_
timestamp 0
transform -1 0 5770 0 1 6010
box -6 -8 86 248
use NOR2X1  _7704_
timestamp 0
transform -1 0 5510 0 1 6010
box -6 -8 86 248
use NAND2X1  _7705_
timestamp 0
transform 1 0 5550 0 1 6010
box -6 -8 86 248
use NAND2X1  _7706_
timestamp 0
transform -1 0 5390 0 1 6010
box -6 -8 86 248
use OAI21X1  _7707_
timestamp 0
transform -1 0 5130 0 1 6010
box -6 -8 106 248
use INVX1  _7708_
timestamp 0
transform -1 0 6130 0 -1 6010
box -6 -8 66 248
use OAI21X1  _7709_
timestamp 0
transform -1 0 6070 0 1 6010
box -6 -8 106 248
use OAI21X1  _7710_
timestamp 0
transform 1 0 7250 0 1 4090
box -6 -8 106 248
use OAI21X1  _7711_
timestamp 0
transform 1 0 7450 0 1 6010
box -6 -8 106 248
use MUX2X1  _7712_
timestamp 0
transform 1 0 7290 0 1 6010
box -6 -8 126 248
use NAND2X1  _7713_
timestamp 0
transform 1 0 7650 0 -1 6490
box -6 -8 86 248
use OR2X2  _7714_
timestamp 0
transform -1 0 7590 0 -1 6490
box -6 -8 106 248
use NAND2X1  _7715_
timestamp 0
transform 1 0 7370 0 -1 6490
box -6 -8 86 248
use INVX1  _7716_
timestamp 0
transform -1 0 6890 0 1 6490
box -6 -8 66 248
use NOR2X1  _7717_
timestamp 0
transform -1 0 6550 0 1 6490
box -6 -8 86 248
use NAND2X1  _7718_
timestamp 0
transform -1 0 6890 0 -1 6490
box -6 -8 86 248
use NAND2X1  _7719_
timestamp 0
transform 1 0 6570 0 -1 6490
box -6 -8 86 248
use OAI22X1  _7720_
timestamp 0
transform 1 0 6310 0 1 6490
box -6 -8 126 248
use NOR2X1  _7721_
timestamp 0
transform -1 0 5870 0 -1 6490
box -6 -8 86 248
use NAND2X1  _7722_
timestamp 0
transform -1 0 7030 0 -1 6490
box -6 -8 86 248
use INVX1  _7723_
timestamp 0
transform -1 0 6750 0 -1 6490
box -6 -8 66 248
use INVX1  _7724_
timestamp 0
transform -1 0 6750 0 -1 5050
box -6 -8 66 248
use NOR2X1  _7725_
timestamp 0
transform -1 0 7790 0 1 3610
box -6 -8 86 248
use OAI21X1  _7726_
timestamp 0
transform -1 0 7650 0 1 3610
box -6 -8 106 248
use OAI21X1  _7727_
timestamp 0
transform 1 0 7090 0 1 4090
box -6 -8 106 248
use OAI21X1  _7728_
timestamp 0
transform 1 0 7390 0 1 4090
box -6 -8 106 248
use NOR2X1  _7729_
timestamp 0
transform -1 0 6630 0 -1 5530
box -6 -8 86 248
use NAND2X1  _7730_
timestamp 0
transform 1 0 6670 0 -1 5530
box -6 -8 86 248
use INVX1  _7731_
timestamp 0
transform -1 0 6390 0 -1 6010
box -6 -8 66 248
use NOR2X1  _7732_
timestamp 0
transform -1 0 6450 0 1 6010
box -6 -8 86 248
use OAI21X1  _7733_
timestamp 0
transform 1 0 6430 0 -1 6490
box -6 -8 106 248
use AOI21X1  _7734_
timestamp 0
transform -1 0 6390 0 -1 6490
box -6 -8 106 248
use NOR2X1  _7735_
timestamp 0
transform 1 0 6150 0 -1 6490
box -6 -8 86 248
use NAND2X1  _7736_
timestamp 0
transform -1 0 6570 0 1 6010
box -6 -8 86 248
use INVX1  _7737_
timestamp 0
transform -1 0 8170 0 -1 6010
box -6 -8 66 248
use AOI21X1  _7738_
timestamp 0
transform -1 0 7450 0 1 5050
box -6 -8 106 248
use OAI21X1  _7739_
timestamp 0
transform 1 0 7210 0 1 5050
box -6 -8 106 248
use OAI21X1  _7740_
timestamp 0
transform 1 0 6790 0 -1 5530
box -6 -8 106 248
use OR2X2  _7741_
timestamp 0
transform 1 0 7730 0 -1 5530
box -6 -8 106 248
use NAND2X1  _7742_
timestamp 0
transform -1 0 7550 0 -1 5530
box -6 -8 86 248
use NAND2X1  _7743_
timestamp 0
transform 1 0 7590 0 -1 5530
box -6 -8 86 248
use AOI21X1  _7744_
timestamp 0
transform -1 0 6670 0 -1 6010
box -6 -8 106 248
use AND2X2  _7745_
timestamp 0
transform -1 0 7090 0 1 6010
box -6 -8 106 248
use OAI21X1  _7746_
timestamp 0
transform 1 0 7150 0 1 6010
box -6 -8 106 248
use OAI21X1  _7747_
timestamp 0
transform -1 0 6950 0 1 6010
box -6 -8 106 248
use OAI21X1  _7748_
timestamp 0
transform 1 0 7610 0 1 5530
box -6 -8 106 248
use INVX1  _7749_
timestamp 0
transform -1 0 8210 0 -1 5530
box -6 -8 66 248
use OAI21X1  _7750_
timestamp 0
transform 1 0 8190 0 -1 3610
box -6 -8 106 248
use OAI21X1  _7751_
timestamp 0
transform 1 0 8870 0 -1 4570
box -6 -8 106 248
use OR2X2  _7752_
timestamp 0
transform -1 0 8810 0 -1 4570
box -6 -8 106 248
use NAND2X1  _7753_
timestamp 0
transform 1 0 8310 0 1 4090
box -6 -8 86 248
use OR2X2  _7754_
timestamp 0
transform -1 0 8250 0 1 5530
box -6 -8 106 248
use NAND2X1  _7755_
timestamp 0
transform 1 0 8290 0 1 5530
box -6 -8 86 248
use NAND2X1  _7756_
timestamp 0
transform -1 0 8110 0 1 5530
box -6 -8 86 248
use INVX1  _7757_
timestamp 0
transform -1 0 7810 0 1 5530
box -6 -8 66 248
use NOR2X1  _7758_
timestamp 0
transform 1 0 7490 0 1 5530
box -6 -8 86 248
use NAND2X1  _7759_
timestamp 0
transform 1 0 7350 0 1 5530
box -6 -8 86 248
use NAND2X1  _7760_
timestamp 0
transform 1 0 7190 0 -1 5530
box -6 -8 86 248
use OAI22X1  _7761_
timestamp 0
transform 1 0 7310 0 -1 5530
box -6 -8 126 248
use NAND2X1  _7762_
timestamp 0
transform -1 0 6510 0 -1 6010
box -6 -8 86 248
use INVX1  _7763_
timestamp 0
transform -1 0 7570 0 -1 6010
box -6 -8 66 248
use NAND2X1  _7764_
timestamp 0
transform -1 0 7690 0 -1 6010
box -6 -8 86 248
use OAI21X1  _7765_
timestamp 0
transform 1 0 7870 0 1 5530
box -6 -8 106 248
use INVX1  _7766_
timestamp 0
transform 1 0 7870 0 -1 6010
box -6 -8 66 248
use OAI21X1  _7767_
timestamp 0
transform 1 0 7730 0 -1 6010
box -6 -8 106 248
use OAI21X1  _7768_
timestamp 0
transform 1 0 7910 0 -1 3610
box -6 -8 106 248
use NOR2X1  _7769_
timestamp 0
transform 1 0 7970 0 1 3610
box -6 -8 86 248
use NAND2X1  _7770_
timestamp 0
transform 1 0 7870 0 -1 4090
box -6 -8 86 248
use OAI21X1  _7771_
timestamp 0
transform -1 0 7930 0 1 3610
box -6 -8 106 248
use NAND2X1  _7772_
timestamp 0
transform -1 0 7810 0 -1 4090
box -6 -8 86 248
use NAND2X1  _7773_
timestamp 0
transform 1 0 7630 0 1 5050
box -6 -8 86 248
use OR2X2  _7774_
timestamp 0
transform -1 0 7590 0 1 5050
box -6 -8 106 248
use NAND2X1  _7775_
timestamp 0
transform 1 0 6950 0 -1 5530
box -6 -8 86 248
use INVX1  _7776_
timestamp 0
transform 1 0 7070 0 -1 5530
box -6 -8 66 248
use NOR2X1  _7777_
timestamp 0
transform 1 0 7370 0 -1 6010
box -6 -8 86 248
use NAND2X1  _7778_
timestamp 0
transform -1 0 7310 0 -1 6010
box -6 -8 86 248
use NAND2X1  _7779_
timestamp 0
transform 1 0 7110 0 -1 6010
box -6 -8 86 248
use OAI21X1  _7780_
timestamp 0
transform -1 0 7050 0 -1 6010
box -6 -8 106 248
use INVX1  _7781_
timestamp 0
transform 1 0 5550 0 1 5530
box -6 -8 66 248
use NAND2X1  _7782_
timestamp 0
transform 1 0 6670 0 1 5530
box -6 -8 86 248
use INVX1  _7783_
timestamp 0
transform 1 0 5150 0 1 5050
box -6 -8 66 248
use NAND2X1  _7784_
timestamp 0
transform -1 0 4990 0 -1 5530
box -6 -8 86 248
use OR2X2  _7785_
timestamp 0
transform -1 0 4850 0 -1 5530
box -6 -8 106 248
use NAND2X1  _7786_
timestamp 0
transform 1 0 5030 0 -1 5530
box -6 -8 86 248
use NOR2X1  _7787_
timestamp 0
transform -1 0 5250 0 -1 5530
box -6 -8 86 248
use INVX1  _7788_
timestamp 0
transform 1 0 5210 0 1 5530
box -6 -8 66 248
use NAND2X1  _7789_
timestamp 0
transform 1 0 5310 0 -1 5530
box -6 -8 86 248
use NAND2X1  _7790_
timestamp 0
transform 1 0 5650 0 1 5530
box -6 -8 86 248
use OR2X2  _7791_
timestamp 0
transform -1 0 6190 0 1 5530
box -6 -8 106 248
use AOI21X1  _7792_
timestamp 0
transform -1 0 6030 0 1 5530
box -6 -8 106 248
use AOI22X1  _7793_
timestamp 0
transform 1 0 5770 0 1 5530
box -6 -8 126 248
use NAND2X1  _7794_
timestamp 0
transform -1 0 8570 0 -1 5050
box -6 -8 86 248
use NOR2X1  _7795_
timestamp 0
transform -1 0 7070 0 -1 4570
box -6 -8 86 248
use INVX1  _7796_
timestamp 0
transform 1 0 7130 0 -1 4570
box -6 -8 66 248
use NAND3X1  _7797_
timestamp 0
transform 1 0 7390 0 -1 4570
box -6 -8 106 248
use INVX1  _7798_
timestamp 0
transform -1 0 7390 0 -1 5050
box -6 -8 66 248
use AOI21X1  _7799_
timestamp 0
transform -1 0 7350 0 -1 4570
box -6 -8 106 248
use NOR2X1  _7800_
timestamp 0
transform -1 0 7290 0 -1 5050
box -6 -8 86 248
use OAI21X1  _7801_
timestamp 0
transform -1 0 6610 0 1 5530
box -6 -8 106 248
use NOR2X1  _7802_
timestamp 0
transform 1 0 6790 0 1 5530
box -6 -8 86 248
use AOI21X1  _7803_
timestamp 0
transform -1 0 7030 0 1 5530
box -6 -8 106 248
use NAND3X1  _7804_
timestamp 0
transform -1 0 7310 0 1 5530
box -6 -8 106 248
use OAI21X1  _7805_
timestamp 0
transform -1 0 7170 0 1 5530
box -6 -8 106 248
use NOR2X1  _7806_
timestamp 0
transform -1 0 7530 0 -1 5050
box -6 -8 86 248
use NAND2X1  _7807_
timestamp 0
transform -1 0 7830 0 1 5050
box -6 -8 86 248
use NAND2X1  _7808_
timestamp 0
transform 1 0 8230 0 1 5050
box -6 -8 86 248
use OAI21X1  _7809_
timestamp 0
transform 1 0 8470 0 1 5050
box -6 -8 106 248
use AOI21X1  _7810_
timestamp 0
transform -1 0 7170 0 -1 5050
box -6 -8 106 248
use OR2X2  _7811_
timestamp 0
transform -1 0 8130 0 1 4570
box -6 -8 106 248
use NAND2X1  _7812_
timestamp 0
transform 1 0 8170 0 1 4570
box -6 -8 86 248
use NAND2X1  _7813_
timestamp 0
transform 1 0 7910 0 1 4570
box -6 -8 86 248
use AND2X2  _7814_
timestamp 0
transform -1 0 6650 0 -1 5050
box -6 -8 106 248
use OAI21X1  _7815_
timestamp 0
transform -1 0 6510 0 -1 5050
box -6 -8 106 248
use OAI22X1  _7816_
timestamp 0
transform 1 0 6230 0 -1 5050
box -6 -8 126 248
use NAND2X1  _7817_
timestamp 0
transform 1 0 5950 0 1 4570
box -6 -8 86 248
use OAI21X1  _7818_
timestamp 0
transform 1 0 7490 0 1 4570
box -6 -8 106 248
use NAND3X1  _7819_
timestamp 0
transform -1 0 7850 0 1 4570
box -6 -8 106 248
use INVX1  _7820_
timestamp 0
transform 1 0 7650 0 1 4570
box -6 -8 66 248
use AOI21X1  _7821_
timestamp 0
transform -1 0 7430 0 1 4570
box -6 -8 106 248
use INVX1  _7822_
timestamp 0
transform 1 0 7090 0 -1 4090
box -6 -8 66 248
use NAND2X1  _7823_
timestamp 0
transform 1 0 6950 0 -1 4090
box -6 -8 86 248
use NAND2X1  _7824_
timestamp 0
transform -1 0 6550 0 -1 4570
box -6 -8 86 248
use NAND2X1  _7825_
timestamp 0
transform -1 0 6430 0 -1 4570
box -6 -8 86 248
use AND2X2  _7826_
timestamp 0
transform -1 0 6130 0 -1 4570
box -6 -8 106 248
use OAI21X1  _7827_
timestamp 0
transform 1 0 6190 0 -1 4570
box -6 -8 106 248
use OAI21X1  _7828_
timestamp 0
transform -1 0 5990 0 -1 4570
box -6 -8 106 248
use NAND2X1  _7829_
timestamp 0
transform 1 0 6070 0 1 4570
box -6 -8 86 248
use OAI21X1  _7830_
timestamp 0
transform 1 0 6350 0 1 4570
box -6 -8 106 248
use OAI21X1  _7831_
timestamp 0
transform -1 0 6290 0 1 4570
box -6 -8 106 248
use NAND2X1  _7832_
timestamp 0
transform 1 0 6790 0 1 3610
box -6 -8 86 248
use NAND2X1  _7833_
timestamp 0
transform 1 0 8390 0 -1 4090
box -6 -8 86 248
use NOR2X1  _7834_
timestamp 0
transform 1 0 6930 0 1 3610
box -6 -8 86 248
use NAND2X1  _7835_
timestamp 0
transform -1 0 8710 0 1 1210
box -6 -8 86 248
use OAI21X1  _7836_
timestamp 0
transform -1 0 8850 0 1 1210
box -6 -8 106 248
use NAND2X1  _7837_
timestamp 0
transform 1 0 6930 0 -1 250
box -6 -8 86 248
use OAI21X1  _7838_
timestamp 0
transform -1 0 7030 0 1 250
box -6 -8 106 248
use INVX1  _7839_
timestamp 0
transform -1 0 10590 0 1 2650
box -6 -8 66 248
use OR2X2  _7840_
timestamp 0
transform -1 0 7630 0 1 4090
box -6 -8 106 248
use OAI21X1  _7841_
timestamp 0
transform 1 0 9630 0 -1 3130
box -6 -8 106 248
use OAI21X1  _7842_
timestamp 0
transform -1 0 10010 0 -1 3130
box -6 -8 106 248
use INVX1  _7843_
timestamp 0
transform -1 0 8870 0 -1 3610
box -6 -8 66 248
use OAI21X1  _7844_
timestamp 0
transform 1 0 9310 0 -1 3610
box -6 -8 106 248
use OAI21X1  _7845_
timestamp 0
transform 1 0 9150 0 -1 3610
box -6 -8 106 248
use NAND2X1  _7846_
timestamp 0
transform -1 0 6750 0 1 4570
box -6 -8 86 248
use NAND2X1  _7847_
timestamp 0
transform -1 0 10710 0 1 2650
box -6 -8 86 248
use OAI21X1  _7848_
timestamp 0
transform 1 0 10750 0 1 2650
box -6 -8 106 248
use NAND2X1  _7849_
timestamp 0
transform 1 0 9790 0 -1 3130
box -6 -8 86 248
use OAI21X1  _7850_
timestamp 0
transform 1 0 9590 0 1 3130
box -6 -8 106 248
use AND2X2  _7851_
timestamp 0
transform -1 0 6270 0 1 4090
box -6 -8 106 248
use NAND2X1  _7852_
timestamp 0
transform 1 0 11150 0 -1 2170
box -6 -8 86 248
use OAI21X1  _7853_
timestamp 0
transform 1 0 11010 0 -1 2170
box -6 -8 106 248
use NAND2X1  _7854_
timestamp 0
transform 1 0 8930 0 -1 1690
box -6 -8 86 248
use OAI21X1  _7855_
timestamp 0
transform -1 0 8890 0 -1 1690
box -6 -8 106 248
use OAI21X1  _7856_
timestamp 0
transform 1 0 8950 0 1 3130
box -6 -8 106 248
use OAI21X1  _7857_
timestamp 0
transform -1 0 9190 0 1 3130
box -6 -8 106 248
use OAI21X1  _7858_
timestamp 0
transform -1 0 8890 0 1 3130
box -6 -8 106 248
use OAI21X1  _7859_
timestamp 0
transform -1 0 8730 0 1 3130
box -6 -8 106 248
use NAND2X1  _7860_
timestamp 0
transform -1 0 9070 0 -1 3130
box -6 -8 86 248
use OAI21X1  _7861_
timestamp 0
transform -1 0 9230 0 -1 3130
box -6 -8 106 248
use NAND2X1  _7862_
timestamp 0
transform 1 0 10250 0 1 2650
box -6 -8 86 248
use OAI21X1  _7863_
timestamp 0
transform 1 0 10110 0 1 2650
box -6 -8 106 248
use NAND2X1  _7864_
timestamp 0
transform -1 0 7310 0 -1 730
box -6 -8 86 248
use OAI21X1  _7865_
timestamp 0
transform -1 0 7190 0 -1 730
box -6 -8 106 248
use NAND2X1  _7866_
timestamp 0
transform 1 0 7290 0 -1 250
box -6 -8 86 248
use OAI21X1  _7867_
timestamp 0
transform 1 0 7150 0 -1 250
box -6 -8 106 248
use INVX1  _7868_
timestamp 0
transform -1 0 6870 0 1 3130
box -6 -8 66 248
use OAI21X1  _7869_
timestamp 0
transform -1 0 7010 0 1 3130
box -6 -8 106 248
use OAI21X1  _7870_
timestamp 0
transform -1 0 7170 0 1 3130
box -6 -8 106 248
use INVX1  _7871_
timestamp 0
transform -1 0 7030 0 -1 3130
box -6 -8 66 248
use OAI21X1  _7872_
timestamp 0
transform -1 0 8050 0 -1 3130
box -6 -8 106 248
use OAI21X1  _7873_
timestamp 0
transform 1 0 7550 0 -1 3130
box -6 -8 106 248
use NAND2X1  _7874_
timestamp 0
transform 1 0 6510 0 1 3130
box -6 -8 86 248
use OAI21X1  _7875_
timestamp 0
transform -1 0 6750 0 1 3130
box -6 -8 106 248
use NAND2X1  _7876_
timestamp 0
transform 1 0 6690 0 -1 3130
box -6 -8 86 248
use OAI21X1  _7877_
timestamp 0
transform -1 0 6930 0 -1 3130
box -6 -8 106 248
use NAND2X1  _7878_
timestamp 0
transform -1 0 6350 0 -1 250
box -6 -8 86 248
use OAI21X1  _7879_
timestamp 0
transform 1 0 6130 0 -1 250
box -6 -8 106 248
use NAND2X1  _7880_
timestamp 0
transform -1 0 6170 0 1 250
box -6 -8 86 248
use OAI21X1  _7881_
timestamp 0
transform -1 0 6310 0 1 250
box -6 -8 106 248
use OAI21X1  _7882_
timestamp 0
transform -1 0 7290 0 -1 3610
box -6 -8 106 248
use OAI21X1  _7883_
timestamp 0
transform 1 0 7030 0 -1 3610
box -6 -8 106 248
use OAI21X1  _7884_
timestamp 0
transform -1 0 7330 0 1 3130
box -6 -8 106 248
use OAI21X1  _7885_
timestamp 0
transform -1 0 7470 0 1 3130
box -6 -8 106 248
use NAND2X1  _7886_
timestamp 0
transform -1 0 8170 0 -1 3130
box -6 -8 86 248
use OAI21X1  _7887_
timestamp 0
transform 1 0 8230 0 -1 3130
box -6 -8 106 248
use NAND2X1  _7888_
timestamp 0
transform -1 0 7410 0 -1 3610
box -6 -8 86 248
use OAI21X1  _7889_
timestamp 0
transform -1 0 7570 0 -1 3610
box -6 -8 106 248
use NAND2X1  _7890_
timestamp 0
transform 1 0 7350 0 -1 4090
box -6 -8 86 248
use OAI21X1  _7891_
timestamp 0
transform 1 0 7210 0 -1 4090
box -6 -8 106 248
use NAND2X1  _7892_
timestamp 0
transform 1 0 8510 0 1 3130
box -6 -8 86 248
use OAI21X1  _7893_
timestamp 0
transform 1 0 8370 0 1 3130
box -6 -8 106 248
use INVX1  _7894_
timestamp 0
transform 1 0 8370 0 1 5050
box -6 -8 66 248
use OAI21X1  _7895_
timestamp 0
transform 1 0 8070 0 -1 4570
box -6 -8 106 248
use OAI21X1  _7896_
timestamp 0
transform -1 0 8330 0 -1 4570
box -6 -8 106 248
use INVX1  _7897_
timestamp 0
transform -1 0 7010 0 -1 5050
box -6 -8 66 248
use OAI21X1  _7898_
timestamp 0
transform 1 0 7930 0 -1 4570
box -6 -8 106 248
use OAI21X1  _7899_
timestamp 0
transform 1 0 7550 0 -1 4570
box -6 -8 106 248
use NAND2X1  _7900_
timestamp 0
transform -1 0 8030 0 -1 5050
box -6 -8 86 248
use OAI21X1  _7901_
timestamp 0
transform -1 0 8190 0 -1 5050
box -6 -8 106 248
use NAND2X1  _7902_
timestamp 0
transform 1 0 5070 0 -1 5050
box -6 -8 86 248
use OAI21X1  _7903_
timestamp 0
transform -1 0 5030 0 -1 5050
box -6 -8 106 248
use NAND2X1  _7904_
timestamp 0
transform -1 0 7950 0 -1 5530
box -6 -8 86 248
use OAI21X1  _7905_
timestamp 0
transform -1 0 8090 0 -1 5530
box -6 -8 106 248
use NAND2X1  _7906_
timestamp 0
transform 1 0 8870 0 1 5050
box -6 -8 86 248
use OAI21X1  _7907_
timestamp 0
transform 1 0 8490 0 -1 5530
box -6 -8 106 248
use OAI21X1  _7908_
timestamp 0
transform -1 0 8410 0 1 4570
box -6 -8 106 248
use OAI21X1  _7909_
timestamp 0
transform -1 0 7910 0 -1 5050
box -6 -8 106 248
use OAI21X1  _7910_
timestamp 0
transform 1 0 6790 0 1 4570
box -6 -8 106 248
use OAI21X1  _7911_
timestamp 0
transform -1 0 7050 0 1 4570
box -6 -8 106 248
use NAND2X1  _7912_
timestamp 0
transform 1 0 7070 0 1 5050
box -6 -8 86 248
use OAI21X1  _7913_
timestamp 0
transform 1 0 6810 0 1 5050
box -6 -8 106 248
use NAND2X1  _7914_
timestamp 0
transform 1 0 6950 0 1 5050
box -6 -8 86 248
use OAI21X1  _7915_
timestamp 0
transform 1 0 6190 0 -1 6010
box -6 -8 106 248
use DFFPOSX1  _7916_
timestamp 0
transform -1 0 7030 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _7917_
timestamp 0
transform -1 0 6790 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _7918_
timestamp 0
transform -1 0 8070 0 -1 6490
box -6 -8 246 248
use DFFPOSX1  _7919_
timestamp 0
transform 1 0 6070 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _7920_
timestamp 0
transform -1 0 6230 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _7921_
timestamp 0
transform 1 0 5370 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _7922_
timestamp 0
transform 1 0 5690 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _7923_
timestamp 0
transform 1 0 5170 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _7924_
timestamp 0
transform 1 0 4470 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _7925_
timestamp 0
transform 1 0 5710 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _7926_
timestamp 0
transform 1 0 5070 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _7927_
timestamp 0
transform 1 0 5530 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _7928_
timestamp 0
transform 1 0 4710 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _7929_
timestamp 0
transform -1 0 8570 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _7930_
timestamp 0
transform 1 0 8390 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _7931_
timestamp 0
transform -1 0 9210 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _7932_
timestamp 0
transform -1 0 9750 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _7933_
timestamp 0
transform -1 0 11110 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _7934_
timestamp 0
transform -1 0 10010 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _7935_
timestamp 0
transform -1 0 9370 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _7936_
timestamp 0
transform -1 0 10490 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _7937_
timestamp 0
transform -1 0 10670 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _7938_
timestamp 0
transform -1 0 10550 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _7939_
timestamp 0
transform -1 0 10110 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _7940_
timestamp 0
transform -1 0 10150 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _7941_
timestamp 0
transform 1 0 5530 0 -1 5530
box -6 -8 246 248
use DFFPOSX1  _7942_
timestamp 0
transform 1 0 4930 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _7943_
timestamp 0
transform 1 0 5890 0 1 6490
box -6 -8 246 248
use DFFPOSX1  _7944_
timestamp 0
transform -1 0 6110 0 -1 6490
box -6 -8 246 248
use DFFPOSX1  _7945_
timestamp 0
transform -1 0 6810 0 1 6010
box -6 -8 246 248
use DFFPOSX1  _7946_
timestamp 0
transform -1 0 8170 0 1 5050
box -6 -8 246 248
use DFFPOSX1  _7947_
timestamp 0
transform -1 0 6910 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _7948_
timestamp 0
transform 1 0 5270 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _7949_
timestamp 0
transform -1 0 8810 0 1 5050
box -6 -8 246 248
use DFFPOSX1  _7950_
timestamp 0
transform -1 0 5790 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _7951_
timestamp 0
transform 1 0 5610 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _7952_
timestamp 0
transform -1 0 5910 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _7953_
timestamp 0
transform 1 0 8850 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _7954_
timestamp 0
transform 1 0 7030 0 1 250
box -6 -8 246 248
use DFFPOSX1  _7955_
timestamp 0
transform -1 0 10410 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _7956_
timestamp 0
transform 1 0 8870 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _7957_
timestamp 0
transform 1 0 10850 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _7958_
timestamp 0
transform 1 0 9690 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _7959_
timestamp 0
transform -1 0 10810 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _7960_
timestamp 0
transform -1 0 8630 0 -1 1690
box -6 -8 246 248
use DFFPOSX1  _7961_
timestamp 0
transform 1 0 9190 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _7962_
timestamp 0
transform 1 0 8530 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _7963_
timestamp 0
transform -1 0 9570 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _7964_
timestamp 0
transform -1 0 10050 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _7965_
timestamp 0
transform 1 0 6650 0 1 250
box -6 -8 246 248
use DFFPOSX1  _7966_
timestamp 0
transform 1 0 6630 0 -1 250
box -6 -8 246 248
use DFFPOSX1  _7967_
timestamp 0
transform 1 0 7650 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _7968_
timestamp 0
transform -1 0 7510 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _7969_
timestamp 0
transform -1 0 6470 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _7970_
timestamp 0
transform -1 0 6650 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _7971_
timestamp 0
transform -1 0 6090 0 -1 250
box -6 -8 246 248
use DFFPOSX1  _7972_
timestamp 0
transform 1 0 6310 0 1 250
box -6 -8 246 248
use DFFPOSX1  _7973_
timestamp 0
transform 1 0 6750 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _7974_
timestamp 0
transform -1 0 7270 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _7975_
timestamp 0
transform 1 0 7590 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _7976_
timestamp 0
transform 1 0 7270 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _7977_
timestamp 0
transform 1 0 6410 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _7978_
timestamp 0
transform -1 0 8330 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _7979_
timestamp 0
transform -1 0 8570 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _7980_
timestamp 0
transform 1 0 7650 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _7981_
timestamp 0
transform -1 0 8430 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _7982_
timestamp 0
transform 1 0 4390 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _7983_
timestamp 0
transform -1 0 8410 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _7984_
timestamp 0
transform -1 0 8450 0 -1 5530
box -6 -8 246 248
use DFFPOSX1  _7985_
timestamp 0
transform -1 0 7770 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _7986_
timestamp 0
transform -1 0 7290 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _7987_
timestamp 0
transform -1 0 6750 0 1 5050
box -6 -8 246 248
use DFFPOSX1  _7988_
timestamp 0
transform -1 0 6310 0 1 6010
box -6 -8 246 248
use DFFPOSX1  _7989_
timestamp 0
transform -1 0 12190 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _7990_
timestamp 0
transform 1 0 8410 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _7991_
timestamp 0
transform 1 0 8890 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _7992_
timestamp 0
transform -1 0 5110 0 1 5050
box -6 -8 246 248
use DFFPOSX1  _7993_
timestamp 0
transform 1 0 4630 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _7994_
timestamp 0
transform 1 0 5490 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _7995_
timestamp 0
transform 1 0 5730 0 1 4090
box -6 -8 246 248
use INVX1  _7996_
timestamp 0
transform -1 0 6290 0 1 7930
box -6 -8 66 248
use INVX2  _7997_
timestamp 0
transform -1 0 5250 0 -1 7930
box -6 -8 66 248
use NOR2X1  _7998_
timestamp 0
transform -1 0 5030 0 -1 7930
box -6 -8 86 248
use INVX2  _7999_
timestamp 0
transform 1 0 5010 0 -1 8410
box -6 -8 66 248
use NOR2X1  _8000_
timestamp 0
transform 1 0 4370 0 -1 6970
box -6 -8 86 248
use INVX4  _8001_
timestamp 0
transform 1 0 4230 0 -1 7450
box -6 -8 86 248
use NOR2X1  _8002_
timestamp 0
transform -1 0 4590 0 1 6970
box -6 -8 86 248
use OAI21X1  _8003_
timestamp 0
transform -1 0 4750 0 1 7450
box -6 -8 106 248
use INVX2  _8004_
timestamp 0
transform -1 0 4570 0 -1 7450
box -6 -8 66 248
use AND2X2  _8005_
timestamp 0
transform -1 0 4470 0 -1 7450
box -6 -8 106 248
use AOI22X1  _8006_
timestamp 0
transform -1 0 5410 0 1 7930
box -6 -8 126 248
use OAI21X1  _8007_
timestamp 0
transform 1 0 4510 0 1 7450
box -6 -8 106 248
use NOR2X1  _8008_
timestamp 0
transform 1 0 5070 0 -1 7930
box -6 -8 86 248
use AOI22X1  _8009_
timestamp 0
transform 1 0 4330 0 1 7450
box -6 -8 126 248
use OAI21X1  _8010_
timestamp 0
transform -1 0 3890 0 1 7450
box -6 -8 106 248
use INVX1  _8011_
timestamp 0
transform -1 0 5510 0 -1 6490
box -6 -8 66 248
use OAI21X1  _8012_
timestamp 0
transform -1 0 4130 0 1 6490
box -6 -8 106 248
use AOI21X1  _8013_
timestamp 0
transform -1 0 4270 0 1 6490
box -6 -8 106 248
use INVX1  _8014_
timestamp 0
transform 1 0 6590 0 -1 7450
box -6 -8 66 248
use NAND2X1  _8015_
timestamp 0
transform -1 0 5110 0 -1 7450
box -6 -8 86 248
use OAI21X1  _8016_
timestamp 0
transform 1 0 4890 0 -1 7450
box -6 -8 106 248
use OAI21X1  _8017_
timestamp 0
transform 1 0 4890 0 1 6970
box -6 -8 106 248
use AOI22X1  _8018_
timestamp 0
transform -1 0 5010 0 1 7930
box -6 -8 126 248
use NAND2X1  _8019_
timestamp 0
transform -1 0 4590 0 -1 6970
box -6 -8 86 248
use INVX1  _8020_
timestamp 0
transform 1 0 3310 0 -1 7930
box -6 -8 66 248
use OAI21X1  _8021_
timestamp 0
transform 1 0 4390 0 -1 7930
box -6 -8 106 248
use AOI21X1  _8022_
timestamp 0
transform -1 0 4350 0 -1 7930
box -6 -8 106 248
use INVX1  _8023_
timestamp 0
transform 1 0 3350 0 1 8410
box -6 -8 66 248
use NAND2X1  _8024_
timestamp 0
transform 1 0 3010 0 1 7930
box -6 -8 86 248
use OAI21X1  _8025_
timestamp 0
transform -1 0 3510 0 1 7930
box -6 -8 106 248
use OAI21X1  _8026_
timestamp 0
transform -1 0 3670 0 1 7930
box -6 -8 106 248
use AOI22X1  _8027_
timestamp 0
transform -1 0 4350 0 -1 8890
box -6 -8 126 248
use NAND2X1  _8028_
timestamp 0
transform -1 0 3790 0 1 7930
box -6 -8 86 248
use INVX1  _8029_
timestamp 0
transform 1 0 3390 0 1 6970
box -6 -8 66 248
use OAI21X1  _8030_
timestamp 0
transform 1 0 3810 0 -1 7450
box -6 -8 106 248
use AOI21X1  _8031_
timestamp 0
transform -1 0 3770 0 -1 7450
box -6 -8 106 248
use INVX1  _8032_
timestamp 0
transform 1 0 2890 0 1 7930
box -6 -8 66 248
use NAND2X1  _8033_
timestamp 0
transform 1 0 3150 0 1 7930
box -6 -8 86 248
use OAI21X1  _8034_
timestamp 0
transform -1 0 3370 0 1 7930
box -6 -8 106 248
use OAI21X1  _8035_
timestamp 0
transform -1 0 3470 0 1 7450
box -6 -8 106 248
use AOI22X1  _8036_
timestamp 0
transform -1 0 4490 0 1 7930
box -6 -8 126 248
use NAND2X1  _8037_
timestamp 0
transform -1 0 3590 0 1 7450
box -6 -8 86 248
use INVX1  _8038_
timestamp 0
transform 1 0 3110 0 1 6970
box -6 -8 66 248
use OAI21X1  _8039_
timestamp 0
transform 1 0 4110 0 1 6970
box -6 -8 106 248
use AOI21X1  _8040_
timestamp 0
transform 1 0 3870 0 1 6970
box -6 -8 106 248
use INVX1  _8041_
timestamp 0
transform 1 0 4470 0 -1 8410
box -6 -8 66 248
use NAND2X1  _8042_
timestamp 0
transform 1 0 4690 0 -1 7930
box -6 -8 86 248
use OAI21X1  _8043_
timestamp 0
transform 1 0 4550 0 -1 7930
box -6 -8 106 248
use OAI21X1  _8044_
timestamp 0
transform -1 0 3830 0 1 6970
box -6 -8 106 248
use AOI22X1  _8045_
timestamp 0
transform 1 0 3950 0 -1 7930
box -6 -8 126 248
use NAND2X1  _8046_
timestamp 0
transform -1 0 3690 0 1 6970
box -6 -8 86 248
use INVX1  _8047_
timestamp 0
transform 1 0 2790 0 -1 7930
box -6 -8 66 248
use NOR2X1  _8048_
timestamp 0
transform -1 0 3650 0 -1 6970
box -6 -8 86 248
use OAI21X1  _8049_
timestamp 0
transform 1 0 3950 0 -1 7450
box -6 -8 106 248
use AOI22X1  _8050_
timestamp 0
transform 1 0 4590 0 -1 8410
box -6 -8 126 248
use OAI21X1  _8051_
timestamp 0
transform 1 0 3630 0 1 7450
box -6 -8 106 248
use AOI22X1  _8052_
timestamp 0
transform 1 0 3070 0 1 7450
box -6 -8 126 248
use OAI21X1  _8053_
timestamp 0
transform 1 0 2930 0 1 7450
box -6 -8 106 248
use INVX1  _8054_
timestamp 0
transform 1 0 4630 0 1 8890
box -6 -8 66 248
use INVX1  _8055_
timestamp 0
transform -1 0 5470 0 1 9850
box -6 -8 66 248
use INVX8  _8056_
timestamp 0
transform -1 0 1410 0 1 9370
box -6 -8 126 248
use INVX8  _8057_
timestamp 0
transform 1 0 1590 0 -1 9370
box -6 -8 126 248
use INVX1  _8058_
timestamp 0
transform 1 0 2390 0 1 11290
box -6 -8 66 248
use NAND2X1  _8059_
timestamp 0
transform 1 0 2650 0 1 11290
box -6 -8 86 248
use OAI21X1  _8060_
timestamp 0
transform 1 0 2510 0 1 11290
box -6 -8 106 248
use INVX1  _8061_
timestamp 0
transform 1 0 3510 0 1 10330
box -6 -8 66 248
use NAND2X1  _8062_
timestamp 0
transform -1 0 4030 0 1 10330
box -6 -8 86 248
use OAI21X1  _8063_
timestamp 0
transform 1 0 3790 0 1 10330
box -6 -8 106 248
use MUX2X1  _8064_
timestamp 0
transform 1 0 3630 0 1 10330
box -6 -8 126 248
use INVX1  _8065_
timestamp 0
transform 1 0 4170 0 1 9370
box -6 -8 66 248
use NAND2X1  _8066_
timestamp 0
transform 1 0 3810 0 -1 9850
box -6 -8 86 248
use OAI21X1  _8067_
timestamp 0
transform -1 0 4130 0 1 9370
box -6 -8 106 248
use INVX1  _8068_
timestamp 0
transform -1 0 2890 0 1 8890
box -6 -8 66 248
use NAND2X1  _8069_
timestamp 0
transform -1 0 3030 0 1 8890
box -6 -8 86 248
use OAI21X1  _8070_
timestamp 0
transform -1 0 3170 0 1 8890
box -6 -8 106 248
use MUX2X1  _8071_
timestamp 0
transform 1 0 3850 0 1 9370
box -6 -8 126 248
use MUX2X1  _8072_
timestamp 0
transform 1 0 3830 0 -1 10330
box -6 -8 126 248
use NOR2X1  _8073_
timestamp 0
transform -1 0 5210 0 1 9850
box -6 -8 86 248
use NAND2X1  _8074_
timestamp 0
transform 1 0 5270 0 1 9850
box -6 -8 86 248
use INVX1  _8075_
timestamp 0
transform -1 0 5190 0 -1 9850
box -6 -8 66 248
use NAND2X1  _8076_
timestamp 0
transform 1 0 5590 0 1 9370
box -6 -8 86 248
use OAI21X1  _8077_
timestamp 0
transform -1 0 4590 0 -1 10810
box -6 -8 106 248
use INVX2  _8078_
timestamp 0
transform -1 0 4450 0 -1 10810
box -6 -8 66 248
use OAI21X1  _8079_
timestamp 0
transform -1 0 5090 0 -1 9850
box -6 -8 106 248
use OAI21X1  _8080_
timestamp 0
transform 1 0 4730 0 1 8890
box -6 -8 106 248
use INVX8  _8081_
timestamp 0
transform 1 0 6870 0 -1 7930
box -6 -8 126 248
use NAND2X1  _8082_
timestamp 0
transform 1 0 4890 0 -1 8410
box -6 -8 86 248
use NOR2X1  _8083_
timestamp 0
transform 1 0 5250 0 1 10330
box -6 -8 86 248
use MUX2X1  _8084_
timestamp 0
transform -1 0 3010 0 1 9850
box -6 -8 126 248
use MUX2X1  _8085_
timestamp 0
transform -1 0 3170 0 1 9850
box -6 -8 126 248
use MUX2X1  _8086_
timestamp 0
transform -1 0 2750 0 -1 9850
box -6 -8 126 248
use INVX2  _8087_
timestamp 0
transform -1 0 3770 0 -1 8890
box -6 -8 66 248
use NAND2X1  _8088_
timestamp 0
transform 1 0 3690 0 -1 9850
box -6 -8 86 248
use AOI21X1  _8089_
timestamp 0
transform -1 0 3630 0 -1 9850
box -6 -8 106 248
use NAND3X1  _8090_
timestamp 0
transform 1 0 3270 0 -1 9370
box -6 -8 106 248
use NAND3X1  _8091_
timestamp 0
transform 1 0 3170 0 1 9370
box -6 -8 106 248
use NAND3X1  _8092_
timestamp 0
transform 1 0 3310 0 1 9370
box -6 -8 106 248
use OAI22X1  _8093_
timestamp 0
transform -1 0 3490 0 -1 9850
box -6 -8 126 248
use INVX1  _8094_
timestamp 0
transform -1 0 5810 0 1 10330
box -6 -8 66 248
use INVX8  _8095_
timestamp 0
transform -1 0 190 0 -1 8890
box -6 -8 126 248
use INVX1  _8096_
timestamp 0
transform -1 0 2810 0 -1 10810
box -6 -8 66 248
use NAND2X1  _8097_
timestamp 0
transform -1 0 2570 0 -1 9850
box -6 -8 86 248
use OAI21X1  _8098_
timestamp 0
transform -1 0 2830 0 -1 10330
box -6 -8 106 248
use INVX1  _8099_
timestamp 0
transform 1 0 3130 0 1 10330
box -6 -8 66 248
use NAND2X1  _8100_
timestamp 0
transform 1 0 3390 0 1 10330
box -6 -8 86 248
use OAI21X1  _8101_
timestamp 0
transform 1 0 3230 0 1 10330
box -6 -8 106 248
use MUX2X1  _8102_
timestamp 0
transform 1 0 3030 0 -1 10330
box -6 -8 126 248
use INVX1  _8103_
timestamp 0
transform -1 0 3290 0 1 9850
box -6 -8 66 248
use NAND2X1  _8104_
timestamp 0
transform 1 0 3350 0 -1 10330
box -6 -8 86 248
use OAI21X1  _8105_
timestamp 0
transform 1 0 3210 0 -1 10330
box -6 -8 106 248
use INVX1  _8106_
timestamp 0
transform -1 0 2710 0 -1 9370
box -6 -8 66 248
use NAND2X1  _8107_
timestamp 0
transform -1 0 2330 0 -1 9370
box -6 -8 86 248
use OAI21X1  _8108_
timestamp 0
transform -1 0 2470 0 -1 9370
box -6 -8 106 248
use MUX2X1  _8109_
timestamp 0
transform 1 0 3470 0 -1 10330
box -6 -8 126 248
use MUX2X1  _8110_
timestamp 0
transform -1 0 3770 0 -1 10330
box -6 -8 126 248
use NAND3X1  _8111_
timestamp 0
transform 1 0 4790 0 -1 10330
box -6 -8 106 248
use MUX2X1  _8112_
timestamp 0
transform -1 0 2270 0 1 9370
box -6 -8 126 248
use MUX2X1  _8113_
timestamp 0
transform -1 0 2450 0 -1 9850
box -6 -8 126 248
use MUX2X1  _8114_
timestamp 0
transform 1 0 2170 0 -1 9850
box -6 -8 126 248
use MUX2X1  _8115_
timestamp 0
transform -1 0 3630 0 1 9850
box -6 -8 126 248
use MUX2X1  _8116_
timestamp 0
transform 1 0 3190 0 -1 9850
box -6 -8 126 248
use MUX2X1  _8117_
timestamp 0
transform -1 0 3470 0 1 9850
box -6 -8 126 248
use MUX2X1  _8118_
timestamp 0
transform 1 0 3790 0 1 9850
box -6 -8 126 248
use OAI21X1  _8119_
timestamp 0
transform 1 0 4850 0 1 9850
box -6 -8 106 248
use AOI21X1  _8120_
timestamp 0
transform 1 0 5090 0 -1 10330
box -6 -8 106 248
use INVX1  _8121_
timestamp 0
transform 1 0 5370 0 -1 10330
box -6 -8 66 248
use NAND3X1  _8122_
timestamp 0
transform -1 0 5050 0 -1 10330
box -6 -8 106 248
use AND2X2  _8123_
timestamp 0
transform -1 0 5090 0 1 9850
box -6 -8 106 248
use OAI21X1  _8124_
timestamp 0
transform -1 0 4930 0 -1 9850
box -6 -8 106 248
use OR2X2  _8125_
timestamp 0
transform -1 0 4770 0 -1 9850
box -6 -8 106 248
use AOI21X1  _8126_
timestamp 0
transform -1 0 4630 0 -1 9850
box -6 -8 106 248
use OAI21X1  _8127_
timestamp 0
transform 1 0 4750 0 -1 8410
box -6 -8 106 248
use INVX1  _8128_
timestamp 0
transform 1 0 7050 0 1 6490
box -6 -8 66 248
use NAND2X1  _8129_
timestamp 0
transform 1 0 7230 0 -1 6490
box -6 -8 86 248
use OAI21X1  _8130_
timestamp 0
transform 1 0 7070 0 -1 6490
box -6 -8 106 248
use NAND2X1  _8131_
timestamp 0
transform 1 0 4530 0 1 9370
box -6 -8 86 248
use AOI21X1  _8132_
timestamp 0
transform 1 0 5230 0 -1 10330
box -6 -8 106 248
use MUX2X1  _8133_
timestamp 0
transform -1 0 2030 0 -1 8890
box -6 -8 126 248
use MUX2X1  _8134_
timestamp 0
transform -1 0 2110 0 -1 9850
box -6 -8 126 248
use MUX2X1  _8135_
timestamp 0
transform 1 0 4090 0 -1 9850
box -6 -8 126 248
use NAND2X1  _8136_
timestamp 0
transform -1 0 4170 0 1 9850
box -6 -8 86 248
use OAI22X1  _8137_
timestamp 0
transform 1 0 4210 0 1 9850
box -6 -8 126 248
use AOI21X1  _8138_
timestamp 0
transform 1 0 4390 0 1 9850
box -6 -8 106 248
use AOI21X1  _8139_
timestamp 0
transform -1 0 4790 0 1 9850
box -6 -8 106 248
use NAND2X1  _8140_
timestamp 0
transform 1 0 4670 0 -1 10330
box -6 -8 86 248
use INVX1  _8141_
timestamp 0
transform -1 0 4350 0 -1 10330
box -6 -8 66 248
use OAI21X1  _8142_
timestamp 0
transform 1 0 4530 0 -1 10330
box -6 -8 106 248
use NAND2X1  _8143_
timestamp 0
transform 1 0 4410 0 -1 10330
box -6 -8 86 248
use AOI21X1  _8144_
timestamp 0
transform 1 0 4970 0 1 10330
box -6 -8 106 248
use NAND3X1  _8145_
timestamp 0
transform -1 0 4930 0 1 10330
box -6 -8 106 248
use INVX1  _8146_
timestamp 0
transform -1 0 4850 0 -1 10810
box -6 -8 66 248
use OR2X2  _8147_
timestamp 0
transform 1 0 5050 0 -1 10810
box -6 -8 106 248
use NOR2X1  _8148_
timestamp 0
transform 1 0 5310 0 -1 10810
box -6 -8 86 248
use INVX1  _8149_
timestamp 0
transform -1 0 5250 0 -1 10810
box -6 -8 66 248
use OAI21X1  _8150_
timestamp 0
transform 1 0 4910 0 -1 10810
box -6 -8 106 248
use AOI21X1  _8151_
timestamp 0
transform -1 0 5210 0 1 10330
box -6 -8 106 248
use INVX2  _8152_
timestamp 0
transform -1 0 1150 0 -1 9370
box -6 -8 66 248
use OAI21X1  _8153_
timestamp 0
transform 1 0 3950 0 -1 9850
box -6 -8 106 248
use OAI21X1  _8154_
timestamp 0
transform 1 0 4370 0 1 9370
box -6 -8 106 248
use INVX1  _8155_
timestamp 0
transform 1 0 3590 0 1 11290
box -6 -8 66 248
use INVX2  _8156_
timestamp 0
transform -1 0 4330 0 1 9370
box -6 -8 66 248
use OAI21X1  _8157_
timestamp 0
transform -1 0 4750 0 -1 10810
box -6 -8 106 248
use INVX1  _8158_
timestamp 0
transform 1 0 2970 0 -1 11770
box -6 -8 66 248
use INVX1  _8159_
timestamp 0
transform -1 0 2630 0 -1 11770
box -6 -8 66 248
use NAND3X1  _8160_
timestamp 0
transform -1 0 4650 0 1 9850
box -6 -8 106 248
use INVX1  _8161_
timestamp 0
transform -1 0 1950 0 1 7930
box -6 -8 66 248
use NAND2X1  _8162_
timestamp 0
transform -1 0 1650 0 -1 7450
box -6 -8 86 248
use OAI21X1  _8163_
timestamp 0
transform -1 0 1690 0 1 7450
box -6 -8 106 248
use NAND2X1  _8164_
timestamp 0
transform 1 0 1870 0 1 9370
box -6 -8 86 248
use OAI21X1  _8165_
timestamp 0
transform 1 0 1590 0 1 9370
box -6 -8 106 248
use NOR2X1  _8166_
timestamp 0
transform -1 0 1450 0 -1 10330
box -6 -8 86 248
use NOR2X1  _8167_
timestamp 0
transform 1 0 5990 0 1 10330
box -6 -8 86 248
use AOI22X1  _8168_
timestamp 0
transform -1 0 2990 0 -1 10330
box -6 -8 126 248
use OAI21X1  _8169_
timestamp 0
transform 1 0 1610 0 1 9850
box -6 -8 106 248
use NAND3X1  _8170_
timestamp 0
transform 1 0 1430 0 -1 11770
box -6 -8 106 248
use INVX1  _8171_
timestamp 0
transform 1 0 770 0 1 11290
box -6 -8 66 248
use INVX1  _8172_
timestamp 0
transform 1 0 1030 0 1 11290
box -6 -8 66 248
use OAI21X1  _8173_
timestamp 0
transform 1 0 870 0 1 11290
box -6 -8 106 248
use NAND3X1  _8174_
timestamp 0
transform 1 0 2010 0 -1 11770
box -6 -8 106 248
use AOI21X1  _8175_
timestamp 0
transform 1 0 2150 0 -1 11770
box -6 -8 106 248
use INVX1  _8176_
timestamp 0
transform 1 0 2390 0 1 11770
box -6 -8 66 248
use NAND2X1  _8177_
timestamp 0
transform -1 0 2530 0 -1 11770
box -6 -8 86 248
use AOI21X1  _8178_
timestamp 0
transform 1 0 2670 0 -1 11770
box -6 -8 106 248
use OAI21X1  _8179_
timestamp 0
transform -1 0 2930 0 -1 11770
box -6 -8 106 248
use AOI22X1  _8180_
timestamp 0
transform -1 0 3530 0 1 11290
box -6 -8 126 248
use AOI21X1  _8181_
timestamp 0
transform -1 0 2410 0 -1 11770
box -6 -8 106 248
use INVX1  _8182_
timestamp 0
transform 1 0 1750 0 1 11770
box -6 -8 66 248
use INVX1  _8183_
timestamp 0
transform -1 0 770 0 -1 6970
box -6 -8 66 248
use NAND2X1  _8184_
timestamp 0
transform -1 0 530 0 -1 6970
box -6 -8 86 248
use OAI21X1  _8185_
timestamp 0
transform -1 0 670 0 -1 6970
box -6 -8 106 248
use NAND2X1  _8186_
timestamp 0
transform -1 0 1830 0 1 9370
box -6 -8 86 248
use OAI21X1  _8187_
timestamp 0
transform 1 0 710 0 1 9370
box -6 -8 106 248
use NAND2X1  _8188_
timestamp 0
transform 1 0 1690 0 -1 9850
box -6 -8 86 248
use OAI21X1  _8189_
timestamp 0
transform -1 0 810 0 -1 9850
box -6 -8 106 248
use INVX2  _8190_
timestamp 0
transform 1 0 750 0 -1 11290
box -6 -8 66 248
use OAI21X1  _8191_
timestamp 0
transform 1 0 830 0 -1 11770
box -6 -8 106 248
use OR2X2  _8192_
timestamp 0
transform -1 0 390 0 -1 12250
box -6 -8 106 248
use NOR2X1  _8193_
timestamp 0
transform -1 0 950 0 -1 11290
box -6 -8 86 248
use OAI21X1  _8194_
timestamp 0
transform -1 0 730 0 1 11290
box -6 -8 106 248
use NAND3X1  _8195_
timestamp 0
transform 1 0 730 0 1 11770
box -6 -8 106 248
use NOR2X1  _8196_
timestamp 0
transform 1 0 590 0 -1 12250
box -6 -8 86 248
use AND2X2  _8197_
timestamp 0
transform 1 0 430 0 -1 12250
box -6 -8 106 248
use OAI21X1  _8198_
timestamp 0
transform 1 0 730 0 -1 12250
box -6 -8 106 248
use NAND2X1  _8199_
timestamp 0
transform 1 0 1010 0 1 11770
box -6 -8 86 248
use AOI21X1  _8200_
timestamp 0
transform 1 0 1150 0 -1 11770
box -6 -8 106 248
use OAI21X1  _8201_
timestamp 0
transform 1 0 1290 0 -1 11770
box -6 -8 106 248
use AOI22X1  _8202_
timestamp 0
transform -1 0 2930 0 1 8410
box -6 -8 126 248
use OAI21X1  _8203_
timestamp 0
transform -1 0 1090 0 -1 11770
box -6 -8 106 248
use INVX1  _8204_
timestamp 0
transform -1 0 1470 0 1 11770
box -6 -8 66 248
use NAND3X1  _8205_
timestamp 0
transform -1 0 590 0 1 11290
box -6 -8 106 248
use NAND2X1  _8206_
timestamp 0
transform -1 0 870 0 1 6970
box -6 -8 86 248
use INVX1  _8207_
timestamp 0
transform 1 0 1050 0 1 7930
box -6 -8 66 248
use AOI21X1  _8208_
timestamp 0
transform -1 0 870 0 -1 9370
box -6 -8 106 248
use NAND2X1  _8209_
timestamp 0
transform 1 0 1070 0 1 9850
box -6 -8 86 248
use OAI21X1  _8210_
timestamp 0
transform 1 0 570 0 -1 9850
box -6 -8 106 248
use NAND3X1  _8211_
timestamp 0
transform -1 0 150 0 1 11290
box -6 -8 106 248
use NOR3X1  _8212_
timestamp 0
transform -1 0 870 0 1 10810
box -6 -8 186 248
use INVX1  _8213_
timestamp 0
transform -1 0 570 0 -1 11290
box -6 -8 66 248
use OAI21X1  _8214_
timestamp 0
transform -1 0 470 0 -1 11290
box -6 -8 106 248
use NAND3X1  _8215_
timestamp 0
transform 1 0 70 0 -1 11770
box -6 -8 106 248
use AOI21X1  _8216_
timestamp 0
transform 1 0 50 0 1 11770
box -6 -8 106 248
use INVX1  _8217_
timestamp 0
transform 1 0 210 0 1 11770
box -6 -8 66 248
use NAND2X1  _8218_
timestamp 0
transform 1 0 190 0 1 11290
box -6 -8 86 248
use AND2X2  _8219_
timestamp 0
transform 1 0 1150 0 -1 11290
box -6 -8 106 248
use OAI21X1  _8220_
timestamp 0
transform -1 0 1090 0 -1 11290
box -6 -8 106 248
use OAI21X1  _8221_
timestamp 0
transform 1 0 1290 0 -1 11290
box -6 -8 106 248
use OAI21X1  _8222_
timestamp 0
transform -1 0 2610 0 1 7930
box -6 -8 106 248
use INVX1  _8223_
timestamp 0
transform -1 0 2210 0 1 7930
box -6 -8 66 248
use INVX1  _8224_
timestamp 0
transform 1 0 530 0 -1 10810
box -6 -8 66 248
use NAND3X1  _8225_
timestamp 0
transform 1 0 610 0 -1 11290
box -6 -8 106 248
use AOI21X1  _8226_
timestamp 0
transform -1 0 730 0 -1 9370
box -6 -8 106 248
use NAND2X1  _8227_
timestamp 0
transform 1 0 430 0 -1 9850
box -6 -8 86 248
use OAI21X1  _8228_
timestamp 0
transform -1 0 390 0 -1 9850
box -6 -8 106 248
use NAND3X1  _8229_
timestamp 0
transform -1 0 170 0 -1 10810
box -6 -8 106 248
use INVX1  _8230_
timestamp 0
transform 1 0 170 0 1 10810
box -6 -8 66 248
use OAI21X1  _8231_
timestamp 0
transform -1 0 430 0 1 11290
box -6 -8 106 248
use NAND2X1  _8232_
timestamp 0
transform 1 0 270 0 1 10810
box -6 -8 86 248
use NAND3X1  _8233_
timestamp 0
transform 1 0 370 0 -1 10810
box -6 -8 106 248
use NAND3X1  _8234_
timestamp 0
transform -1 0 170 0 -1 11290
box -6 -8 106 248
use NAND2X1  _8235_
timestamp 0
transform 1 0 390 0 1 10810
box -6 -8 86 248
use NAND3X1  _8236_
timestamp 0
transform 1 0 530 0 1 10810
box -6 -8 106 248
use NAND2X1  _8237_
timestamp 0
transform 1 0 730 0 1 10330
box -6 -8 86 248
use AOI21X1  _8238_
timestamp 0
transform -1 0 690 0 1 11770
box -6 -8 106 248
use NOR2X1  _8239_
timestamp 0
transform -1 0 530 0 1 11770
box -6 -8 86 248
use OAI21X1  _8240_
timestamp 0
transform -1 0 770 0 -1 11770
box -6 -8 106 248
use NAND2X1  _8241_
timestamp 0
transform 1 0 550 0 -1 11770
box -6 -8 86 248
use AOI21X1  _8242_
timestamp 0
transform 1 0 1150 0 1 10330
box -6 -8 106 248
use OAI21X1  _8243_
timestamp 0
transform 1 0 1230 0 -1 10330
box -6 -8 106 248
use AOI22X1  _8244_
timestamp 0
transform -1 0 2110 0 1 7930
box -6 -8 126 248
use INVX1  _8245_
timestamp 0
transform -1 0 2870 0 -1 8410
box -6 -8 66 248
use AOI21X1  _8246_
timestamp 0
transform -1 0 330 0 -1 10810
box -6 -8 106 248
use AND2X2  _8247_
timestamp 0
transform -1 0 970 0 1 11770
box -6 -8 106 248
use NAND3X1  _8248_
timestamp 0
transform 1 0 230 0 -1 11770
box -6 -8 106 248
use AOI21X1  _8249_
timestamp 0
transform -1 0 410 0 1 11770
box -6 -8 106 248
use OAI21X1  _8250_
timestamp 0
transform -1 0 490 0 -1 11770
box -6 -8 106 248
use AOI21X1  _8251_
timestamp 0
transform 1 0 450 0 1 10330
box -6 -8 106 248
use INVX1  _8252_
timestamp 0
transform -1 0 250 0 -1 9850
box -6 -8 66 248
use NAND3X1  _8253_
timestamp 0
transform -1 0 330 0 -1 11290
box -6 -8 106 248
use INVX1  _8254_
timestamp 0
transform 1 0 690 0 1 6970
box -6 -8 66 248
use NOR2X1  _8255_
timestamp 0
transform -1 0 890 0 -1 8890
box -6 -8 86 248
use INVX1  _8256_
timestamp 0
transform 1 0 910 0 1 8890
box -6 -8 66 248
use OAI21X1  _8257_
timestamp 0
transform -1 0 970 0 1 9370
box -6 -8 106 248
use NAND3X1  _8258_
timestamp 0
transform 1 0 390 0 1 9850
box -6 -8 106 248
use INVX1  _8259_
timestamp 0
transform -1 0 110 0 1 9850
box -6 -8 66 248
use OAI21X1  _8260_
timestamp 0
transform 1 0 190 0 1 10330
box -6 -8 106 248
use NAND2X1  _8261_
timestamp 0
transform 1 0 150 0 1 9850
box -6 -8 86 248
use NAND3X1  _8262_
timestamp 0
transform 1 0 550 0 1 9850
box -6 -8 106 248
use NAND3X1  _8263_
timestamp 0
transform 1 0 50 0 -1 10330
box -6 -8 106 248
use NAND2X1  _8264_
timestamp 0
transform -1 0 350 0 1 9850
box -6 -8 86 248
use NAND3X1  _8265_
timestamp 0
transform 1 0 210 0 -1 10330
box -6 -8 106 248
use NAND2X1  _8266_
timestamp 0
transform 1 0 810 0 -1 10330
box -6 -8 86 248
use INVX1  _8267_
timestamp 0
transform -1 0 890 0 1 9850
box -6 -8 66 248
use NOR2X1  _8268_
timestamp 0
transform -1 0 770 0 1 9850
box -6 -8 86 248
use OAI21X1  _8269_
timestamp 0
transform -1 0 970 0 1 10330
box -6 -8 106 248
use OAI21X1  _8270_
timestamp 0
transform 1 0 930 0 1 9850
box -6 -8 106 248
use OAI21X1  _8271_
timestamp 0
transform -1 0 2610 0 -1 8410
box -6 -8 106 248
use INVX1  _8272_
timestamp 0
transform -1 0 2250 0 1 8410
box -6 -8 66 248
use OAI21X1  _8273_
timestamp 0
transform 1 0 1010 0 1 9370
box -6 -8 106 248
use OAI21X1  _8274_
timestamp 0
transform -1 0 2770 0 -1 8410
box -6 -8 106 248
use INVX1  _8275_
timestamp 0
transform -1 0 2350 0 1 8410
box -6 -8 66 248
use OAI21X1  _8276_
timestamp 0
transform 1 0 930 0 -1 10330
box -6 -8 106 248
use NOR2X1  _8277_
timestamp 0
transform -1 0 1110 0 1 10330
box -6 -8 86 248
use AOI21X1  _8278_
timestamp 0
transform 1 0 1070 0 -1 10330
box -6 -8 106 248
use INVX1  _8279_
timestamp 0
transform -1 0 470 0 -1 8890
box -6 -8 66 248
use OR2X2  _8280_
timestamp 0
transform -1 0 150 0 -1 9850
box -6 -8 106 248
use OAI21X1  _8281_
timestamp 0
transform -1 0 670 0 1 9370
box -6 -8 106 248
use NAND3X1  _8282_
timestamp 0
transform 1 0 190 0 1 8890
box -6 -8 106 248
use NOR2X1  _8283_
timestamp 0
transform -1 0 130 0 1 9370
box -6 -8 86 248
use INVX1  _8284_
timestamp 0
transform -1 0 130 0 -1 9370
box -6 -8 66 248
use OAI21X1  _8285_
timestamp 0
transform -1 0 150 0 1 8890
box -6 -8 106 248
use NAND3X1  _8286_
timestamp 0
transform -1 0 350 0 -1 8890
box -6 -8 106 248
use NAND3X1  _8287_
timestamp 0
transform 1 0 170 0 -1 9370
box -6 -8 106 248
use OAI21X1  _8288_
timestamp 0
transform 1 0 350 0 1 8890
box -6 -8 106 248
use NAND3X1  _8289_
timestamp 0
transform 1 0 490 0 1 8890
box -6 -8 106 248
use AND2X2  _8290_
timestamp 0
transform 1 0 510 0 -1 8890
box -6 -8 106 248
use INVX1  _8291_
timestamp 0
transform 1 0 1070 0 -1 8410
box -6 -8 66 248
use AOI21X1  _8292_
timestamp 0
transform 1 0 1410 0 -1 8410
box -6 -8 106 248
use OAI21X1  _8293_
timestamp 0
transform 1 0 1570 0 -1 8410
box -6 -8 106 248
use AOI22X1  _8294_
timestamp 0
transform -1 0 2130 0 1 8410
box -6 -8 126 248
use NAND2X1  _8295_
timestamp 0
transform 1 0 330 0 1 10330
box -6 -8 86 248
use AND2X2  _8296_
timestamp 0
transform 1 0 370 0 -1 10330
box -6 -8 106 248
use AND2X2  _8297_
timestamp 0
transform 1 0 590 0 1 10330
box -6 -8 106 248
use NAND3X1  _8298_
timestamp 0
transform -1 0 770 0 -1 10330
box -6 -8 106 248
use OAI21X1  _8299_
timestamp 0
transform -1 0 610 0 -1 10330
box -6 -8 106 248
use INVX1  _8300_
timestamp 0
transform 1 0 650 0 1 8890
box -6 -8 66 248
use AOI21X1  _8301_
timestamp 0
transform 1 0 650 0 -1 8890
box -6 -8 106 248
use INVX1  _8302_
timestamp 0
transform -1 0 1070 0 1 8410
box -6 -8 66 248
use NOR3X1  _8303_
timestamp 0
transform 1 0 190 0 1 9370
box -6 -8 186 248
use INVX1  _8304_
timestamp 0
transform -1 0 250 0 1 8410
box -6 -8 66 248
use OAI21X1  _8305_
timestamp 0
transform 1 0 770 0 1 8890
box -6 -8 106 248
use NAND3X1  _8306_
timestamp 0
transform 1 0 50 0 1 8410
box -6 -8 106 248
use INVX1  _8307_
timestamp 0
transform -1 0 110 0 -1 8410
box -6 -8 66 248
use OAI21X1  _8308_
timestamp 0
transform -1 0 410 0 1 8410
box -6 -8 106 248
use NAND3X1  _8309_
timestamp 0
transform -1 0 550 0 1 8410
box -6 -8 106 248
use NAND3X1  _8310_
timestamp 0
transform 1 0 170 0 -1 8410
box -6 -8 106 248
use OAI21X1  _8311_
timestamp 0
transform 1 0 310 0 -1 8410
box -6 -8 106 248
use NAND3X1  _8312_
timestamp 0
transform 1 0 470 0 -1 8410
box -6 -8 106 248
use AND2X2  _8313_
timestamp 0
transform 1 0 610 0 -1 8410
box -6 -8 106 248
use AND2X2  _8314_
timestamp 0
transform 1 0 1150 0 1 7930
box -6 -8 106 248
use OAI21X1  _8315_
timestamp 0
transform 1 0 1310 0 1 7930
box -6 -8 106 248
use OAI21X1  _8316_
timestamp 0
transform 1 0 1450 0 1 7930
box -6 -8 106 248
use OAI21X1  _8317_
timestamp 0
transform -1 0 3330 0 1 6970
box -6 -8 106 248
use INVX1  _8318_
timestamp 0
transform 1 0 470 0 1 7450
box -6 -8 66 248
use OAI21X1  _8319_
timestamp 0
transform 1 0 470 0 -1 9370
box -6 -8 106 248
use INVX1  _8320_
timestamp 0
transform 1 0 490 0 1 7930
box -6 -8 66 248
use AOI21X1  _8321_
timestamp 0
transform -1 0 290 0 1 7930
box -6 -8 106 248
use NAND3X1  _8322_
timestamp 0
transform 1 0 350 0 1 7930
box -6 -8 106 248
use NAND2X1  _8323_
timestamp 0
transform -1 0 250 0 -1 7930
box -6 -8 86 248
use NAND2X1  _8324_
timestamp 0
transform -1 0 690 0 1 7930
box -6 -8 86 248
use OAI21X1  _8325_
timestamp 0
transform 1 0 290 0 -1 7930
box -6 -8 106 248
use NAND2X1  _8326_
timestamp 0
transform -1 0 510 0 -1 7930
box -6 -8 86 248
use INVX1  _8327_
timestamp 0
transform -1 0 130 0 -1 7930
box -6 -8 66 248
use AND2X2  _8328_
timestamp 0
transform -1 0 290 0 1 7450
box -6 -8 106 248
use NAND2X1  _8329_
timestamp 0
transform -1 0 150 0 1 7450
box -6 -8 86 248
use NAND3X1  _8330_
timestamp 0
transform -1 0 430 0 1 7450
box -6 -8 106 248
use NAND2X1  _8331_
timestamp 0
transform -1 0 650 0 -1 7930
box -6 -8 86 248
use AOI21X1  _8332_
timestamp 0
transform 1 0 590 0 1 8410
box -6 -8 106 248
use AOI21X1  _8333_
timestamp 0
transform 1 0 730 0 1 8410
box -6 -8 106 248
use NAND3X1  _8334_
timestamp 0
transform 1 0 750 0 1 7930
box -6 -8 106 248
use AOI21X1  _8335_
timestamp 0
transform 1 0 890 0 1 7930
box -6 -8 106 248
use AND2X2  _8336_
timestamp 0
transform 1 0 710 0 -1 7930
box -6 -8 106 248
use NAND3X1  _8337_
timestamp 0
transform 1 0 750 0 -1 8410
box -6 -8 106 248
use OAI21X1  _8338_
timestamp 0
transform 1 0 910 0 -1 8410
box -6 -8 106 248
use OAI21X1  _8339_
timestamp 0
transform 1 0 990 0 -1 7930
box -6 -8 106 248
use OR2X2  _8340_
timestamp 0
transform 1 0 1130 0 -1 7930
box -6 -8 106 248
use AOI22X1  _8341_
timestamp 0
transform -1 0 3030 0 -1 7930
box -6 -8 126 248
use NAND2X1  _8342_
timestamp 0
transform 1 0 3530 0 -1 7450
box -6 -8 86 248
use INVX1  _8343_
timestamp 0
transform -1 0 650 0 1 7450
box -6 -8 66 248
use NAND2X1  _8344_
timestamp 0
transform -1 0 770 0 -1 7450
box -6 -8 86 248
use INVX1  _8345_
timestamp 0
transform 1 0 810 0 -1 7450
box -6 -8 66 248
use NAND2X1  _8346_
timestamp 0
transform 1 0 570 0 -1 7450
box -6 -8 86 248
use NAND2X1  _8347_
timestamp 0
transform -1 0 510 0 -1 7450
box -6 -8 86 248
use INVX1  _8348_
timestamp 0
transform -1 0 250 0 1 6970
box -6 -8 66 248
use NAND2X1  _8349_
timestamp 0
transform -1 0 270 0 -1 7450
box -6 -8 86 248
use NAND2X1  _8350_
timestamp 0
transform -1 0 150 0 -1 7450
box -6 -8 86 248
use NAND2X1  _8351_
timestamp 0
transform 1 0 310 0 -1 7450
box -6 -8 86 248
use INVX1  _8352_
timestamp 0
transform -1 0 750 0 1 7450
box -6 -8 66 248
use NOR3X1  _8353_
timestamp 0
transform 1 0 810 0 1 7450
box -6 -8 186 248
use AOI21X1  _8354_
timestamp 0
transform -1 0 950 0 -1 7930
box -6 -8 106 248
use OAI21X1  _8355_
timestamp 0
transform 1 0 1290 0 -1 7930
box -6 -8 106 248
use OAI21X1  _8356_
timestamp 0
transform 1 0 1430 0 -1 7930
box -6 -8 106 248
use NAND2X1  _8357_
timestamp 0
transform -1 0 3250 0 -1 7450
box -6 -8 86 248
use NAND2X1  _8358_
timestamp 0
transform 1 0 3410 0 -1 8410
box -6 -8 86 248
use INVX1  _8359_
timestamp 0
transform 1 0 4590 0 1 10330
box -6 -8 66 248
use NAND2X1  _8360_
timestamp 0
transform -1 0 4410 0 1 10330
box -6 -8 86 248
use OAI21X1  _8361_
timestamp 0
transform -1 0 4550 0 1 10330
box -6 -8 106 248
use NAND2X1  _8362_
timestamp 0
transform 1 0 4150 0 -1 10330
box -6 -8 86 248
use NOR2X1  _8363_
timestamp 0
transform 1 0 5850 0 1 10330
box -6 -8 86 248
use NOR2X1  _8364_
timestamp 0
transform -1 0 5310 0 -1 9850
box -6 -8 86 248
use AOI22X1  _8365_
timestamp 0
transform 1 0 5730 0 -1 10330
box -6 -8 126 248
use NAND3X1  _8366_
timestamp 0
transform -1 0 4090 0 -1 10330
box -6 -8 106 248
use NAND2X1  _8367_
timestamp 0
transform 1 0 790 0 -1 10810
box -6 -8 86 248
use OAI21X1  _8368_
timestamp 0
transform 1 0 630 0 -1 10810
box -6 -8 106 248
use NAND2X1  _8369_
timestamp 0
transform 1 0 1290 0 1 11770
box -6 -8 86 248
use OAI21X1  _8370_
timestamp 0
transform -1 0 1230 0 1 11770
box -6 -8 106 248
use MUX2X1  _8371_
timestamp 0
transform 1 0 1290 0 -1 10810
box -6 -8 126 248
use NAND2X1  _8372_
timestamp 0
transform -1 0 1830 0 -1 10810
box -6 -8 86 248
use AND2X2  _8373_
timestamp 0
transform -1 0 2830 0 1 9850
box -6 -8 106 248
use NOR2X1  _8374_
timestamp 0
transform -1 0 2790 0 1 8890
box -6 -8 86 248
use NAND2X1  _8375_
timestamp 0
transform 1 0 1170 0 -1 10810
box -6 -8 86 248
use NAND2X1  _8376_
timestamp 0
transform -1 0 990 0 -1 10810
box -6 -8 86 248
use NAND2X1  _8377_
timestamp 0
transform -1 0 1130 0 -1 10810
box -6 -8 86 248
use OAI21X1  _8378_
timestamp 0
transform 1 0 2030 0 1 9850
box -6 -8 106 248
use OAI21X1  _8379_
timestamp 0
transform 1 0 2890 0 -1 8890
box -6 -8 106 248
use OAI21X1  _8380_
timestamp 0
transform 1 0 2970 0 1 8410
box -6 -8 106 248
use NAND2X1  _8381_
timestamp 0
transform -1 0 2870 0 1 7450
box -6 -8 86 248
use NOR2X1  _8382_
timestamp 0
transform -1 0 2830 0 -1 8890
box -6 -8 86 248
use NAND2X1  _8383_
timestamp 0
transform 1 0 1850 0 1 11770
box -6 -8 86 248
use OAI21X1  _8384_
timestamp 0
transform -1 0 1950 0 -1 11770
box -6 -8 106 248
use NAND2X1  _8385_
timestamp 0
transform -1 0 5450 0 1 10330
box -6 -8 86 248
use OAI21X1  _8386_
timestamp 0
transform -1 0 5610 0 1 10330
box -6 -8 106 248
use MUX2X1  _8387_
timestamp 0
transform 1 0 2970 0 1 10330
box -6 -8 126 248
use NAND2X1  _8388_
timestamp 0
transform 1 0 1910 0 1 9850
box -6 -8 86 248
use NAND2X1  _8389_
timestamp 0
transform -1 0 410 0 -1 9370
box -6 -8 86 248
use OAI21X1  _8390_
timestamp 0
transform -1 0 510 0 1 9370
box -6 -8 106 248
use INVX1  _8391_
timestamp 0
transform 1 0 870 0 -1 9850
box -6 -8 66 248
use NAND2X1  _8392_
timestamp 0
transform -1 0 990 0 1 10810
box -6 -8 86 248
use OAI21X1  _8393_
timestamp 0
transform -1 0 1150 0 1 10810
box -6 -8 106 248
use NAND2X1  _8394_
timestamp 0
transform -1 0 1190 0 -1 9850
box -6 -8 86 248
use OAI21X1  _8395_
timestamp 0
transform -1 0 1070 0 -1 9850
box -6 -8 106 248
use OAI21X1  _8396_
timestamp 0
transform 1 0 1770 0 1 9850
box -6 -8 106 248
use NAND3X1  _8397_
timestamp 0
transform 1 0 2510 0 -1 9370
box -6 -8 106 248
use MUX2X1  _8398_
timestamp 0
transform 1 0 1250 0 -1 9850
box -6 -8 126 248
use MUX2X1  _8399_
timestamp 0
transform -1 0 1930 0 -1 9850
box -6 -8 126 248
use OAI21X1  _8400_
timestamp 0
transform -1 0 2730 0 1 9370
box -6 -8 106 248
use AOI21X1  _8401_
timestamp 0
transform 1 0 2550 0 1 8890
box -6 -8 106 248
use INVX1  _8402_
timestamp 0
transform 1 0 2650 0 -1 8890
box -6 -8 66 248
use NAND3X1  _8403_
timestamp 0
transform -1 0 2510 0 1 8890
box -6 -8 106 248
use AND2X2  _8404_
timestamp 0
transform -1 0 2610 0 -1 8890
box -6 -8 106 248
use NAND2X1  _8405_
timestamp 0
transform -1 0 2490 0 1 8410
box -6 -8 86 248
use OR2X2  _8406_
timestamp 0
transform 1 0 2530 0 1 8410
box -6 -8 106 248
use AOI21X1  _8407_
timestamp 0
transform 1 0 2670 0 1 8410
box -6 -8 106 248
use OAI21X1  _8408_
timestamp 0
transform -1 0 2730 0 1 7450
box -6 -8 106 248
use NAND2X1  _8409_
timestamp 0
transform -1 0 3650 0 -1 7930
box -6 -8 86 248
use AOI21X1  _8410_
timestamp 0
transform -1 0 2470 0 -1 8890
box -6 -8 106 248
use NAND2X1  _8411_
timestamp 0
transform 1 0 2330 0 1 9850
box -6 -8 86 248
use NAND2X1  _8412_
timestamp 0
transform -1 0 1110 0 1 8890
box -6 -8 86 248
use OAI21X1  _8413_
timestamp 0
transform 1 0 1150 0 1 8890
box -6 -8 106 248
use NAND2X1  _8414_
timestamp 0
transform -1 0 1370 0 1 10330
box -6 -8 86 248
use OAI21X1  _8415_
timestamp 0
transform -1 0 1530 0 1 10330
box -6 -8 106 248
use NAND2X1  _8416_
timestamp 0
transform 1 0 4070 0 1 10330
box -6 -8 86 248
use NAND2X1  _8417_
timestamp 0
transform 1 0 1470 0 -1 10810
box -6 -8 86 248
use NAND2X1  _8418_
timestamp 0
transform -1 0 1650 0 1 10330
box -6 -8 86 248
use AOI21X1  _8419_
timestamp 0
transform 1 0 1630 0 -1 10330
box -6 -8 106 248
use INVX1  _8420_
timestamp 0
transform 1 0 2070 0 -1 10330
box -6 -8 66 248
use NAND3X1  _8421_
timestamp 0
transform 1 0 2310 0 -1 10330
box -6 -8 106 248
use AOI21X1  _8422_
timestamp 0
transform 1 0 2190 0 1 9850
box -6 -8 106 248
use OAI21X1  _8423_
timestamp 0
transform -1 0 2690 0 1 9850
box -6 -8 106 248
use NAND3X1  _8424_
timestamp 0
transform -1 0 2430 0 1 9370
box -6 -8 106 248
use INVX1  _8425_
timestamp 0
transform 1 0 1990 0 -1 9370
box -6 -8 66 248
use AOI21X1  _8426_
timestamp 0
transform 1 0 2470 0 1 9370
box -6 -8 106 248
use NOR2X1  _8427_
timestamp 0
transform -1 0 2210 0 1 8890
box -6 -8 86 248
use AND2X2  _8428_
timestamp 0
transform 1 0 2250 0 1 8890
box -6 -8 106 248
use NOR2X1  _8429_
timestamp 0
transform -1 0 2170 0 -1 8890
box -6 -8 86 248
use OAI21X1  _8430_
timestamp 0
transform 1 0 2210 0 -1 8890
box -6 -8 106 248
use OAI21X1  _8431_
timestamp 0
transform 1 0 3430 0 -1 7930
box -6 -8 106 248
use OAI21X1  _8432_
timestamp 0
transform -1 0 2190 0 -1 9370
box -6 -8 106 248
use INVX1  _8433_
timestamp 0
transform -1 0 1810 0 -1 9370
box -6 -8 66 248
use NAND2X1  _8434_
timestamp 0
transform -1 0 970 0 1 8410
box -6 -8 86 248
use OAI21X1  _8435_
timestamp 0
transform -1 0 1030 0 -1 8890
box -6 -8 106 248
use MUX2X1  _8436_
timestamp 0
transform 1 0 930 0 -1 9370
box -6 -8 126 248
use NOR2X1  _8437_
timestamp 0
transform -1 0 1490 0 -1 9850
box -6 -8 86 248
use NAND2X1  _8438_
timestamp 0
transform -1 0 2930 0 1 10330
box -6 -8 86 248
use NAND2X1  _8439_
timestamp 0
transform 1 0 1710 0 1 10330
box -6 -8 86 248
use NAND2X1  _8440_
timestamp 0
transform -1 0 1910 0 1 10330
box -6 -8 86 248
use OR2X2  _8441_
timestamp 0
transform -1 0 2070 0 1 10330
box -6 -8 106 248
use OAI21X1  _8442_
timestamp 0
transform -1 0 2270 0 -1 10330
box -6 -8 106 248
use OR2X2  _8443_
timestamp 0
transform 1 0 2270 0 1 10330
box -6 -8 106 248
use OAI21X1  _8444_
timestamp 0
transform 1 0 2110 0 1 10330
box -6 -8 106 248
use AOI21X1  _8445_
timestamp 0
transform 1 0 2550 0 1 10330
box -6 -8 106 248
use INVX1  _8446_
timestamp 0
transform -1 0 2670 0 -1 10330
box -6 -8 66 248
use NAND3X1  _8447_
timestamp 0
transform -1 0 2510 0 1 10330
box -6 -8 106 248
use NAND2X1  _8448_
timestamp 0
transform -1 0 2550 0 -1 10330
box -6 -8 86 248
use OR2X2  _8449_
timestamp 0
transform 1 0 1850 0 -1 9370
box -6 -8 106 248
use NAND2X1  _8450_
timestamp 0
transform 1 0 1870 0 1 8890
box -6 -8 86 248
use NAND2X1  _8451_
timestamp 0
transform 1 0 1990 0 1 8890
box -6 -8 86 248
use AOI22X1  _8452_
timestamp 0
transform -1 0 2510 0 -1 7930
box -6 -8 126 248
use AOI21X1  _8453_
timestamp 0
transform 1 0 2710 0 1 10330
box -6 -8 106 248
use NAND2X1  _8454_
timestamp 0
transform -1 0 1110 0 1 7450
box -6 -8 86 248
use OAI21X1  _8455_
timestamp 0
transform 1 0 1170 0 1 7450
box -6 -8 106 248
use NAND2X1  _8456_
timestamp 0
transform -1 0 1530 0 1 8890
box -6 -8 86 248
use OAI21X1  _8457_
timestamp 0
transform -1 0 1670 0 1 8890
box -6 -8 106 248
use NAND2X1  _8458_
timestamp 0
transform 1 0 1730 0 1 8890
box -6 -8 86 248
use OAI21X1  _8459_
timestamp 0
transform 1 0 1590 0 -1 10810
box -6 -8 106 248
use INVX1  _8460_
timestamp 0
transform 1 0 2210 0 1 10810
box -6 -8 66 248
use NAND3X1  _8461_
timestamp 0
transform -1 0 2550 0 1 9850
box -6 -8 106 248
use OAI21X1  _8462_
timestamp 0
transform -1 0 1990 0 -1 10810
box -6 -8 106 248
use OR2X2  _8463_
timestamp 0
transform 1 0 2610 0 -1 10810
box -6 -8 106 248
use NOR2X1  _8464_
timestamp 0
transform 1 0 2030 0 -1 10810
box -6 -8 86 248
use OAI21X1  _8465_
timestamp 0
transform 1 0 2470 0 -1 10810
box -6 -8 106 248
use NAND3X1  _8466_
timestamp 0
transform -1 0 3230 0 -1 10810
box -6 -8 106 248
use OR2X2  _8467_
timestamp 0
transform 1 0 2170 0 -1 10810
box -6 -8 106 248
use OAI21X1  _8468_
timestamp 0
transform -1 0 2410 0 -1 10810
box -6 -8 106 248
use NAND3X1  _8469_
timestamp 0
transform 1 0 2990 0 -1 10810
box -6 -8 106 248
use NAND2X1  _8470_
timestamp 0
transform 1 0 3450 0 -1 10810
box -6 -8 86 248
use OR2X2  _8471_
timestamp 0
transform 1 0 4250 0 -1 10810
box -6 -8 106 248
use NAND2X1  _8472_
timestamp 0
transform -1 0 4210 0 -1 10810
box -6 -8 86 248
use NAND2X1  _8473_
timestamp 0
transform 1 0 4190 0 1 10330
box -6 -8 86 248
use AOI22X1  _8474_
timestamp 0
transform -1 0 4410 0 -1 8410
box -6 -8 126 248
use INVX1  _8475_
timestamp 0
transform 1 0 4550 0 1 10810
box -6 -8 66 248
use OAI21X1  _8476_
timestamp 0
transform -1 0 4070 0 -1 10810
box -6 -8 106 248
use NAND2X1  _8477_
timestamp 0
transform -1 0 2410 0 1 10810
box -6 -8 86 248
use NOR2X1  _8478_
timestamp 0
transform -1 0 1290 0 -1 8890
box -6 -8 86 248
use AOI21X1  _8479_
timestamp 0
transform 1 0 1310 0 1 8890
box -6 -8 106 248
use NAND2X1  _8480_
timestamp 0
transform -1 0 1390 0 1 9850
box -6 -8 86 248
use OAI21X1  _8481_
timestamp 0
transform -1 0 1550 0 1 9850
box -6 -8 106 248
use INVX1  _8482_
timestamp 0
transform 1 0 1950 0 1 10810
box -6 -8 66 248
use NAND3X1  _8483_
timestamp 0
transform 1 0 2450 0 1 10810
box -6 -8 106 248
use NOR2X1  _8484_
timestamp 0
transform 1 0 1930 0 -1 10330
box -6 -8 86 248
use NAND3X1  _8485_
timestamp 0
transform -1 0 1870 0 -1 10330
box -6 -8 106 248
use OAI21X1  _8486_
timestamp 0
transform -1 0 1690 0 1 10810
box -6 -8 106 248
use NAND2X1  _8487_
timestamp 0
transform -1 0 1530 0 1 10810
box -6 -8 86 248
use AOI21X1  _8488_
timestamp 0
transform 1 0 2730 0 1 10810
box -6 -8 106 248
use INVX1  _8489_
timestamp 0
transform 1 0 3470 0 1 10810
box -6 -8 66 248
use NAND3X1  _8490_
timestamp 0
transform -1 0 2690 0 1 10810
box -6 -8 106 248
use NAND2X1  _8491_
timestamp 0
transform 1 0 3590 0 1 10810
box -6 -8 86 248
use NOR2X1  _8492_
timestamp 0
transform -1 0 4070 0 1 10810
box -6 -8 86 248
use AND2X2  _8493_
timestamp 0
transform 1 0 4130 0 1 10810
box -6 -8 106 248
use OAI21X1  _8494_
timestamp 0
transform 1 0 4270 0 1 10810
box -6 -8 106 248
use OAI21X1  _8495_
timestamp 0
transform -1 0 4510 0 1 10810
box -6 -8 106 248
use INVX1  _8496_
timestamp 0
transform -1 0 4310 0 1 7930
box -6 -8 66 248
use NAND3X1  _8497_
timestamp 0
transform -1 0 2150 0 1 10810
box -6 -8 106 248
use AOI21X1  _8498_
timestamp 0
transform 1 0 1350 0 -1 8890
box -6 -8 106 248
use NAND2X1  _8499_
timestamp 0
transform -1 0 1530 0 -1 9370
box -6 -8 86 248
use OAI21X1  _8500_
timestamp 0
transform -1 0 1590 0 -1 10330
box -6 -8 106 248
use NAND3X1  _8501_
timestamp 0
transform 1 0 2250 0 -1 11290
box -6 -8 106 248
use NOR3X1  _8502_
timestamp 0
transform -1 0 1910 0 1 10810
box -6 -8 186 248
use INVX1  _8503_
timestamp 0
transform -1 0 1650 0 -1 11290
box -6 -8 66 248
use OAI21X1  _8504_
timestamp 0
transform 1 0 2090 0 -1 11290
box -6 -8 106 248
use NAND2X1  _8505_
timestamp 0
transform -1 0 2490 0 -1 11290
box -6 -8 86 248
use NAND2X1  _8506_
timestamp 0
transform -1 0 2750 0 -1 11290
box -6 -8 86 248
use NAND3X1  _8507_
timestamp 0
transform 1 0 2530 0 -1 11290
box -6 -8 106 248
use NAND2X1  _8508_
timestamp 0
transform -1 0 3150 0 -1 11290
box -6 -8 86 248
use AOI21X1  _8509_
timestamp 0
transform 1 0 2850 0 -1 10810
box -6 -8 106 248
use NOR2X1  _8510_
timestamp 0
transform -1 0 2970 0 1 10810
box -6 -8 86 248
use OAI21X1  _8511_
timestamp 0
transform -1 0 3950 0 1 10810
box -6 -8 106 248
use NAND2X1  _8512_
timestamp 0
transform 1 0 3730 0 1 10810
box -6 -8 86 248
use NOR2X1  _8513_
timestamp 0
transform 1 0 3450 0 -1 11290
box -6 -8 86 248
use AND2X2  _8514_
timestamp 0
transform 1 0 3190 0 -1 11290
box -6 -8 106 248
use AND2X2  _8515_
timestamp 0
transform 1 0 3290 0 -1 10810
box -6 -8 106 248
use NAND3X1  _8516_
timestamp 0
transform -1 0 3410 0 1 10810
box -6 -8 106 248
use AOI21X1  _8517_
timestamp 0
transform 1 0 3030 0 1 10810
box -6 -8 106 248
use OAI21X1  _8518_
timestamp 0
transform -1 0 3270 0 1 10810
box -6 -8 106 248
use NOR2X1  _8519_
timestamp 0
transform 1 0 3330 0 -1 11290
box -6 -8 86 248
use OAI21X1  _8520_
timestamp 0
transform 1 0 3590 0 -1 11290
box -6 -8 106 248
use NAND2X1  _8521_
timestamp 0
transform -1 0 4030 0 1 9850
box -6 -8 86 248
use OAI21X1  _8522_
timestamp 0
transform -1 0 4190 0 1 7930
box -6 -8 106 248
use INVX1  _8523_
timestamp 0
transform -1 0 4450 0 -1 11290
box -6 -8 66 248
use INVX1  _8524_
timestamp 0
transform -1 0 2850 0 1 11290
box -6 -8 66 248
use NAND2X1  _8525_
timestamp 0
transform 1 0 1830 0 -1 11290
box -6 -8 86 248
use NOR2X1  _8526_
timestamp 0
transform -1 0 1190 0 1 8410
box -6 -8 86 248
use INVX1  _8527_
timestamp 0
transform 1 0 1250 0 1 8410
box -6 -8 66 248
use OAI21X1  _8528_
timestamp 0
transform 1 0 1190 0 -1 9370
box -6 -8 106 248
use NAND3X1  _8529_
timestamp 0
transform 1 0 1250 0 1 11290
box -6 -8 106 248
use INVX1  _8530_
timestamp 0
transform 1 0 1130 0 1 11290
box -6 -8 66 248
use OAI21X1  _8531_
timestamp 0
transform -1 0 2050 0 -1 11290
box -6 -8 106 248
use NAND2X1  _8532_
timestamp 0
transform -1 0 1610 0 1 11290
box -6 -8 86 248
use NAND3X1  _8533_
timestamp 0
transform 1 0 1650 0 1 11290
box -6 -8 106 248
use NAND3X1  _8534_
timestamp 0
transform 1 0 1810 0 1 11290
box -6 -8 106 248
use NAND2X1  _8535_
timestamp 0
transform 1 0 1390 0 1 11290
box -6 -8 86 248
use NAND3X1  _8536_
timestamp 0
transform -1 0 2070 0 1 11290
box -6 -8 106 248
use NAND2X1  _8537_
timestamp 0
transform -1 0 2190 0 1 11290
box -6 -8 86 248
use OAI21X1  _8538_
timestamp 0
transform -1 0 2990 0 1 11290
box -6 -8 106 248
use NOR2X1  _8539_
timestamp 0
transform 1 0 3050 0 1 11290
box -6 -8 86 248
use INVX1  _8540_
timestamp 0
transform 1 0 3730 0 -1 11290
box -6 -8 66 248
use AOI21X1  _8541_
timestamp 0
transform 1 0 3850 0 -1 11290
box -6 -8 106 248
use AOI22X1  _8542_
timestamp 0
transform -1 0 4110 0 -1 11290
box -6 -8 126 248
use OAI21X1  _8543_
timestamp 0
transform -1 0 2350 0 1 11290
box -6 -8 106 248
use NOR2X1  _8544_
timestamp 0
transform -1 0 3010 0 -1 11290
box -6 -8 86 248
use AOI21X1  _8545_
timestamp 0
transform -1 0 2890 0 -1 11290
box -6 -8 106 248
use INVX1  _8546_
timestamp 0
transform -1 0 2230 0 -1 8410
box -6 -8 66 248
use NAND3X1  _8547_
timestamp 0
transform 1 0 1690 0 -1 11290
box -6 -8 106 248
use INVX1  _8548_
timestamp 0
transform -1 0 1710 0 -1 8890
box -6 -8 66 248
use OAI21X1  _8549_
timestamp 0
transform -1 0 1590 0 -1 8890
box -6 -8 106 248
use INVX1  _8550_
timestamp 0
transform -1 0 1710 0 1 8410
box -6 -8 66 248
use NAND3X1  _8551_
timestamp 0
transform 1 0 1730 0 -1 8410
box -6 -8 106 248
use OAI21X1  _8552_
timestamp 0
transform 1 0 1430 0 -1 11290
box -6 -8 106 248
use NAND2X1  _8553_
timestamp 0
transform 1 0 1890 0 -1 8410
box -6 -8 86 248
use AOI21X1  _8554_
timestamp 0
transform 1 0 2010 0 -1 8410
box -6 -8 106 248
use NAND3X1  _8555_
timestamp 0
transform 1 0 1770 0 -1 8890
box -6 -8 106 248
use NAND2X1  _8556_
timestamp 0
transform 1 0 1750 0 1 8410
box -6 -8 86 248
use AOI21X1  _8557_
timestamp 0
transform 1 0 1870 0 1 8410
box -6 -8 106 248
use OAI21X1  _8558_
timestamp 0
transform 1 0 2050 0 1 6970
box -6 -8 106 248
use INVX1  _8559_
timestamp 0
transform 1 0 2190 0 1 6970
box -6 -8 66 248
use OR2X2  _8560_
timestamp 0
transform 1 0 1890 0 1 6970
box -6 -8 106 248
use OAI21X1  _8561_
timestamp 0
transform 1 0 2550 0 1 6970
box -6 -8 106 248
use OAI22X1  _8562_
timestamp 0
transform -1 0 2810 0 1 6970
box -6 -8 126 248
use NAND2X1  _8563_
timestamp 0
transform 1 0 3050 0 -1 7450
box -6 -8 86 248
use NOR2X1  _8564_
timestamp 0
transform 1 0 2430 0 1 6970
box -6 -8 86 248
use NOR2X1  _8565_
timestamp 0
transform 1 0 2310 0 1 6970
box -6 -8 86 248
use OAI21X1  _8566_
timestamp 0
transform -1 0 1610 0 1 8410
box -6 -8 106 248
use INVX1  _8567_
timestamp 0
transform 1 0 1730 0 -1 7930
box -6 -8 66 248
use OAI21X1  _8568_
timestamp 0
transform -1 0 1850 0 1 7930
box -6 -8 106 248
use NAND2X1  _8569_
timestamp 0
transform -1 0 1910 0 -1 7930
box -6 -8 86 248
use OR2X2  _8570_
timestamp 0
transform 1 0 1970 0 -1 7930
box -6 -8 106 248
use NAND3X1  _8571_
timestamp 0
transform 1 0 2250 0 -1 7930
box -6 -8 106 248
use NAND2X1  _8572_
timestamp 0
transform 1 0 2130 0 -1 7930
box -6 -8 86 248
use NAND2X1  _8573_
timestamp 0
transform -1 0 1810 0 1 7450
box -6 -8 86 248
use NAND2X1  _8574_
timestamp 0
transform -1 0 2310 0 -1 7450
box -6 -8 86 248
use AND2X2  _8575_
timestamp 0
transform 1 0 2350 0 -1 7450
box -6 -8 106 248
use OAI21X1  _8576_
timestamp 0
transform 1 0 2490 0 -1 7450
box -6 -8 106 248
use OAI21X1  _8577_
timestamp 0
transform 1 0 2650 0 -1 7450
box -6 -8 106 248
use INVX1  _8578_
timestamp 0
transform -1 0 4070 0 1 6970
box -6 -8 66 248
use INVX1  _8579_
timestamp 0
transform -1 0 2170 0 -1 7450
box -6 -8 66 248
use AOI21X1  _8580_
timestamp 0
transform -1 0 1910 0 -1 7450
box -6 -8 106 248
use NOR2X1  _8581_
timestamp 0
transform -1 0 1930 0 1 7450
box -6 -8 86 248
use NAND3X1  _8582_
timestamp 0
transform -1 0 2090 0 1 7450
box -6 -8 106 248
use OAI21X1  _8583_
timestamp 0
transform -1 0 2050 0 -1 7450
box -6 -8 106 248
use OAI21X1  _8584_
timestamp 0
transform -1 0 1470 0 1 8410
box -6 -8 106 248
use INVX1  _8585_
timestamp 0
transform -1 0 1370 0 -1 8410
box -6 -8 66 248
use OR2X2  _8586_
timestamp 0
transform -1 0 1710 0 1 7930
box -6 -8 106 248
use OAI21X1  _8587_
timestamp 0
transform -1 0 1670 0 -1 7930
box -6 -8 106 248
use NAND2X1  _8588_
timestamp 0
transform 1 0 1330 0 1 6970
box -6 -8 86 248
use OR2X2  _8589_
timestamp 0
transform 1 0 1610 0 1 6970
box -6 -8 106 248
use NAND3X1  _8590_
timestamp 0
transform 1 0 1450 0 1 6970
box -6 -8 106 248
use AND2X2  _8591_
timestamp 0
transform -1 0 1170 0 1 6970
box -6 -8 106 248
use NOR2X1  _8592_
timestamp 0
transform 1 0 1210 0 1 6970
box -6 -8 86 248
use OAI21X1  _8593_
timestamp 0
transform 1 0 1230 0 -1 6970
box -6 -8 106 248
use NAND2X1  _8594_
timestamp 0
transform 1 0 1370 0 -1 6970
box -6 -8 86 248
use AND2X2  _8595_
timestamp 0
transform 1 0 1750 0 -1 6970
box -6 -8 106 248
use NOR2X1  _8596_
timestamp 0
transform 1 0 1910 0 -1 6970
box -6 -8 86 248
use NOR2X1  _8597_
timestamp 0
transform 1 0 2030 0 -1 6970
box -6 -8 86 248
use AOI22X1  _8598_
timestamp 0
transform -1 0 3830 0 -1 6970
box -6 -8 126 248
use NAND2X1  _8599_
timestamp 0
transform 1 0 2830 0 -1 6970
box -6 -8 86 248
use INVX1  _8600_
timestamp 0
transform 1 0 1490 0 -1 6970
box -6 -8 66 248
use AOI21X1  _8601_
timestamp 0
transform -1 0 1710 0 -1 6970
box -6 -8 106 248
use NAND2X1  _8602_
timestamp 0
transform 1 0 570 0 1 6970
box -6 -8 86 248
use NOR2X1  _8603_
timestamp 0
transform 1 0 450 0 1 6970
box -6 -8 86 248
use AOI21X1  _8604_
timestamp 0
transform -1 0 390 0 1 6970
box -6 -8 106 248
use NOR2X1  _8605_
timestamp 0
transform 1 0 310 0 -1 6970
box -6 -8 86 248
use AND2X2  _8606_
timestamp 0
transform 1 0 2150 0 -1 6970
box -6 -8 106 248
use OAI21X1  _8607_
timestamp 0
transform 1 0 2290 0 -1 6970
box -6 -8 106 248
use OAI21X1  _8608_
timestamp 0
transform 1 0 2450 0 -1 6970
box -6 -8 106 248
use OAI21X1  _8609_
timestamp 0
transform 1 0 5990 0 -1 9850
box -6 -8 106 248
use OAI21X1  _8610_
timestamp 0
transform -1 0 6150 0 1 9850
box -6 -8 106 248
use INVX1  _8611_
timestamp 0
transform -1 0 5690 0 -1 9850
box -6 -8 66 248
use NOR2X1  _8612_
timestamp 0
transform 1 0 5870 0 -1 9850
box -6 -8 86 248
use NAND2X1  _8613_
timestamp 0
transform 1 0 5750 0 -1 9850
box -6 -8 86 248
use NAND2X1  _8614_
timestamp 0
transform 1 0 5710 0 1 9370
box -6 -8 86 248
use NAND2X1  _8615_
timestamp 0
transform -1 0 4710 0 -1 7450
box -6 -8 86 248
use OAI21X1  _8616_
timestamp 0
transform -1 0 4850 0 -1 7450
box -6 -8 106 248
use NAND2X1  _8617_
timestamp 0
transform 1 0 6650 0 -1 8410
box -6 -8 86 248
use INVX1  _8618_
timestamp 0
transform 1 0 6470 0 1 9370
box -6 -8 66 248
use NOR2X1  _8619_
timestamp 0
transform 1 0 6810 0 1 10330
box -6 -8 86 248
use AOI21X1  _8620_
timestamp 0
transform 1 0 6670 0 1 10330
box -6 -8 106 248
use NOR2X1  _8621_
timestamp 0
transform 1 0 6350 0 1 9850
box -6 -8 86 248
use OAI21X1  _8622_
timestamp 0
transform 1 0 6210 0 1 9850
box -6 -8 106 248
use AND2X2  _8623_
timestamp 0
transform 1 0 6430 0 -1 9850
box -6 -8 106 248
use OR2X2  _8624_
timestamp 0
transform -1 0 6250 0 -1 9850
box -6 -8 106 248
use OR2X2  _8625_
timestamp 0
transform 1 0 6190 0 1 9370
box -6 -8 106 248
use OAI21X1  _8626_
timestamp 0
transform -1 0 6390 0 -1 9850
box -6 -8 106 248
use NAND2X1  _8627_
timestamp 0
transform 1 0 6350 0 1 9370
box -6 -8 86 248
use NOR2X1  _8628_
timestamp 0
transform -1 0 6470 0 -1 9370
box -6 -8 86 248
use NAND2X1  _8629_
timestamp 0
transform 1 0 6270 0 -1 9370
box -6 -8 86 248
use NAND2X1  _8630_
timestamp 0
transform 1 0 6990 0 1 8410
box -6 -8 86 248
use OAI21X1  _8631_
timestamp 0
transform -1 0 6950 0 1 8410
box -6 -8 106 248
use INVX1  _8632_
timestamp 0
transform -1 0 6150 0 1 9370
box -6 -8 66 248
use OAI21X1  _8633_
timestamp 0
transform 1 0 6110 0 -1 9370
box -6 -8 106 248
use OAI21X1  _8634_
timestamp 0
transform 1 0 5290 0 1 9370
box -6 -8 106 248
use OAI21X1  _8635_
timestamp 0
transform -1 0 5670 0 -1 9370
box -6 -8 106 248
use MUX2X1  _8636_
timestamp 0
transform 1 0 5410 0 -1 9370
box -6 -8 126 248
use NAND2X1  _8637_
timestamp 0
transform 1 0 5110 0 1 8890
box -6 -8 86 248
use OR2X2  _8638_
timestamp 0
transform -1 0 5150 0 -1 8890
box -6 -8 106 248
use NAND2X1  _8639_
timestamp 0
transform -1 0 5290 0 -1 8890
box -6 -8 86 248
use INVX1  _8640_
timestamp 0
transform 1 0 6090 0 -1 8890
box -6 -8 66 248
use NOR2X1  _8641_
timestamp 0
transform -1 0 6690 0 1 8410
box -6 -8 86 248
use NAND2X1  _8642_
timestamp 0
transform 1 0 6730 0 1 8410
box -6 -8 86 248
use NAND2X1  _8643_
timestamp 0
transform -1 0 6830 0 1 7930
box -6 -8 86 248
use OAI22X1  _8644_
timestamp 0
transform 1 0 6590 0 1 7930
box -6 -8 126 248
use NOR2X1  _8645_
timestamp 0
transform 1 0 6110 0 1 7930
box -6 -8 86 248
use NAND2X1  _8646_
timestamp 0
transform 1 0 6470 0 1 8410
box -6 -8 86 248
use INVX1  _8647_
timestamp 0
transform -1 0 6350 0 -1 8410
box -6 -8 66 248
use INVX1  _8648_
timestamp 0
transform 1 0 5830 0 1 8410
box -6 -8 66 248
use NOR2X1  _8649_
timestamp 0
transform 1 0 5710 0 -1 9370
box -6 -8 86 248
use OAI21X1  _8650_
timestamp 0
transform -1 0 5590 0 1 8890
box -6 -8 106 248
use OAI21X1  _8651_
timestamp 0
transform 1 0 6090 0 -1 7930
box -6 -8 106 248
use OAI21X1  _8652_
timestamp 0
transform 1 0 5370 0 1 8410
box -6 -8 106 248
use NOR2X1  _8653_
timestamp 0
transform 1 0 6070 0 1 8410
box -6 -8 86 248
use NAND2X1  _8654_
timestamp 0
transform -1 0 6010 0 1 8410
box -6 -8 86 248
use INVX1  _8655_
timestamp 0
transform -1 0 6270 0 1 8410
box -6 -8 66 248
use NOR2X1  _8656_
timestamp 0
transform 1 0 6170 0 -1 8410
box -6 -8 86 248
use OAI21X1  _8657_
timestamp 0
transform 1 0 6030 0 -1 8410
box -6 -8 106 248
use AOI21X1  _8658_
timestamp 0
transform -1 0 5990 0 -1 8410
box -6 -8 106 248
use NOR2X1  _8659_
timestamp 0
transform -1 0 6070 0 1 7930
box -6 -8 86 248
use NAND2X1  _8660_
timestamp 0
transform -1 0 7350 0 1 7930
box -6 -8 86 248
use INVX1  _8661_
timestamp 0
transform 1 0 7150 0 1 9850
box -6 -8 66 248
use AOI21X1  _8662_
timestamp 0
transform 1 0 6470 0 1 9850
box -6 -8 106 248
use OAI21X1  _8663_
timestamp 0
transform 1 0 6630 0 1 9850
box -6 -8 106 248
use OAI21X1  _8664_
timestamp 0
transform 1 0 6770 0 1 9850
box -6 -8 106 248
use OR2X2  _8665_
timestamp 0
transform 1 0 6990 0 -1 9850
box -6 -8 106 248
use NAND2X1  _8666_
timestamp 0
transform 1 0 6850 0 -1 9850
box -6 -8 86 248
use NAND2X1  _8667_
timestamp 0
transform -1 0 6890 0 1 9370
box -6 -8 86 248
use AOI21X1  _8668_
timestamp 0
transform 1 0 6310 0 1 8410
box -6 -8 106 248
use AND2X2  _8669_
timestamp 0
transform 1 0 7350 0 -1 8410
box -6 -8 106 248
use OAI21X1  _8670_
timestamp 0
transform 1 0 7210 0 -1 8410
box -6 -8 106 248
use OAI21X1  _8671_
timestamp 0
transform 1 0 7390 0 1 7930
box -6 -8 106 248
use OAI21X1  _8672_
timestamp 0
transform 1 0 7390 0 1 8410
box -6 -8 106 248
use INVX1  _8673_
timestamp 0
transform 1 0 7430 0 1 10330
box -6 -8 66 248
use OAI21X1  _8674_
timestamp 0
transform 1 0 5890 0 -1 10330
box -6 -8 106 248
use OAI21X1  _8675_
timestamp 0
transform -1 0 6370 0 1 10330
box -6 -8 106 248
use OR2X2  _8676_
timestamp 0
transform -1 0 6210 0 1 10330
box -6 -8 106 248
use NAND2X1  _8677_
timestamp 0
transform 1 0 6150 0 -1 10330
box -6 -8 86 248
use OR2X2  _8678_
timestamp 0
transform 1 0 7470 0 -1 10330
box -6 -8 106 248
use NAND2X1  _8679_
timestamp 0
transform -1 0 7430 0 -1 10330
box -6 -8 86 248
use NAND2X1  _8680_
timestamp 0
transform -1 0 7330 0 1 9850
box -6 -8 86 248
use INVX1  _8681_
timestamp 0
transform 1 0 7290 0 -1 9850
box -6 -8 66 248
use NOR2X1  _8682_
timestamp 0
transform 1 0 6790 0 -1 8410
box -6 -8 86 248
use NAND2X1  _8683_
timestamp 0
transform 1 0 7490 0 -1 8410
box -6 -8 86 248
use NAND2X1  _8684_
timestamp 0
transform -1 0 7670 0 -1 7930
box -6 -8 86 248
use OAI22X1  _8685_
timestamp 0
transform 1 0 6610 0 1 7450
box -6 -8 126 248
use NAND2X1  _8686_
timestamp 0
transform -1 0 7010 0 -1 8410
box -6 -8 86 248
use INVX1  _8687_
timestamp 0
transform -1 0 6730 0 -1 8890
box -6 -8 66 248
use NAND2X1  _8688_
timestamp 0
transform -1 0 6850 0 -1 8890
box -6 -8 86 248
use OAI21X1  _8689_
timestamp 0
transform 1 0 7150 0 -1 9850
box -6 -8 106 248
use INVX1  _8690_
timestamp 0
transform 1 0 6830 0 -1 9370
box -6 -8 66 248
use OAI21X1  _8691_
timestamp 0
transform 1 0 6890 0 1 8890
box -6 -8 106 248
use OAI21X1  _8692_
timestamp 0
transform -1 0 5330 0 1 8890
box -6 -8 106 248
use NOR2X1  _8693_
timestamp 0
transform 1 0 5630 0 1 8890
box -6 -8 86 248
use NAND2X1  _8694_
timestamp 0
transform -1 0 5990 0 1 8890
box -6 -8 86 248
use OAI21X1  _8695_
timestamp 0
transform 1 0 5750 0 1 8890
box -6 -8 106 248
use NAND2X1  _8696_
timestamp 0
transform 1 0 6050 0 1 8890
box -6 -8 86 248
use NAND2X1  _8697_
timestamp 0
transform 1 0 6190 0 -1 8890
box -6 -8 86 248
use OR2X2  _8698_
timestamp 0
transform 1 0 6190 0 1 8890
box -6 -8 106 248
use NAND2X1  _8699_
timestamp 0
transform -1 0 6410 0 1 8890
box -6 -8 86 248
use INVX1  _8700_
timestamp 0
transform -1 0 6370 0 -1 8890
box -6 -8 66 248
use NOR2X1  _8701_
timestamp 0
transform 1 0 6430 0 -1 8890
box -6 -8 86 248
use NAND2X1  _8702_
timestamp 0
transform 1 0 6550 0 -1 8890
box -6 -8 86 248
use NAND2X1  _8703_
timestamp 0
transform 1 0 7130 0 1 8410
box -6 -8 86 248
use OAI21X1  _8704_
timestamp 0
transform -1 0 7150 0 -1 8410
box -6 -8 106 248
use INVX1  _8705_
timestamp 0
transform 1 0 6230 0 -1 7450
box -6 -8 66 248
use NAND2X1  _8706_
timestamp 0
transform 1 0 7250 0 1 8410
box -6 -8 86 248
use INVX1  _8707_
timestamp 0
transform -1 0 6610 0 -1 10330
box -6 -8 66 248
use NAND2X1  _8708_
timestamp 0
transform 1 0 6670 0 -1 10330
box -6 -8 86 248
use OR2X2  _8709_
timestamp 0
transform 1 0 6790 0 -1 10330
box -6 -8 106 248
use NAND2X1  _8710_
timestamp 0
transform 1 0 6950 0 -1 10330
box -6 -8 86 248
use NOR2X1  _8711_
timestamp 0
transform 1 0 7070 0 -1 10330
box -6 -8 86 248
use INVX1  _8712_
timestamp 0
transform -1 0 6750 0 1 9370
box -6 -8 66 248
use NAND2X1  _8713_
timestamp 0
transform 1 0 7210 0 -1 10330
box -6 -8 86 248
use NAND2X1  _8714_
timestamp 0
transform -1 0 6650 0 1 9370
box -6 -8 86 248
use OR2X2  _8715_
timestamp 0
transform 1 0 7430 0 -1 7930
box -6 -8 106 248
use AOI21X1  _8716_
timestamp 0
transform -1 0 7370 0 -1 7930
box -6 -8 106 248
use AOI22X1  _8717_
timestamp 0
transform 1 0 6450 0 1 7450
box -6 -8 126 248
use NAND2X1  _8718_
timestamp 0
transform 1 0 6050 0 1 7450
box -6 -8 86 248
use NOR2X1  _8719_
timestamp 0
transform -1 0 6550 0 -1 7930
box -6 -8 86 248
use INVX1  _8720_
timestamp 0
transform 1 0 6610 0 -1 7930
box -6 -8 66 248
use NAND3X1  _8721_
timestamp 0
transform 1 0 5530 0 1 7450
box -6 -8 106 248
use INVX1  _8722_
timestamp 0
transform 1 0 5730 0 -1 7450
box -6 -8 66 248
use AOI21X1  _8723_
timestamp 0
transform -1 0 5490 0 1 7450
box -6 -8 106 248
use NOR2X1  _8724_
timestamp 0
transform 1 0 5430 0 -1 7450
box -6 -8 86 248
use OAI21X1  _8725_
timestamp 0
transform 1 0 6530 0 -1 9370
box -6 -8 106 248
use NOR2X1  _8726_
timestamp 0
transform -1 0 6530 0 1 8890
box -6 -8 86 248
use AOI21X1  _8727_
timestamp 0
transform -1 0 6790 0 -1 9370
box -6 -8 106 248
use NAND3X1  _8728_
timestamp 0
transform -1 0 6830 0 1 8890
box -6 -8 106 248
use OAI21X1  _8729_
timestamp 0
transform -1 0 6690 0 1 8890
box -6 -8 106 248
use NOR2X1  _8730_
timestamp 0
transform 1 0 5970 0 -1 7450
box -6 -8 86 248
use NAND2X1  _8731_
timestamp 0
transform -1 0 6170 0 -1 7450
box -6 -8 86 248
use NAND2X1  _8732_
timestamp 0
transform -1 0 6270 0 1 7450
box -6 -8 86 248
use OAI21X1  _8733_
timestamp 0
transform -1 0 6010 0 1 7450
box -6 -8 106 248
use AOI21X1  _8734_
timestamp 0
transform -1 0 5670 0 -1 7450
box -6 -8 106 248
use OR2X2  _8735_
timestamp 0
transform 1 0 5830 0 -1 7450
box -6 -8 106 248
use NAND2X1  _8736_
timestamp 0
transform 1 0 6050 0 1 6970
box -6 -8 86 248
use NAND2X1  _8737_
timestamp 0
transform 1 0 5910 0 1 6970
box -6 -8 86 248
use AND2X2  _8738_
timestamp 0
transform 1 0 5590 0 -1 6970
box -6 -8 106 248
use OAI21X1  _8739_
timestamp 0
transform -1 0 5550 0 -1 6970
box -6 -8 106 248
use OAI22X1  _8740_
timestamp 0
transform 1 0 5410 0 1 6490
box -6 -8 126 248
use NAND2X1  _8741_
timestamp 0
transform -1 0 4930 0 1 6490
box -6 -8 86 248
use OAI21X1  _8742_
timestamp 0
transform 1 0 5770 0 1 6970
box -6 -8 106 248
use NAND3X1  _8743_
timestamp 0
transform 1 0 6170 0 1 6970
box -6 -8 106 248
use INVX1  _8744_
timestamp 0
transform -1 0 6390 0 1 6970
box -6 -8 66 248
use AOI21X1  _8745_
timestamp 0
transform -1 0 5390 0 -1 6970
box -6 -8 106 248
use INVX1  _8746_
timestamp 0
transform 1 0 5290 0 1 6970
box -6 -8 66 248
use NAND2X1  _8747_
timestamp 0
transform -1 0 4990 0 -1 6970
box -6 -8 86 248
use NAND2X1  _8748_
timestamp 0
transform 1 0 5410 0 1 6970
box -6 -8 86 248
use NAND2X1  _8749_
timestamp 0
transform 1 0 5030 0 -1 6970
box -6 -8 86 248
use AND2X2  _8750_
timestamp 0
transform -1 0 5210 0 1 6490
box -6 -8 106 248
use OAI21X1  _8751_
timestamp 0
transform 1 0 5270 0 1 6490
box -6 -8 106 248
use OAI21X1  _8752_
timestamp 0
transform -1 0 5070 0 1 6490
box -6 -8 106 248
use NAND2X1  _8753_
timestamp 0
transform 1 0 4330 0 1 6490
box -6 -8 86 248
use OAI21X1  _8754_
timestamp 0
transform -1 0 5250 0 -1 6970
box -6 -8 106 248
use OAI21X1  _8755_
timestamp 0
transform -1 0 4790 0 1 6490
box -6 -8 106 248
use NAND2X1  _8756_
timestamp 0
transform 1 0 4110 0 -1 7450
box -6 -8 86 248
use NAND2X1  _8757_
timestamp 0
transform 1 0 3930 0 1 7450
box -6 -8 86 248
use NOR2X1  _8758_
timestamp 0
transform -1 0 4150 0 1 7450
box -6 -8 86 248
use NAND2X1  _8759_
timestamp 0
transform -1 0 3030 0 -1 6970
box -6 -8 86 248
use OAI21X1  _8760_
timestamp 0
transform 1 0 1070 0 -1 6970
box -6 -8 106 248
use NAND2X1  _8761_
timestamp 0
transform -1 0 1830 0 1 6970
box -6 -8 86 248
use OAI21X1  _8762_
timestamp 0
transform 1 0 910 0 1 6970
box -6 -8 106 248
use INVX1  _8763_
timestamp 0
transform 1 0 4310 0 1 8410
box -6 -8 66 248
use OR2X2  _8764_
timestamp 0
transform -1 0 5330 0 1 8410
box -6 -8 106 248
use OAI21X1  _8765_
timestamp 0
transform -1 0 4110 0 1 8410
box -6 -8 106 248
use OAI21X1  _8766_
timestamp 0
transform -1 0 4250 0 1 8410
box -6 -8 106 248
use INVX1  _8767_
timestamp 0
transform -1 0 5050 0 -1 9370
box -6 -8 66 248
use OAI21X1  _8768_
timestamp 0
transform -1 0 5190 0 1 8410
box -6 -8 106 248
use OAI21X1  _8769_
timestamp 0
transform 1 0 4950 0 1 8410
box -6 -8 106 248
use NAND2X1  _8770_
timestamp 0
transform 1 0 5250 0 -1 8410
box -6 -8 86 248
use NAND2X1  _8771_
timestamp 0
transform -1 0 3510 0 -1 8890
box -6 -8 86 248
use OAI21X1  _8772_
timestamp 0
transform -1 0 3670 0 -1 8890
box -6 -8 106 248
use NAND2X1  _8773_
timestamp 0
transform -1 0 4850 0 1 9370
box -6 -8 86 248
use OAI21X1  _8774_
timestamp 0
transform -1 0 4990 0 1 9370
box -6 -8 106 248
use AND2X2  _8775_
timestamp 0
transform 1 0 5390 0 -1 8410
box -6 -8 106 248
use NAND2X1  _8776_
timestamp 0
transform -1 0 3870 0 1 8890
box -6 -8 86 248
use OAI21X1  _8777_
timestamp 0
transform 1 0 3830 0 -1 10810
box -6 -8 106 248
use NAND2X1  _8778_
timestamp 0
transform -1 0 2850 0 1 9370
box -6 -8 86 248
use OAI21X1  _8779_
timestamp 0
transform -1 0 2910 0 -1 9850
box -6 -8 106 248
use OAI21X1  _8780_
timestamp 0
transform -1 0 4050 0 -1 8890
box -6 -8 106 248
use OAI21X1  _8781_
timestamp 0
transform 1 0 3810 0 -1 8890
box -6 -8 106 248
use OAI21X1  _8782_
timestamp 0
transform -1 0 5350 0 -1 9370
box -6 -8 106 248
use OAI21X1  _8783_
timestamp 0
transform 1 0 5090 0 -1 9370
box -6 -8 106 248
use NAND2X1  _8784_
timestamp 0
transform 1 0 3310 0 -1 8890
box -6 -8 86 248
use OAI21X1  _8785_
timestamp 0
transform 1 0 3150 0 -1 8890
box -6 -8 106 248
use NAND2X1  _8786_
timestamp 0
transform 1 0 3150 0 -1 9370
box -6 -8 86 248
use OAI21X1  _8787_
timestamp 0
transform 1 0 3010 0 -1 9370
box -6 -8 106 248
use NAND2X1  _8788_
timestamp 0
transform -1 0 1770 0 -1 7450
box -6 -8 86 248
use OAI21X1  _8789_
timestamp 0
transform 1 0 1170 0 -1 7450
box -6 -8 106 248
use NAND2X1  _8790_
timestamp 0
transform -1 0 1550 0 1 7450
box -6 -8 86 248
use OAI21X1  _8791_
timestamp 0
transform 1 0 1330 0 1 7450
box -6 -8 106 248
use INVX1  _8792_
timestamp 0
transform 1 0 5650 0 1 10330
box -6 -8 66 248
use OAI21X1  _8793_
timestamp 0
transform -1 0 4510 0 1 8410
box -6 -8 106 248
use OAI21X1  _8794_
timestamp 0
transform -1 0 4910 0 1 8410
box -6 -8 106 248
use INVX1  _8795_
timestamp 0
transform 1 0 3690 0 1 8890
box -6 -8 66 248
use OAI21X1  _8796_
timestamp 0
transform -1 0 3950 0 1 8410
box -6 -8 106 248
use OAI21X1  _8797_
timestamp 0
transform 1 0 3690 0 1 8410
box -6 -8 106 248
use NAND2X1  _8798_
timestamp 0
transform 1 0 5290 0 1 10810
box -6 -8 86 248
use OAI21X1  _8799_
timestamp 0
transform 1 0 5130 0 1 10810
box -6 -8 106 248
use NAND2X1  _8800_
timestamp 0
transform 1 0 3450 0 1 9370
box -6 -8 86 248
use OAI21X1  _8801_
timestamp 0
transform -1 0 3690 0 1 9370
box -6 -8 106 248
use NAND2X1  _8802_
timestamp 0
transform -1 0 2570 0 1 11770
box -6 -8 86 248
use OAI21X1  _8803_
timestamp 0
transform 1 0 2230 0 1 11770
box -6 -8 106 248
use NAND2X1  _8804_
timestamp 0
transform -1 0 1790 0 -1 11770
box -6 -8 86 248
use OAI21X1  _8805_
timestamp 0
transform 1 0 1570 0 -1 11770
box -6 -8 106 248
use OAI21X1  _8806_
timestamp 0
transform 1 0 4210 0 -1 9370
box -6 -8 106 248
use OAI21X1  _8807_
timestamp 0
transform -1 0 4690 0 -1 9370
box -6 -8 106 248
use OAI21X1  _8808_
timestamp 0
transform -1 0 4150 0 -1 9370
box -6 -8 106 248
use OAI21X1  _8809_
timestamp 0
transform 1 0 3890 0 -1 9370
box -6 -8 106 248
use NAND2X1  _8810_
timestamp 0
transform 1 0 5670 0 1 9850
box -6 -8 86 248
use OAI21X1  _8811_
timestamp 0
transform 1 0 5510 0 1 9850
box -6 -8 106 248
use NAND2X1  _8812_
timestamp 0
transform 1 0 5590 0 -1 10810
box -6 -8 86 248
use OAI21X1  _8813_
timestamp 0
transform 1 0 5450 0 -1 10810
box -6 -8 106 248
use NAND2X1  _8814_
timestamp 0
transform -1 0 4710 0 -1 6970
box -6 -8 86 248
use OAI21X1  _8815_
timestamp 0
transform -1 0 4870 0 -1 6970
box -6 -8 106 248
use NAND2X1  _8816_
timestamp 0
transform -1 0 5390 0 -1 7450
box -6 -8 86 248
use OAI21X1  _8817_
timestamp 0
transform 1 0 5170 0 -1 7450
box -6 -8 106 248
use INVX1  _8818_
timestamp 0
transform -1 0 5590 0 -1 8410
box -6 -8 66 248
use OAI21X1  _8819_
timestamp 0
transform 1 0 5530 0 -1 7930
box -6 -8 106 248
use OAI21X1  _8820_
timestamp 0
transform 1 0 5470 0 1 7930
box -6 -8 106 248
use INVX1  _8821_
timestamp 0
transform -1 0 6090 0 -1 10330
box -6 -8 66 248
use OAI21X1  _8822_
timestamp 0
transform 1 0 5690 0 -1 7930
box -6 -8 106 248
use OAI21X1  _8823_
timestamp 0
transform 1 0 5610 0 1 7930
box -6 -8 106 248
use NAND2X1  _8824_
timestamp 0
transform -1 0 5810 0 -1 8890
box -6 -8 86 248
use OAI21X1  _8825_
timestamp 0
transform 1 0 5350 0 -1 8890
box -6 -8 106 248
use NAND2X1  _8826_
timestamp 0
transform -1 0 6510 0 -1 10330
box -6 -8 86 248
use OAI21X1  _8827_
timestamp 0
transform 1 0 6290 0 -1 10330
box -6 -8 106 248
use NAND2X1  _8828_
timestamp 0
transform 1 0 6570 0 -1 9850
box -6 -8 86 248
use OAI21X1  _8829_
timestamp 0
transform -1 0 6810 0 -1 9850
box -6 -8 106 248
use NAND2X1  _8830_
timestamp 0
transform 1 0 6930 0 1 10330
box -6 -8 86 248
use OAI21X1  _8831_
timestamp 0
transform -1 0 7150 0 1 10330
box -6 -8 106 248
use OAI21X1  _8832_
timestamp 0
transform 1 0 4770 0 -1 8890
box -6 -8 106 248
use OAI21X1  _8833_
timestamp 0
transform -1 0 5010 0 -1 8890
box -6 -8 106 248
use OAI21X1  _8834_
timestamp 0
transform 1 0 5530 0 1 8410
box -6 -8 106 248
use OAI21X1  _8835_
timestamp 0
transform 1 0 5670 0 1 8410
box -6 -8 106 248
use NAND2X1  _8836_
timestamp 0
transform -1 0 5430 0 -1 9850
box -6 -8 86 248
use OAI21X1  _8837_
timestamp 0
transform -1 0 5590 0 -1 9850
box -6 -8 106 248
use NAND2X1  _8838_
timestamp 0
transform 1 0 5990 0 -1 9370
box -6 -8 86 248
use OAI21X1  _8839_
timestamp 0
transform -1 0 5950 0 -1 9370
box -6 -8 106 248
use DFFPOSX1  _8840_
timestamp 0
transform -1 0 4590 0 1 8890
box -6 -8 246 248
use DFFPOSX1  _8841_
timestamp 0
transform -1 0 4850 0 1 7930
box -6 -8 246 248
use DFFPOSX1  _8842_
timestamp 0
transform 1 0 6550 0 1 6490
box -6 -8 246 248
use DFFPOSX1  _8843_
timestamp 0
transform 1 0 4110 0 1 8890
box -6 -8 246 248
use DFFPOSX1  _8844_
timestamp 0
transform 1 0 3130 0 1 11290
box -6 -8 246 248
use DFFPOSX1  _8845_
timestamp 0
transform 1 0 3070 0 1 8410
box -6 -8 246 248
use DFFPOSX1  _8846_
timestamp 0
transform 1 0 2610 0 1 7930
box -6 -8 246 248
use DFFPOSX1  _8847_
timestamp 0
transform 1 0 2210 0 1 7930
box -6 -8 246 248
use DFFPOSX1  _8848_
timestamp 0
transform 1 0 2870 0 -1 8410
box -6 -8 246 248
use DFFPOSX1  _8849_
timestamp 0
transform 1 0 2230 0 -1 8410
box -6 -8 246 248
use DFFPOSX1  _8850_
timestamp 0
transform 1 0 3030 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _8851_
timestamp 0
transform 1 0 3030 0 -1 7930
box -6 -8 246 248
use DFFPOSX1  _8852_
timestamp 0
transform 1 0 3250 0 -1 7450
box -6 -8 246 248
use DFFPOSX1  _8853_
timestamp 0
transform 1 0 3110 0 -1 8410
box -6 -8 246 248
use DFFPOSX1  _8854_
timestamp 0
transform 1 0 2330 0 1 7450
box -6 -8 246 248
use DFFPOSX1  _8855_
timestamp 0
transform 1 0 3650 0 -1 7930
box -6 -8 246 248
use DFFPOSX1  _8856_
timestamp 0
transform 1 0 2510 0 -1 7930
box -6 -8 246 248
use DFFPOSX1  _8857_
timestamp 0
transform 1 0 3990 0 -1 8410
box -6 -8 246 248
use DFFPOSX1  _8858_
timestamp 0
transform -1 0 4850 0 1 10810
box -6 -8 246 248
use DFFPOSX1  _8859_
timestamp 0
transform 1 0 3790 0 1 7930
box -6 -8 246 248
use DFFPOSX1  _8860_
timestamp 0
transform 1 0 4110 0 -1 11290
box -6 -8 246 248
use DFFPOSX1  _8861_
timestamp 0
transform 1 0 2810 0 1 6970
box -6 -8 246 248
use DFFPOSX1  _8862_
timestamp 0
transform 1 0 2750 0 -1 7450
box -6 -8 246 248
use DFFPOSX1  _8863_
timestamp 0
transform 1 0 3830 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _8864_
timestamp 0
transform 1 0 2550 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _8865_
timestamp 0
transform -1 0 5110 0 1 7450
box -6 -8 246 248
use DFFPOSX1  _8866_
timestamp 0
transform -1 0 6590 0 -1 8410
box -6 -8 246 248
use DFFPOSX1  _8867_
timestamp 0
transform -1 0 6530 0 1 7930
box -6 -8 246 248
use DFFPOSX1  _8868_
timestamp 0
transform -1 0 5950 0 1 7930
box -6 -8 246 248
use DFFPOSX1  _8869_
timestamp 0
transform -1 0 8050 0 -1 7930
box -6 -8 246 248
use DFFPOSX1  _8870_
timestamp 0
transform -1 0 6750 0 1 6970
box -6 -8 246 248
use DFFPOSX1  _8871_
timestamp 0
transform -1 0 7210 0 1 7930
box -6 -8 246 248
use DFFPOSX1  _8872_
timestamp 0
transform -1 0 6530 0 -1 7450
box -6 -8 246 248
use DFFPOSX1  _8873_
timestamp 0
transform -1 0 5870 0 1 7450
box -6 -8 246 248
use DFFPOSX1  _8874_
timestamp 0
transform -1 0 5750 0 -1 6490
box -6 -8 246 248
use DFFPOSX1  _8875_
timestamp 0
transform -1 0 5170 0 -1 6490
box -6 -8 246 248
use DFFPOSX1  _8876_
timestamp 0
transform -1 0 4650 0 1 6490
box -6 -8 246 248
use DFFPOSX1  _8877_
timestamp 0
transform -1 0 1010 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _8878_
timestamp 0
transform 1 0 10 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _8879_
timestamp 0
transform -1 0 3990 0 -1 8410
box -6 -8 246 248
use DFFPOSX1  _8880_
timestamp 0
transform -1 0 4590 0 -1 8890
box -6 -8 246 248
use DFFPOSX1  _8881_
timestamp 0
transform -1 0 3650 0 1 8890
box -6 -8 246 248
use DFFPOSX1  _8882_
timestamp 0
transform -1 0 5230 0 1 9370
box -6 -8 246 248
use DFFPOSX1  _8883_
timestamp 0
transform -1 0 3770 0 -1 10810
box -6 -8 246 248
use DFFPOSX1  _8884_
timestamp 0
transform 1 0 2910 0 -1 9850
box -6 -8 246 248
use DFFPOSX1  _8885_
timestamp 0
transform 1 0 3870 0 1 8890
box -6 -8 246 248
use DFFPOSX1  _8886_
timestamp 0
transform -1 0 4930 0 -1 9370
box -6 -8 246 248
use DFFPOSX1  _8887_
timestamp 0
transform -1 0 3410 0 1 8890
box -6 -8 246 248
use DFFPOSX1  _8888_
timestamp 0
transform -1 0 2950 0 -1 9370
box -6 -8 246 248
use DFFPOSX1  _8889_
timestamp 0
transform -1 0 1110 0 -1 7450
box -6 -8 246 248
use DFFPOSX1  _8890_
timestamp 0
transform -1 0 1510 0 -1 7450
box -6 -8 246 248
use DFFPOSX1  _8891_
timestamp 0
transform -1 0 4750 0 1 8410
box -6 -8 246 248
use DFFPOSX1  _8892_
timestamp 0
transform -1 0 3650 0 1 8410
box -6 -8 246 248
use DFFPOSX1  _8893_
timestamp 0
transform -1 0 5090 0 1 10810
box -6 -8 246 248
use DFFPOSX1  _8894_
timestamp 0
transform -1 0 3610 0 -1 9370
box -6 -8 246 248
use DFFPOSX1  _8895_
timestamp 0
transform -1 0 2170 0 1 11770
box -6 -8 246 248
use DFFPOSX1  _8896_
timestamp 0
transform -1 0 1710 0 1 11770
box -6 -8 246 248
use DFFPOSX1  _8897_
timestamp 0
transform -1 0 4550 0 -1 9370
box -6 -8 246 248
use DFFPOSX1  _8898_
timestamp 0
transform -1 0 3850 0 -1 9370
box -6 -8 246 248
use DFFPOSX1  _8899_
timestamp 0
transform 1 0 5430 0 -1 10330
box -6 -8 246 248
use DFFPOSX1  _8900_
timestamp 0
transform 1 0 5670 0 -1 10810
box -6 -8 246 248
use DFFPOSX1  _8901_
timestamp 0
transform 1 0 4990 0 1 6970
box -6 -8 246 248
use DFFPOSX1  _8902_
timestamp 0
transform 1 0 5110 0 1 7450
box -6 -8 246 248
use DFFPOSX1  _8903_
timestamp 0
transform -1 0 6030 0 -1 7930
box -6 -8 246 248
use DFFPOSX1  _8904_
timestamp 0
transform 1 0 6190 0 -1 7930
box -6 -8 246 248
use DFFPOSX1  _8905_
timestamp 0
transform 1 0 5450 0 -1 8890
box -6 -8 246 248
use DFFPOSX1  _8906_
timestamp 0
transform 1 0 6370 0 1 10330
box -6 -8 246 248
use DFFPOSX1  _8907_
timestamp 0
transform 1 0 6870 0 1 9850
box -6 -8 246 248
use DFFPOSX1  _8908_
timestamp 0
transform 1 0 7150 0 1 10330
box -6 -8 246 248
use DFFPOSX1  _8909_
timestamp 0
transform 1 0 4830 0 1 8890
box -6 -8 246 248
use DFFPOSX1  _8910_
timestamp 0
transform 1 0 5590 0 -1 8410
box -6 -8 246 248
use DFFPOSX1  _8911_
timestamp 0
transform 1 0 5750 0 1 9850
box -6 -8 246 248
use DFFPOSX1  _8912_
timestamp 0
transform 1 0 5790 0 1 9370
box -6 -8 246 248
use DFFPOSX1  _8913_
timestamp 0
transform -1 0 5730 0 1 6970
box -6 -8 246 248
use DFFPOSX1  _8914_
timestamp 0
transform 1 0 5010 0 1 7930
box -6 -8 246 248
use DFFPOSX1  _8915_
timestamp 0
transform 1 0 5250 0 -1 7930
box -6 -8 246 248
use DFFPOSX1  _8916_
timestamp 0
transform -1 0 4830 0 1 6970
box -6 -8 246 248
use DFFPOSX1  _8917_
timestamp 0
transform -1 0 4310 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _8918_
timestamp 0
transform -1 0 4450 0 1 6970
box -6 -8 246 248
use DFFPOSX1  _8919_
timestamp 0
transform 1 0 3270 0 -1 6970
box -6 -8 246 248
use INVX1  _8920_
timestamp 0
transform 1 0 290 0 1 6490
box -6 -8 66 248
use INVX2  _8921_
timestamp 0
transform -1 0 2890 0 -1 5050
box -6 -8 66 248
use NOR2X1  _8922_
timestamp 0
transform -1 0 3010 0 -1 5050
box -6 -8 86 248
use INVX2  _8923_
timestamp 0
transform -1 0 4250 0 -1 4570
box -6 -8 66 248
use NOR2X1  _8924_
timestamp 0
transform -1 0 4150 0 -1 5530
box -6 -8 86 248
use INVX4  _8925_
timestamp 0
transform 1 0 4990 0 1 4570
box -6 -8 86 248
use NOR2X1  _8926_
timestamp 0
transform -1 0 4390 0 -1 5050
box -6 -8 86 248
use OAI21X1  _8927_
timestamp 0
transform 1 0 4190 0 -1 5530
box -6 -8 106 248
use INVX2  _8928_
timestamp 0
transform 1 0 4570 0 1 5050
box -6 -8 66 248
use AND2X2  _8929_
timestamp 0
transform -1 0 4710 0 1 4570
box -6 -8 106 248
use AOI22X1  _8930_
timestamp 0
transform 1 0 4490 0 1 5530
box -6 -8 126 248
use OAI21X1  _8931_
timestamp 0
transform 1 0 4210 0 1 5530
box -6 -8 106 248
use NOR2X1  _8932_
timestamp 0
transform 1 0 4010 0 1 4570
box -6 -8 86 248
use AOI22X1  _8933_
timestamp 0
transform 1 0 4030 0 1 5530
box -6 -8 126 248
use OAI21X1  _8934_
timestamp 0
transform 1 0 3750 0 1 5530
box -6 -8 106 248
use INVX1  _8935_
timestamp 0
transform 1 0 3650 0 1 5530
box -6 -8 66 248
use OAI21X1  _8936_
timestamp 0
transform 1 0 4350 0 -1 5530
box -6 -8 106 248
use AOI21X1  _8937_
timestamp 0
transform 1 0 4490 0 -1 5530
box -6 -8 106 248
use INVX1  _8938_
timestamp 0
transform 1 0 4930 0 1 6010
box -6 -8 66 248
use NAND2X1  _8939_
timestamp 0
transform -1 0 4710 0 -1 5530
box -6 -8 86 248
use OAI21X1  _8940_
timestamp 0
transform -1 0 5050 0 1 5530
box -6 -8 106 248
use OAI21X1  _8941_
timestamp 0
transform -1 0 4890 0 1 5530
box -6 -8 106 248
use AOI22X1  _8942_
timestamp 0
transform 1 0 3110 0 1 5530
box -6 -8 126 248
use NAND2X1  _8943_
timestamp 0
transform 1 0 4670 0 1 5530
box -6 -8 86 248
use INVX1  _8944_
timestamp 0
transform 1 0 5190 0 1 1690
box -6 -8 66 248
use OAI21X1  _8945_
timestamp 0
transform 1 0 5630 0 -1 2650
box -6 -8 106 248
use AOI21X1  _8946_
timestamp 0
transform 1 0 5470 0 -1 2650
box -6 -8 106 248
use INVX1  _8947_
timestamp 0
transform 1 0 6250 0 1 2650
box -6 -8 66 248
use NAND2X1  _8948_
timestamp 0
transform -1 0 6130 0 -1 2650
box -6 -8 86 248
use OAI21X1  _8949_
timestamp 0
transform 1 0 5690 0 1 2650
box -6 -8 106 248
use OAI21X1  _8950_
timestamp 0
transform -1 0 5490 0 1 2650
box -6 -8 106 248
use AOI22X1  _8951_
timestamp 0
transform -1 0 4150 0 -1 4570
box -6 -8 126 248
use NAND2X1  _8952_
timestamp 0
transform 1 0 4790 0 -1 4570
box -6 -8 86 248
use INVX1  _8953_
timestamp 0
transform -1 0 5130 0 1 3130
box -6 -8 66 248
use OAI21X1  _8954_
timestamp 0
transform -1 0 5990 0 -1 2650
box -6 -8 106 248
use AOI21X1  _8955_
timestamp 0
transform 1 0 5610 0 -1 3130
box -6 -8 106 248
use INVX1  _8956_
timestamp 0
transform 1 0 4990 0 1 3610
box -6 -8 66 248
use NAND2X1  _8957_
timestamp 0
transform -1 0 5030 0 1 3130
box -6 -8 86 248
use OAI21X1  _8958_
timestamp 0
transform -1 0 5070 0 -1 3610
box -6 -8 106 248
use OAI21X1  _8959_
timestamp 0
transform -1 0 5230 0 -1 3610
box -6 -8 106 248
use AOI22X1  _8960_
timestamp 0
transform 1 0 4710 0 -1 4090
box -6 -8 126 248
use NAND2X1  _8961_
timestamp 0
transform 1 0 5090 0 1 3610
box -6 -8 86 248
use INVX1  _8962_
timestamp 0
transform 1 0 3610 0 -1 730
box -6 -8 66 248
use OAI21X1  _8963_
timestamp 0
transform -1 0 4910 0 -1 2650
box -6 -8 106 248
use AOI21X1  _8964_
timestamp 0
transform 1 0 4550 0 -1 2650
box -6 -8 106 248
use INVX1  _8965_
timestamp 0
transform -1 0 5890 0 -1 2170
box -6 -8 66 248
use NAND2X1  _8966_
timestamp 0
transform 1 0 5770 0 -1 2650
box -6 -8 86 248
use OAI21X1  _8967_
timestamp 0
transform -1 0 5650 0 1 2650
box -6 -8 106 248
use OAI21X1  _8968_
timestamp 0
transform 1 0 5230 0 1 2650
box -6 -8 106 248
use AOI22X1  _8969_
timestamp 0
transform -1 0 4130 0 1 3610
box -6 -8 126 248
use NAND2X1  _8970_
timestamp 0
transform -1 0 4930 0 -1 3610
box -6 -8 86 248
use INVX1  _8971_
timestamp 0
transform 1 0 5990 0 1 2170
box -6 -8 66 248
use NOR2X1  _8972_
timestamp 0
transform -1 0 4490 0 -1 2650
box -6 -8 86 248
use OAI21X1  _8973_
timestamp 0
transform 1 0 4630 0 1 2650
box -6 -8 106 248
use AOI22X1  _8974_
timestamp 0
transform 1 0 4250 0 -1 2650
box -6 -8 126 248
use OAI21X1  _8975_
timestamp 0
transform -1 0 4590 0 1 2650
box -6 -8 106 248
use AOI22X1  _8976_
timestamp 0
transform 1 0 4190 0 1 3610
box -6 -8 126 248
use OAI21X1  _8977_
timestamp 0
transform -1 0 4450 0 1 3610
box -6 -8 106 248
use INVX1  _8978_
timestamp 0
transform -1 0 3990 0 -1 4570
box -6 -8 66 248
use INVX1  _8979_
timestamp 0
transform -1 0 2470 0 1 4090
box -6 -8 66 248
use INVX8  _8980_
timestamp 0
transform -1 0 170 0 1 3610
box -6 -8 126 248
use INVX8  _8981_
timestamp 0
transform -1 0 430 0 -1 4090
box -6 -8 126 248
use INVX1  _8982_
timestamp 0
transform 1 0 1470 0 -1 2650
box -6 -8 66 248
use NAND2X1  _8983_
timestamp 0
transform -1 0 1330 0 -1 3130
box -6 -8 86 248
use OAI21X1  _8984_
timestamp 0
transform -1 0 1470 0 -1 3130
box -6 -8 106 248
use INVX1  _8985_
timestamp 0
transform -1 0 1130 0 -1 2170
box -6 -8 66 248
use NAND2X1  _8986_
timestamp 0
transform -1 0 1010 0 1 3130
box -6 -8 86 248
use OAI21X1  _8987_
timestamp 0
transform -1 0 1150 0 1 3130
box -6 -8 106 248
use MUX2X1  _8988_
timestamp 0
transform -1 0 1330 0 1 3130
box -6 -8 126 248
use INVX1  _8989_
timestamp 0
transform 1 0 930 0 -1 4090
box -6 -8 66 248
use NAND2X1  _8990_
timestamp 0
transform -1 0 750 0 -1 4090
box -6 -8 86 248
use OAI21X1  _8991_
timestamp 0
transform -1 0 890 0 -1 4090
box -6 -8 106 248
use INVX1  _8992_
timestamp 0
transform -1 0 1650 0 -1 4090
box -6 -8 66 248
use NAND2X1  _8993_
timestamp 0
transform 1 0 1470 0 -1 4090
box -6 -8 86 248
use OAI21X1  _8994_
timestamp 0
transform -1 0 1510 0 1 3610
box -6 -8 106 248
use MUX2X1  _8995_
timestamp 0
transform 1 0 1090 0 1 3610
box -6 -8 126 248
use MUX2X1  _8996_
timestamp 0
transform 1 0 1250 0 1 3610
box -6 -8 126 248
use NOR2X1  _8997_
timestamp 0
transform -1 0 2590 0 1 4090
box -6 -8 86 248
use NAND2X1  _8998_
timestamp 0
transform -1 0 2350 0 1 4090
box -6 -8 86 248
use INVX1  _8999_
timestamp 0
transform -1 0 2690 0 1 4090
box -6 -8 66 248
use NAND2X1  _9000_
timestamp 0
transform -1 0 550 0 1 3610
box -6 -8 86 248
use OAI21X1  _9001_
timestamp 0
transform 1 0 3570 0 -1 1690
box -6 -8 106 248
use INVX2  _9002_
timestamp 0
transform 1 0 3470 0 1 250
box -6 -8 66 248
use OAI21X1  _9003_
timestamp 0
transform 1 0 2730 0 1 4090
box -6 -8 106 248
use OAI21X1  _9004_
timestamp 0
transform -1 0 3650 0 -1 4570
box -6 -8 106 248
use INVX8  _9005_
timestamp 0
transform 1 0 4550 0 -1 3610
box -6 -8 126 248
use NAND2X1  _9006_
timestamp 0
transform 1 0 4590 0 -1 4090
box -6 -8 86 248
use NOR2X1  _9007_
timestamp 0
transform -1 0 3690 0 1 1690
box -6 -8 86 248
use MUX2X1  _9008_
timestamp 0
transform -1 0 570 0 -1 3130
box -6 -8 126 248
use MUX2X1  _9009_
timestamp 0
transform -1 0 710 0 1 3130
box -6 -8 126 248
use MUX2X1  _9010_
timestamp 0
transform 1 0 410 0 1 3130
box -6 -8 126 248
use INVX2  _9011_
timestamp 0
transform 1 0 50 0 1 5050
box -6 -8 66 248
use NAND2X1  _9012_
timestamp 0
transform -1 0 290 0 1 4090
box -6 -8 86 248
use AOI21X1  _9013_
timestamp 0
transform 1 0 330 0 1 4090
box -6 -8 106 248
use NAND3X1  _9014_
timestamp 0
transform -1 0 730 0 1 4090
box -6 -8 106 248
use NAND3X1  _9015_
timestamp 0
transform -1 0 870 0 1 4090
box -6 -8 106 248
use NAND3X1  _9016_
timestamp 0
transform -1 0 570 0 1 4090
box -6 -8 106 248
use OAI22X1  _9017_
timestamp 0
transform 1 0 490 0 -1 4090
box -6 -8 126 248
use INVX1  _9018_
timestamp 0
transform -1 0 1370 0 1 4570
box -6 -8 66 248
use INVX8  _9019_
timestamp 0
transform -1 0 290 0 1 5050
box -6 -8 126 248
use INVX1  _9020_
timestamp 0
transform -1 0 1130 0 -1 1210
box -6 -8 66 248
use NAND2X1  _9021_
timestamp 0
transform -1 0 910 0 -1 1690
box -6 -8 86 248
use OAI21X1  _9022_
timestamp 0
transform -1 0 1050 0 -1 1690
box -6 -8 106 248
use INVX1  _9023_
timestamp 0
transform -1 0 1730 0 -1 3130
box -6 -8 66 248
use NAND2X1  _9024_
timestamp 0
transform -1 0 1350 0 1 2650
box -6 -8 86 248
use OAI21X1  _9025_
timestamp 0
transform -1 0 1490 0 1 2650
box -6 -8 106 248
use MUX2X1  _9026_
timestamp 0
transform 1 0 1090 0 1 2650
box -6 -8 126 248
use INVX1  _9027_
timestamp 0
transform 1 0 930 0 -1 3610
box -6 -8 66 248
use NAND2X1  _9028_
timestamp 0
transform 1 0 1530 0 1 2650
box -6 -8 86 248
use OAI21X1  _9029_
timestamp 0
transform -1 0 1630 0 -1 3130
box -6 -8 106 248
use INVX1  _9030_
timestamp 0
transform -1 0 1250 0 1 4090
box -6 -8 66 248
use NAND2X1  _9031_
timestamp 0
transform 1 0 1730 0 -1 3610
box -6 -8 86 248
use OAI21X1  _9032_
timestamp 0
transform 1 0 1670 0 1 3130
box -6 -8 106 248
use MUX2X1  _9033_
timestamp 0
transform 1 0 1510 0 1 3130
box -6 -8 126 248
use MUX2X1  _9034_
timestamp 0
transform 1 0 1550 0 -1 3610
box -6 -8 126 248
use NAND3X1  _9035_
timestamp 0
transform 1 0 1550 0 1 3610
box -6 -8 106 248
use MUX2X1  _9036_
timestamp 0
transform 1 0 770 0 1 2650
box -6 -8 126 248
use MUX2X1  _9037_
timestamp 0
transform 1 0 750 0 1 3130
box -6 -8 126 248
use MUX2X1  _9038_
timestamp 0
transform -1 0 910 0 -1 3130
box -6 -8 126 248
use MUX2X1  _9039_
timestamp 0
transform -1 0 890 0 -1 3610
box -6 -8 126 248
use MUX2X1  _9040_
timestamp 0
transform -1 0 1170 0 -1 4090
box -6 -8 126 248
use MUX2X1  _9041_
timestamp 0
transform 1 0 750 0 1 3610
box -6 -8 126 248
use MUX2X1  _9042_
timestamp 0
transform -1 0 1030 0 1 3610
box -6 -8 126 248
use OAI21X1  _9043_
timestamp 0
transform -1 0 1810 0 -1 4090
box -6 -8 106 248
use AOI21X1  _9044_
timestamp 0
transform -1 0 1670 0 1 4090
box -6 -8 106 248
use INVX1  _9045_
timestamp 0
transform 1 0 1870 0 1 4090
box -6 -8 66 248
use NAND3X1  _9046_
timestamp 0
transform 1 0 1710 0 1 4090
box -6 -8 106 248
use AND2X2  _9047_
timestamp 0
transform 1 0 1970 0 1 4090
box -6 -8 106 248
use OAI21X1  _9048_
timestamp 0
transform 1 0 2690 0 -1 4090
box -6 -8 106 248
use OR2X2  _9049_
timestamp 0
transform 1 0 2830 0 -1 4090
box -6 -8 106 248
use AOI21X1  _9050_
timestamp 0
transform 1 0 2990 0 -1 4090
box -6 -8 106 248
use OAI21X1  _9051_
timestamp 0
transform 1 0 4210 0 -1 4090
box -6 -8 106 248
use INVX1  _9052_
timestamp 0
transform 1 0 7550 0 1 6490
box -6 -8 66 248
use NAND2X1  _9053_
timestamp 0
transform -1 0 7010 0 1 6490
box -6 -8 86 248
use OAI21X1  _9054_
timestamp 0
transform 1 0 7150 0 1 6490
box -6 -8 106 248
use NAND2X1  _9055_
timestamp 0
transform -1 0 4070 0 1 4090
box -6 -8 86 248
use AOI21X1  _9056_
timestamp 0
transform -1 0 2210 0 1 4090
box -6 -8 106 248
use MUX2X1  _9057_
timestamp 0
transform -1 0 590 0 1 2650
box -6 -8 126 248
use MUX2X1  _9058_
timestamp 0
transform 1 0 610 0 -1 3130
box -6 -8 126 248
use MUX2X1  _9059_
timestamp 0
transform -1 0 730 0 -1 3610
box -6 -8 126 248
use NAND2X1  _9060_
timestamp 0
transform -1 0 410 0 -1 3610
box -6 -8 86 248
use OAI22X1  _9061_
timestamp 0
transform 1 0 450 0 -1 3610
box -6 -8 126 248
use AOI21X1  _9062_
timestamp 0
transform 1 0 610 0 1 3610
box -6 -8 106 248
use AOI21X1  _9063_
timestamp 0
transform 1 0 1990 0 -1 4090
box -6 -8 106 248
use NAND2X1  _9064_
timestamp 0
transform 1 0 2150 0 -1 4090
box -6 -8 86 248
use INVX1  _9065_
timestamp 0
transform 1 0 2110 0 1 3610
box -6 -8 66 248
use OAI21X1  _9066_
timestamp 0
transform 1 0 1690 0 1 3610
box -6 -8 106 248
use NAND2X1  _9067_
timestamp 0
transform 1 0 1990 0 1 3610
box -6 -8 86 248
use AOI21X1  _9068_
timestamp 0
transform 1 0 2430 0 -1 4090
box -6 -8 106 248
use NAND3X1  _9069_
timestamp 0
transform 1 0 2290 0 -1 4090
box -6 -8 106 248
use INVX1  _9070_
timestamp 0
transform 1 0 3290 0 -1 4090
box -6 -8 66 248
use OR2X2  _9071_
timestamp 0
transform 1 0 3570 0 -1 4090
box -6 -8 106 248
use NOR2X1  _9072_
timestamp 0
transform 1 0 3710 0 -1 4090
box -6 -8 86 248
use INVX1  _9073_
timestamp 0
transform 1 0 3830 0 -1 4090
box -6 -8 66 248
use OAI21X1  _9074_
timestamp 0
transform -1 0 3510 0 -1 4090
box -6 -8 106 248
use AOI21X1  _9075_
timestamp 0
transform 1 0 3930 0 -1 4090
box -6 -8 106 248
use INVX2  _9076_
timestamp 0
transform 1 0 4050 0 -1 3130
box -6 -8 66 248
use OAI21X1  _9077_
timestamp 0
transform 1 0 4390 0 -1 3610
box -6 -8 106 248
use OAI21X1  _9078_
timestamp 0
transform -1 0 4170 0 -1 4090
box -6 -8 106 248
use INVX1  _9079_
timestamp 0
transform 1 0 4890 0 -1 4090
box -6 -8 66 248
use INVX2  _9080_
timestamp 0
transform 1 0 4490 0 1 3610
box -6 -8 66 248
use OAI21X1  _9081_
timestamp 0
transform 1 0 3150 0 -1 4090
box -6 -8 106 248
use INVX1  _9082_
timestamp 0
transform 1 0 3990 0 -1 3610
box -6 -8 66 248
use INVX1  _9083_
timestamp 0
transform -1 0 3010 0 -1 3610
box -6 -8 66 248
use NAND3X1  _9084_
timestamp 0
transform 1 0 1850 0 -1 4090
box -6 -8 106 248
use INVX1  _9085_
timestamp 0
transform 1 0 570 0 -1 1690
box -6 -8 66 248
use NAND2X1  _9086_
timestamp 0
transform -1 0 430 0 -1 1690
box -6 -8 86 248
use OAI21X1  _9087_
timestamp 0
transform -1 0 770 0 -1 1690
box -6 -8 106 248
use NAND2X1  _9088_
timestamp 0
transform -1 0 1030 0 1 2650
box -6 -8 86 248
use OAI21X1  _9089_
timestamp 0
transform 1 0 930 0 -1 2650
box -6 -8 106 248
use NOR2X1  _9090_
timestamp 0
transform -1 0 1730 0 -1 2170
box -6 -8 86 248
use NOR2X1  _9091_
timestamp 0
transform 1 0 1570 0 -1 4570
box -6 -8 86 248
use AOI22X1  _9092_
timestamp 0
transform 1 0 1650 0 1 2650
box -6 -8 126 248
use OAI21X1  _9093_
timestamp 0
transform 1 0 1590 0 -1 2650
box -6 -8 106 248
use NAND3X1  _9094_
timestamp 0
transform 1 0 2650 0 -1 3610
box -6 -8 106 248
use INVX1  _9095_
timestamp 0
transform -1 0 2750 0 1 3130
box -6 -8 66 248
use INVX1  _9096_
timestamp 0
transform -1 0 2850 0 1 3130
box -6 -8 66 248
use OAI21X1  _9097_
timestamp 0
transform -1 0 2890 0 -1 3610
box -6 -8 106 248
use NAND3X1  _9098_
timestamp 0
transform 1 0 3210 0 -1 3610
box -6 -8 106 248
use AOI21X1  _9099_
timestamp 0
transform 1 0 3050 0 -1 3610
box -6 -8 106 248
use INVX1  _9100_
timestamp 0
transform 1 0 3530 0 -1 3610
box -6 -8 66 248
use NAND2X1  _9101_
timestamp 0
transform 1 0 3630 0 -1 3610
box -6 -8 86 248
use AOI21X1  _9102_
timestamp 0
transform 1 0 4110 0 -1 3610
box -6 -8 106 248
use OAI21X1  _9103_
timestamp 0
transform 1 0 4250 0 -1 3610
box -6 -8 106 248
use AOI22X1  _9104_
timestamp 0
transform -1 0 4710 0 1 3610
box -6 -8 126 248
use AOI21X1  _9105_
timestamp 0
transform 1 0 3370 0 -1 3610
box -6 -8 106 248
use INVX1  _9106_
timestamp 0
transform 1 0 3570 0 1 3130
box -6 -8 66 248
use INVX1  _9107_
timestamp 0
transform -1 0 290 0 1 2650
box -6 -8 66 248
use NAND2X1  _9108_
timestamp 0
transform -1 0 470 0 -1 2650
box -6 -8 86 248
use OAI21X1  _9109_
timestamp 0
transform 1 0 510 0 -1 2650
box -6 -8 106 248
use NAND2X1  _9110_
timestamp 0
transform 1 0 670 0 -1 2650
box -6 -8 86 248
use OAI21X1  _9111_
timestamp 0
transform -1 0 890 0 -1 2650
box -6 -8 106 248
use NAND2X1  _9112_
timestamp 0
transform -1 0 1050 0 -1 3130
box -6 -8 86 248
use OAI21X1  _9113_
timestamp 0
transform -1 0 1190 0 -1 3130
box -6 -8 106 248
use INVX2  _9114_
timestamp 0
transform 1 0 3370 0 -1 3130
box -6 -8 66 248
use OAI21X1  _9115_
timestamp 0
transform 1 0 3230 0 1 2650
box -6 -8 106 248
use OR2X2  _9116_
timestamp 0
transform 1 0 3650 0 1 2650
box -6 -8 106 248
use NOR2X1  _9117_
timestamp 0
transform -1 0 3050 0 1 2650
box -6 -8 86 248
use OAI21X1  _9118_
timestamp 0
transform 1 0 3090 0 1 2650
box -6 -8 106 248
use NAND3X1  _9119_
timestamp 0
transform 1 0 3970 0 1 2650
box -6 -8 106 248
use NOR2X1  _9120_
timestamp 0
transform -1 0 3690 0 -1 3130
box -6 -8 86 248
use AND2X2  _9121_
timestamp 0
transform -1 0 3570 0 -1 3130
box -6 -8 106 248
use OAI21X1  _9122_
timestamp 0
transform 1 0 3750 0 -1 3130
box -6 -8 106 248
use NAND2X1  _9123_
timestamp 0
transform 1 0 4370 0 1 2650
box -6 -8 86 248
use AOI21X1  _9124_
timestamp 0
transform 1 0 4950 0 1 2650
box -6 -8 106 248
use OAI21X1  _9125_
timestamp 0
transform 1 0 5090 0 1 2650
box -6 -8 106 248
use AOI22X1  _9126_
timestamp 0
transform -1 0 5970 0 1 2650
box -6 -8 126 248
use OAI21X1  _9127_
timestamp 0
transform -1 0 4390 0 -1 3130
box -6 -8 106 248
use INVX1  _9128_
timestamp 0
transform 1 0 2850 0 -1 3130
box -6 -8 66 248
use NAND3X1  _9129_
timestamp 0
transform 1 0 2970 0 -1 3130
box -6 -8 106 248
use NAND2X1  _9130_
timestamp 0
transform -1 0 530 0 1 2170
box -6 -8 86 248
use INVX1  _9131_
timestamp 0
transform 1 0 590 0 1 2170
box -6 -8 66 248
use AOI21X1  _9132_
timestamp 0
transform 1 0 1010 0 1 2170
box -6 -8 106 248
use NAND2X1  _9133_
timestamp 0
transform -1 0 1170 0 -1 2650
box -6 -8 86 248
use OAI21X1  _9134_
timestamp 0
transform -1 0 1430 0 -1 2650
box -6 -8 106 248
use NAND3X1  _9135_
timestamp 0
transform 1 0 2650 0 1 2650
box -6 -8 106 248
use NOR3X1  _9136_
timestamp 0
transform -1 0 3310 0 -1 3130
box -6 -8 186 248
use INVX1  _9137_
timestamp 0
transform -1 0 2770 0 -1 2650
box -6 -8 66 248
use OAI21X1  _9138_
timestamp 0
transform -1 0 2930 0 -1 2650
box -6 -8 106 248
use NAND3X1  _9139_
timestamp 0
transform 1 0 3390 0 -1 2650
box -6 -8 106 248
use AOI21X1  _9140_
timestamp 0
transform 1 0 3250 0 -1 2650
box -6 -8 106 248
use INVX1  _9141_
timestamp 0
transform -1 0 3610 0 -1 2650
box -6 -8 66 248
use NAND2X1  _9142_
timestamp 0
transform -1 0 3730 0 -1 2650
box -6 -8 86 248
use AND2X2  _9143_
timestamp 0
transform 1 0 4450 0 -1 3130
box -6 -8 106 248
use OAI21X1  _9144_
timestamp 0
transform 1 0 4590 0 -1 3130
box -6 -8 106 248
use OAI21X1  _9145_
timestamp 0
transform 1 0 4750 0 -1 3130
box -6 -8 106 248
use OAI21X1  _9146_
timestamp 0
transform -1 0 4810 0 -1 3610
box -6 -8 106 248
use INVX1  _9147_
timestamp 0
transform -1 0 6390 0 -1 2170
box -6 -8 66 248
use INVX1  _9148_
timestamp 0
transform 1 0 4550 0 1 2170
box -6 -8 66 248
use NAND3X1  _9149_
timestamp 0
transform 1 0 3110 0 -1 2650
box -6 -8 106 248
use AOI21X1  _9150_
timestamp 0
transform 1 0 710 0 1 2170
box -6 -8 106 248
use NAND2X1  _9151_
timestamp 0
transform -1 0 710 0 1 2650
box -6 -8 86 248
use OAI21X1  _9152_
timestamp 0
transform -1 0 970 0 1 2170
box -6 -8 106 248
use NAND3X1  _9153_
timestamp 0
transform 1 0 4110 0 1 2170
box -6 -8 106 248
use INVX1  _9154_
timestamp 0
transform -1 0 3390 0 1 2170
box -6 -8 66 248
use OAI21X1  _9155_
timestamp 0
transform 1 0 2810 0 1 2650
box -6 -8 106 248
use NAND2X1  _9156_
timestamp 0
transform -1 0 3630 0 1 2170
box -6 -8 86 248
use NAND3X1  _9157_
timestamp 0
transform 1 0 4950 0 1 2170
box -6 -8 106 248
use NAND3X1  _9158_
timestamp 0
transform 1 0 3670 0 1 2170
box -6 -8 106 248
use NAND2X1  _9159_
timestamp 0
transform -1 0 3510 0 1 2170
box -6 -8 86 248
use NAND3X1  _9160_
timestamp 0
transform 1 0 3830 0 1 2170
box -6 -8 106 248
use NAND2X1  _9161_
timestamp 0
transform 1 0 5050 0 -1 2170
box -6 -8 86 248
use AOI21X1  _9162_
timestamp 0
transform 1 0 3810 0 1 2650
box -6 -8 106 248
use NOR2X1  _9163_
timestamp 0
transform 1 0 4110 0 1 2650
box -6 -8 86 248
use OAI21X1  _9164_
timestamp 0
transform -1 0 4890 0 1 2650
box -6 -8 106 248
use NAND2X1  _9165_
timestamp 0
transform 1 0 4690 0 -1 2650
box -6 -8 86 248
use AOI21X1  _9166_
timestamp 0
transform 1 0 5170 0 -1 2170
box -6 -8 106 248
use OAI21X1  _9167_
timestamp 0
transform 1 0 5330 0 -1 2170
box -6 -8 106 248
use AOI22X1  _9168_
timestamp 0
transform -1 0 6290 0 -1 2170
box -6 -8 126 248
use INVX1  _9169_
timestamp 0
transform 1 0 5070 0 -1 3130
box -6 -8 66 248
use AOI21X1  _9170_
timestamp 0
transform -1 0 4890 0 1 2170
box -6 -8 106 248
use AND2X2  _9171_
timestamp 0
transform 1 0 4230 0 1 2650
box -6 -8 106 248
use NAND3X1  _9172_
timestamp 0
transform -1 0 4190 0 -1 2650
box -6 -8 106 248
use AOI21X1  _9173_
timestamp 0
transform -1 0 3870 0 -1 2650
box -6 -8 106 248
use OAI21X1  _9174_
timestamp 0
transform -1 0 4030 0 -1 2650
box -6 -8 106 248
use AOI21X1  _9175_
timestamp 0
transform -1 0 4750 0 1 2170
box -6 -8 106 248
use INVX1  _9176_
timestamp 0
transform -1 0 4270 0 -1 2170
box -6 -8 66 248
use NAND3X1  _9177_
timestamp 0
transform -1 0 3070 0 -1 2650
box -6 -8 106 248
use INVX1  _9178_
timestamp 0
transform 1 0 290 0 -1 2650
box -6 -8 66 248
use NOR2X1  _9179_
timestamp 0
transform -1 0 510 0 -1 2170
box -6 -8 86 248
use INVX1  _9180_
timestamp 0
transform 1 0 690 0 -1 2170
box -6 -8 66 248
use OAI21X1  _9181_
timestamp 0
transform -1 0 1610 0 -1 2170
box -6 -8 106 248
use NAND3X1  _9182_
timestamp 0
transform -1 0 3330 0 -1 2170
box -6 -8 106 248
use INVX1  _9183_
timestamp 0
transform -1 0 3450 0 -1 2170
box -6 -8 66 248
use OAI21X1  _9184_
timestamp 0
transform 1 0 3970 0 1 2170
box -6 -8 106 248
use NAND2X1  _9185_
timestamp 0
transform 1 0 3910 0 -1 2170
box -6 -8 86 248
use NAND3X1  _9186_
timestamp 0
transform 1 0 4050 0 -1 2170
box -6 -8 106 248
use NAND3X1  _9187_
timestamp 0
transform 1 0 3490 0 -1 2170
box -6 -8 106 248
use NAND2X1  _9188_
timestamp 0
transform 1 0 3790 0 -1 2170
box -6 -8 86 248
use NAND3X1  _9189_
timestamp 0
transform -1 0 3730 0 -1 2170
box -6 -8 106 248
use NAND2X1  _9190_
timestamp 0
transform -1 0 4230 0 1 1690
box -6 -8 86 248
use INVX1  _9191_
timestamp 0
transform 1 0 4290 0 1 1690
box -6 -8 66 248
use NOR2X1  _9192_
timestamp 0
transform 1 0 4530 0 1 1690
box -6 -8 86 248
use OAI21X1  _9193_
timestamp 0
transform 1 0 4910 0 -1 2170
box -6 -8 106 248
use OAI21X1  _9194_
timestamp 0
transform 1 0 4390 0 1 1690
box -6 -8 106 248
use OAI21X1  _9195_
timestamp 0
transform 1 0 4350 0 -1 1690
box -6 -8 106 248
use INVX1  _9196_
timestamp 0
transform 1 0 4790 0 -1 1690
box -6 -8 66 248
use OAI21X1  _9197_
timestamp 0
transform 1 0 4650 0 1 1690
box -6 -8 106 248
use OAI21X1  _9198_
timestamp 0
transform -1 0 5010 0 -1 3130
box -6 -8 106 248
use INVX1  _9199_
timestamp 0
transform -1 0 5110 0 -1 1690
box -6 -8 66 248
use OAI21X1  _9200_
timestamp 0
transform -1 0 3850 0 1 1690
box -6 -8 106 248
use NOR2X1  _9201_
timestamp 0
transform -1 0 4110 0 1 1690
box -6 -8 86 248
use AOI21X1  _9202_
timestamp 0
transform -1 0 3990 0 1 1690
box -6 -8 106 248
use INVX1  _9203_
timestamp 0
transform -1 0 2450 0 1 1210
box -6 -8 66 248
use OR2X2  _9204_
timestamp 0
transform -1 0 3310 0 -1 1690
box -6 -8 106 248
use OAI21X1  _9205_
timestamp 0
transform 1 0 1190 0 -1 2170
box -6 -8 106 248
use NAND3X1  _9206_
timestamp 0
transform -1 0 2890 0 -1 1690
box -6 -8 106 248
use NOR2X1  _9207_
timestamp 0
transform 1 0 2910 0 1 1690
box -6 -8 86 248
use INVX1  _9208_
timestamp 0
transform 1 0 2650 0 1 1690
box -6 -8 66 248
use OAI21X1  _9209_
timestamp 0
transform -1 0 2850 0 1 1690
box -6 -8 106 248
use NAND3X1  _9210_
timestamp 0
transform 1 0 2510 0 1 1210
box -6 -8 106 248
use NAND3X1  _9211_
timestamp 0
transform 1 0 2930 0 -1 1690
box -6 -8 106 248
use OAI21X1  _9212_
timestamp 0
transform 1 0 3050 0 1 1690
box -6 -8 106 248
use NAND3X1  _9213_
timestamp 0
transform 1 0 3070 0 -1 1690
box -6 -8 106 248
use AND2X2  _9214_
timestamp 0
transform 1 0 4230 0 1 1210
box -6 -8 106 248
use INVX1  _9215_
timestamp 0
transform 1 0 4510 0 1 1210
box -6 -8 66 248
use AOI21X1  _9216_
timestamp 0
transform 1 0 4490 0 -1 1690
box -6 -8 106 248
use OAI21X1  _9217_
timestamp 0
transform 1 0 4650 0 -1 1690
box -6 -8 106 248
use AOI22X1  _9218_
timestamp 0
transform -1 0 5010 0 -1 1690
box -6 -8 126 248
use NAND2X1  _9219_
timestamp 0
transform -1 0 4410 0 -1 2170
box -6 -8 86 248
use AND2X2  _9220_
timestamp 0
transform 1 0 4450 0 -1 2170
box -6 -8 106 248
use AND2X2  _9221_
timestamp 0
transform 1 0 5090 0 1 2170
box -6 -8 106 248
use NAND3X1  _9222_
timestamp 0
transform 1 0 4750 0 -1 2170
box -6 -8 106 248
use OAI21X1  _9223_
timestamp 0
transform -1 0 4690 0 -1 2170
box -6 -8 106 248
use INVX1  _9224_
timestamp 0
transform -1 0 4170 0 1 1210
box -6 -8 66 248
use AOI21X1  _9225_
timestamp 0
transform 1 0 4370 0 1 1210
box -6 -8 106 248
use INVX1  _9226_
timestamp 0
transform -1 0 3730 0 1 1210
box -6 -8 66 248
use NOR3X1  _9227_
timestamp 0
transform 1 0 3350 0 -1 1690
box -6 -8 186 248
use INVX1  _9228_
timestamp 0
transform 1 0 3550 0 1 1210
box -6 -8 66 248
use OAI21X1  _9229_
timestamp 0
transform 1 0 1350 0 -1 2170
box -6 -8 106 248
use NAND3X1  _9230_
timestamp 0
transform 1 0 3410 0 1 1210
box -6 -8 106 248
use INVX1  _9231_
timestamp 0
transform 1 0 3170 0 1 1210
box -6 -8 66 248
use OAI21X1  _9232_
timestamp 0
transform 1 0 3330 0 -1 1210
box -6 -8 106 248
use NAND3X1  _9233_
timestamp 0
transform 1 0 3470 0 -1 1210
box -6 -8 106 248
use NAND3X1  _9234_
timestamp 0
transform 1 0 3790 0 1 1210
box -6 -8 106 248
use OAI21X1  _9235_
timestamp 0
transform -1 0 3370 0 1 1210
box -6 -8 106 248
use NAND3X1  _9236_
timestamp 0
transform 1 0 3950 0 1 1210
box -6 -8 106 248
use AND2X2  _9237_
timestamp 0
transform 1 0 4050 0 -1 1210
box -6 -8 106 248
use AND2X2  _9238_
timestamp 0
transform 1 0 4490 0 -1 1210
box -6 -8 106 248
use OAI21X1  _9239_
timestamp 0
transform 1 0 4610 0 1 1210
box -6 -8 106 248
use OAI21X1  _9240_
timestamp 0
transform 1 0 4750 0 1 1210
box -6 -8 106 248
use OAI21X1  _9241_
timestamp 0
transform -1 0 5290 0 -1 3130
box -6 -8 106 248
use INVX1  _9242_
timestamp 0
transform -1 0 2330 0 1 1210
box -6 -8 66 248
use OAI21X1  _9243_
timestamp 0
transform 1 0 930 0 -1 2170
box -6 -8 106 248
use INVX1  _9244_
timestamp 0
transform 1 0 3430 0 1 730
box -6 -8 66 248
use AOI21X1  _9245_
timestamp 0
transform 1 0 3690 0 1 730
box -6 -8 106 248
use NAND3X1  _9246_
timestamp 0
transform 1 0 3530 0 1 730
box -6 -8 106 248
use NAND2X1  _9247_
timestamp 0
transform -1 0 3790 0 -1 730
box -6 -8 86 248
use NAND2X1  _9248_
timestamp 0
transform -1 0 3390 0 1 730
box -6 -8 86 248
use OAI21X1  _9249_
timestamp 0
transform 1 0 3830 0 1 730
box -6 -8 106 248
use NAND2X1  _9250_
timestamp 0
transform 1 0 3770 0 -1 1210
box -6 -8 86 248
use INVX1  _9251_
timestamp 0
transform 1 0 4110 0 -1 730
box -6 -8 66 248
use AND2X2  _9252_
timestamp 0
transform 1 0 3830 0 -1 730
box -6 -8 106 248
use NAND2X1  _9253_
timestamp 0
transform -1 0 4070 0 -1 730
box -6 -8 86 248
use NAND3X1  _9254_
timestamp 0
transform 1 0 3970 0 1 730
box -6 -8 106 248
use NAND2X1  _9255_
timestamp 0
transform -1 0 4210 0 1 730
box -6 -8 86 248
use AOI21X1  _9256_
timestamp 0
transform 1 0 3610 0 -1 1210
box -6 -8 106 248
use AOI21X1  _9257_
timestamp 0
transform -1 0 4010 0 -1 1210
box -6 -8 106 248
use NAND3X1  _9258_
timestamp 0
transform -1 0 4430 0 -1 1210
box -6 -8 106 248
use AOI21X1  _9259_
timestamp 0
transform 1 0 4410 0 1 730
box -6 -8 106 248
use AND2X2  _9260_
timestamp 0
transform 1 0 4270 0 1 730
box -6 -8 106 248
use NAND3X1  _9261_
timestamp 0
transform 1 0 4190 0 -1 1210
box -6 -8 106 248
use OAI21X1  _9262_
timestamp 0
transform 1 0 4570 0 1 730
box -6 -8 106 248
use OAI21X1  _9263_
timestamp 0
transform 1 0 4710 0 1 730
box -6 -8 106 248
use OR2X2  _9264_
timestamp 0
transform 1 0 4870 0 1 730
box -6 -8 106 248
use AOI22X1  _9265_
timestamp 0
transform -1 0 4910 0 1 1690
box -6 -8 126 248
use NAND2X1  _9266_
timestamp 0
transform 1 0 6230 0 1 2170
box -6 -8 86 248
use INVX1  _9267_
timestamp 0
transform -1 0 4290 0 -1 730
box -6 -8 66 248
use NAND2X1  _9268_
timestamp 0
transform 1 0 50 0 -1 2170
box -6 -8 86 248
use INVX1  _9269_
timestamp 0
transform 1 0 310 0 -1 2170
box -6 -8 66 248
use NAND2X1  _9270_
timestamp 0
transform -1 0 370 0 1 1690
box -6 -8 86 248
use NAND2X1  _9271_
timestamp 0
transform -1 0 130 0 1 1690
box -6 -8 86 248
use INVX1  _9272_
timestamp 0
transform -1 0 3650 0 1 250
box -6 -8 66 248
use NAND2X1  _9273_
timestamp 0
transform 1 0 3830 0 1 250
box -6 -8 86 248
use NAND2X1  _9274_
timestamp 0
transform 1 0 3970 0 1 250
box -6 -8 86 248
use NAND2X1  _9275_
timestamp 0
transform 1 0 4090 0 1 250
box -6 -8 86 248
use INVX1  _9276_
timestamp 0
transform -1 0 4290 0 1 250
box -6 -8 66 248
use NOR3X1  _9277_
timestamp 0
transform 1 0 4470 0 -1 730
box -6 -8 186 248
use AOI21X1  _9278_
timestamp 0
transform -1 0 4430 0 -1 730
box -6 -8 106 248
use OAI21X1  _9279_
timestamp 0
transform 1 0 4350 0 1 250
box -6 -8 106 248
use OAI21X1  _9280_
timestamp 0
transform 1 0 4690 0 -1 730
box -6 -8 106 248
use NAND2X1  _9281_
timestamp 0
transform -1 0 6190 0 1 2170
box -6 -8 86 248
use NAND2X1  _9282_
timestamp 0
transform 1 0 3590 0 1 3610
box -6 -8 86 248
use INVX1  _9283_
timestamp 0
transform 1 0 2570 0 -1 4090
box -6 -8 66 248
use NAND2X1  _9284_
timestamp 0
transform 1 0 2930 0 1 3610
box -6 -8 86 248
use OAI21X1  _9285_
timestamp 0
transform 1 0 2490 0 1 3610
box -6 -8 106 248
use NAND2X1  _9286_
timestamp 0
transform 1 0 2010 0 -1 3610
box -6 -8 86 248
use NOR2X1  _9287_
timestamp 0
transform 1 0 1710 0 1 4570
box -6 -8 86 248
use NOR2X1  _9288_
timestamp 0
transform -1 0 650 0 -1 5050
box -6 -8 86 248
use AOI22X1  _9289_
timestamp 0
transform -1 0 1670 0 1 4570
box -6 -8 126 248
use NAND3X1  _9290_
timestamp 0
transform 1 0 1850 0 -1 3610
box -6 -8 106 248
use NAND2X1  _9291_
timestamp 0
transform -1 0 4350 0 1 2170
box -6 -8 86 248
use OAI21X1  _9292_
timestamp 0
transform -1 0 4490 0 1 2170
box -6 -8 106 248
use NAND2X1  _9293_
timestamp 0
transform -1 0 2470 0 1 2650
box -6 -8 86 248
use OAI21X1  _9294_
timestamp 0
transform -1 0 2610 0 1 2650
box -6 -8 106 248
use MUX2X1  _9295_
timestamp 0
transform -1 0 2510 0 1 2170
box -6 -8 126 248
use NAND2X1  _9296_
timestamp 0
transform -1 0 2010 0 1 2650
box -6 -8 86 248
use AND2X2  _9297_
timestamp 0
transform -1 0 2030 0 -1 3130
box -6 -8 106 248
use NOR2X1  _9298_
timestamp 0
transform 1 0 1850 0 1 3610
box -6 -8 86 248
use NAND2X1  _9299_
timestamp 0
transform 1 0 2550 0 1 2170
box -6 -8 86 248
use NAND2X1  _9300_
timestamp 0
transform 1 0 2810 0 1 2170
box -6 -8 86 248
use NAND2X1  _9301_
timestamp 0
transform 1 0 2670 0 1 2170
box -6 -8 86 248
use OAI21X1  _9302_
timestamp 0
transform 1 0 2010 0 -1 2650
box -6 -8 106 248
use OAI21X1  _9303_
timestamp 0
transform 1 0 2350 0 1 3610
box -6 -8 106 248
use OAI21X1  _9304_
timestamp 0
transform 1 0 3210 0 1 3610
box -6 -8 106 248
use NAND2X1  _9305_
timestamp 0
transform -1 0 3950 0 1 3610
box -6 -8 86 248
use NOR2X1  _9306_
timestamp 0
transform -1 0 2290 0 1 3610
box -6 -8 86 248
use NAND2X1  _9307_
timestamp 0
transform 1 0 3290 0 1 3130
box -6 -8 86 248
use OAI21X1  _9308_
timestamp 0
transform 1 0 3130 0 1 3130
box -6 -8 106 248
use NAND2X1  _9309_
timestamp 0
transform 1 0 1450 0 1 4090
box -6 -8 86 248
use OAI21X1  _9310_
timestamp 0
transform 1 0 1310 0 1 4090
box -6 -8 106 248
use MUX2X1  _9311_
timestamp 0
transform -1 0 1930 0 1 3130
box -6 -8 126 248
use NAND2X1  _9312_
timestamp 0
transform 1 0 1890 0 -1 2650
box -6 -8 86 248
use NAND2X1  _9313_
timestamp 0
transform -1 0 3050 0 -1 2170
box -6 -8 86 248
use OAI21X1  _9314_
timestamp 0
transform -1 0 3190 0 -1 2170
box -6 -8 106 248
use INVX1  _9315_
timestamp 0
transform 1 0 1310 0 1 2170
box -6 -8 66 248
use NAND2X1  _9316_
timestamp 0
transform -1 0 2390 0 -1 2650
box -6 -8 86 248
use OAI21X1  _9317_
timestamp 0
transform -1 0 2550 0 -1 2650
box -6 -8 106 248
use NAND2X1  _9318_
timestamp 0
transform -1 0 1650 0 1 2170
box -6 -8 86 248
use OAI21X1  _9319_
timestamp 0
transform 1 0 1430 0 1 2170
box -6 -8 106 248
use OAI21X1  _9320_
timestamp 0
transform 1 0 1730 0 -1 2650
box -6 -8 106 248
use NAND3X1  _9321_
timestamp 0
transform 1 0 1970 0 1 3130
box -6 -8 106 248
use MUX2X1  _9322_
timestamp 0
transform -1 0 2330 0 1 2170
box -6 -8 126 248
use MUX2X1  _9323_
timestamp 0
transform 1 0 2150 0 -1 2650
box -6 -8 126 248
use OAI21X1  _9324_
timestamp 0
transform -1 0 2330 0 1 2650
box -6 -8 106 248
use AOI21X1  _9325_
timestamp 0
transform 1 0 2230 0 1 3130
box -6 -8 106 248
use INVX1  _9326_
timestamp 0
transform 1 0 2410 0 -1 3610
box -6 -8 66 248
use NAND3X1  _9327_
timestamp 0
transform 1 0 2370 0 1 3130
box -6 -8 106 248
use AND2X2  _9328_
timestamp 0
transform 1 0 2510 0 -1 3610
box -6 -8 106 248
use NAND2X1  _9329_
timestamp 0
transform -1 0 2730 0 1 3610
box -6 -8 86 248
use OR2X2  _9330_
timestamp 0
transform 1 0 2770 0 1 3610
box -6 -8 106 248
use AOI21X1  _9331_
timestamp 0
transform 1 0 3070 0 1 3610
box -6 -8 106 248
use OAI21X1  _9332_
timestamp 0
transform 1 0 3710 0 1 3610
box -6 -8 106 248
use NAND2X1  _9333_
timestamp 0
transform 1 0 4070 0 1 3130
box -6 -8 86 248
use AOI21X1  _9334_
timestamp 0
transform 1 0 2530 0 1 3130
box -6 -8 106 248
use NAND2X1  _9335_
timestamp 0
transform -1 0 2250 0 -1 2170
box -6 -8 86 248
use NAND2X1  _9336_
timestamp 0
transform 1 0 2150 0 1 1210
box -6 -8 86 248
use OAI21X1  _9337_
timestamp 0
transform -1 0 2090 0 1 1210
box -6 -8 106 248
use NAND2X1  _9338_
timestamp 0
transform 1 0 2410 0 1 1690
box -6 -8 86 248
use OAI21X1  _9339_
timestamp 0
transform 1 0 1870 0 1 1690
box -6 -8 106 248
use NAND2X1  _9340_
timestamp 0
transform 1 0 1810 0 1 2650
box -6 -8 86 248
use NAND2X1  _9341_
timestamp 0
transform -1 0 1910 0 1 2170
box -6 -8 86 248
use NAND2X1  _9342_
timestamp 0
transform -1 0 1770 0 1 2170
box -6 -8 86 248
use AOI21X1  _9343_
timestamp 0
transform 1 0 1730 0 1 1690
box -6 -8 106 248
use INVX1  _9344_
timestamp 0
transform 1 0 2010 0 1 1690
box -6 -8 66 248
use NAND3X1  _9345_
timestamp 0
transform 1 0 2250 0 1 1690
box -6 -8 106 248
use AOI21X1  _9346_
timestamp 0
transform 1 0 2070 0 1 2650
box -6 -8 106 248
use OAI21X1  _9347_
timestamp 0
transform -1 0 2130 0 -1 2170
box -6 -8 106 248
use NAND3X1  _9348_
timestamp 0
transform 1 0 2310 0 -1 2170
box -6 -8 106 248
use INVX1  _9349_
timestamp 0
transform 1 0 2750 0 -1 2170
box -6 -8 66 248
use AOI21X1  _9350_
timestamp 0
transform 1 0 2470 0 -1 2170
box -6 -8 106 248
use NOR2X1  _9351_
timestamp 0
transform 1 0 2850 0 -1 2170
box -6 -8 86 248
use AND2X2  _9352_
timestamp 0
transform 1 0 3510 0 1 2650
box -6 -8 106 248
use NOR2X1  _9353_
timestamp 0
transform -1 0 3470 0 1 2650
box -6 -8 86 248
use OAI21X1  _9354_
timestamp 0
transform 1 0 3890 0 -1 3130
box -6 -8 106 248
use OAI21X1  _9355_
timestamp 0
transform 1 0 3930 0 1 3130
box -6 -8 106 248
use OAI21X1  _9356_
timestamp 0
transform -1 0 2710 0 -1 2170
box -6 -8 106 248
use INVX1  _9357_
timestamp 0
transform -1 0 2610 0 1 1690
box -6 -8 66 248
use NAND2X1  _9358_
timestamp 0
transform -1 0 2370 0 -1 1210
box -6 -8 86 248
use OAI21X1  _9359_
timestamp 0
transform 1 0 2150 0 -1 1210
box -6 -8 106 248
use MUX2X1  _9360_
timestamp 0
transform -1 0 1230 0 -1 1690
box -6 -8 126 248
use NOR2X1  _9361_
timestamp 0
transform -1 0 1350 0 -1 1690
box -6 -8 86 248
use NAND2X1  _9362_
timestamp 0
transform 1 0 2090 0 -1 3130
box -6 -8 86 248
use NAND2X1  _9363_
timestamp 0
transform -1 0 2030 0 1 2170
box -6 -8 86 248
use NAND2X1  _9364_
timestamp 0
transform -1 0 2150 0 1 2170
box -6 -8 86 248
use OR2X2  _9365_
timestamp 0
transform 1 0 1410 0 -1 1690
box -6 -8 106 248
use OAI21X1  _9366_
timestamp 0
transform -1 0 2210 0 1 1690
box -6 -8 106 248
use OR2X2  _9367_
timestamp 0
transform 1 0 1970 0 -1 1690
box -6 -8 106 248
use OAI21X1  _9368_
timestamp 0
transform 1 0 1810 0 -1 1690
box -6 -8 106 248
use AOI21X1  _9369_
timestamp 0
transform 1 0 2270 0 -1 1690
box -6 -8 106 248
use INVX1  _9370_
timestamp 0
transform 1 0 2550 0 -1 1690
box -6 -8 66 248
use NAND3X1  _9371_
timestamp 0
transform 1 0 2110 0 -1 1690
box -6 -8 106 248
use NAND2X1  _9372_
timestamp 0
transform 1 0 2670 0 -1 1690
box -6 -8 86 248
use OR2X2  _9373_
timestamp 0
transform 1 0 3330 0 1 1690
box -6 -8 106 248
use NAND2X1  _9374_
timestamp 0
transform -1 0 3290 0 1 1690
box -6 -8 86 248
use NAND2X1  _9375_
timestamp 0
transform 1 0 3470 0 1 1690
box -6 -8 86 248
use AOI22X1  _9376_
timestamp 0
transform -1 0 5610 0 -1 2170
box -6 -8 126 248
use AOI21X1  _9377_
timestamp 0
transform -1 0 2510 0 -1 1690
box -6 -8 106 248
use NAND2X1  _9378_
timestamp 0
transform -1 0 250 0 -1 2170
box -6 -8 86 248
use OAI21X1  _9379_
timestamp 0
transform -1 0 950 0 1 1690
box -6 -8 106 248
use NAND2X1  _9380_
timestamp 0
transform -1 0 1510 0 1 1690
box -6 -8 86 248
use OAI21X1  _9381_
timestamp 0
transform -1 0 1670 0 1 1690
box -6 -8 106 248
use NAND2X1  _9382_
timestamp 0
transform -1 0 1390 0 1 1210
box -6 -8 86 248
use OAI21X1  _9383_
timestamp 0
transform -1 0 1530 0 1 1210
box -6 -8 106 248
use INVX1  _9384_
timestamp 0
transform 1 0 1890 0 -1 1210
box -6 -8 66 248
use NAND3X1  _9385_
timestamp 0
transform -1 0 1870 0 -1 2170
box -6 -8 106 248
use OAI21X1  _9386_
timestamp 0
transform -1 0 1830 0 1 1210
box -6 -8 106 248
use OR2X2  _9387_
timestamp 0
transform -1 0 1830 0 -1 1210
box -6 -8 106 248
use NOR2X1  _9388_
timestamp 0
transform -1 0 1670 0 1 1210
box -6 -8 86 248
use OAI21X1  _9389_
timestamp 0
transform -1 0 1550 0 -1 1210
box -6 -8 106 248
use NAND3X1  _9390_
timestamp 0
transform 1 0 1590 0 -1 1210
box -6 -8 106 248
use OR2X2  _9391_
timestamp 0
transform 1 0 2010 0 -1 1210
box -6 -8 106 248
use OAI21X1  _9392_
timestamp 0
transform -1 0 1850 0 1 730
box -6 -8 106 248
use NAND3X1  _9393_
timestamp 0
transform 1 0 2050 0 1 730
box -6 -8 106 248
use NAND2X1  _9394_
timestamp 0
transform -1 0 2530 0 1 730
box -6 -8 86 248
use OR2X2  _9395_
timestamp 0
transform 1 0 2710 0 1 730
box -6 -8 106 248
use NAND2X1  _9396_
timestamp 0
transform 1 0 2590 0 1 730
box -6 -8 86 248
use NAND2X1  _9397_
timestamp 0
transform 1 0 2710 0 -1 1210
box -6 -8 86 248
use AOI22X1  _9398_
timestamp 0
transform -1 0 5790 0 -1 2170
box -6 -8 126 248
use INVX1  _9399_
timestamp 0
transform 1 0 4230 0 -1 1690
box -6 -8 66 248
use OAI21X1  _9400_
timestamp 0
transform 1 0 2590 0 1 250
box -6 -8 106 248
use NAND2X1  _9401_
timestamp 0
transform -1 0 1890 0 -1 730
box -6 -8 86 248
use NOR2X1  _9402_
timestamp 0
transform -1 0 630 0 1 1690
box -6 -8 86 248
use AOI21X1  _9403_
timestamp 0
transform -1 0 1110 0 1 1690
box -6 -8 106 248
use NAND2X1  _9404_
timestamp 0
transform 1 0 1310 0 1 1690
box -6 -8 86 248
use OAI21X1  _9405_
timestamp 0
transform 1 0 1170 0 1 1690
box -6 -8 106 248
use INVX1  _9406_
timestamp 0
transform 1 0 1590 0 -1 730
box -6 -8 66 248
use NAND3X1  _9407_
timestamp 0
transform 1 0 1950 0 -1 730
box -6 -8 106 248
use NOR2X1  _9408_
timestamp 0
transform -1 0 1630 0 -1 1690
box -6 -8 86 248
use NAND3X1  _9409_
timestamp 0
transform 1 0 1670 0 -1 1690
box -6 -8 106 248
use OAI21X1  _9410_
timestamp 0
transform 1 0 1610 0 1 730
box -6 -8 106 248
use NAND2X1  _9411_
timestamp 0
transform -1 0 1770 0 -1 730
box -6 -8 86 248
use AOI21X1  _9412_
timestamp 0
transform -1 0 1970 0 1 250
box -6 -8 106 248
use INVX1  _9413_
timestamp 0
transform -1 0 2230 0 -1 250
box -6 -8 66 248
use NAND3X1  _9414_
timestamp 0
transform 1 0 2010 0 1 250
box -6 -8 106 248
use NAND2X1  _9415_
timestamp 0
transform -1 0 2370 0 -1 250
box -6 -8 86 248
use NOR2X1  _9416_
timestamp 0
transform -1 0 3110 0 1 250
box -6 -8 86 248
use AND2X2  _9417_
timestamp 0
transform 1 0 3170 0 1 250
box -6 -8 106 248
use OAI21X1  _9418_
timestamp 0
transform 1 0 3310 0 1 250
box -6 -8 106 248
use OAI21X1  _9419_
timestamp 0
transform -1 0 3950 0 -1 1690
box -6 -8 106 248
use INVX1  _9420_
timestamp 0
transform -1 0 5450 0 1 2170
box -6 -8 66 248
use NAND3X1  _9421_
timestamp 0
transform -1 0 1550 0 -1 730
box -6 -8 106 248
use AOI21X1  _9422_
timestamp 0
transform -1 0 790 0 1 1690
box -6 -8 106 248
use NAND2X1  _9423_
timestamp 0
transform -1 0 710 0 1 1210
box -6 -8 86 248
use OAI21X1  _9424_
timestamp 0
transform -1 0 1150 0 1 1210
box -6 -8 106 248
use NAND3X1  _9425_
timestamp 0
transform 1 0 1030 0 1 250
box -6 -8 106 248
use NOR3X1  _9426_
timestamp 0
transform -1 0 1550 0 1 730
box -6 -8 186 248
use INVX1  _9427_
timestamp 0
transform 1 0 930 0 1 250
box -6 -8 66 248
use OAI21X1  _9428_
timestamp 0
transform -1 0 1270 0 1 250
box -6 -8 106 248
use NAND2X1  _9429_
timestamp 0
transform -1 0 1410 0 1 250
box -6 -8 86 248
use NAND2X1  _9430_
timestamp 0
transform 1 0 1450 0 1 250
box -6 -8 86 248
use NAND3X1  _9431_
timestamp 0
transform 1 0 1590 0 1 250
box -6 -8 106 248
use NAND2X1  _9432_
timestamp 0
transform 1 0 1730 0 1 250
box -6 -8 86 248
use AOI21X1  _9433_
timestamp 0
transform -1 0 1990 0 1 730
box -6 -8 106 248
use NOR2X1  _9434_
timestamp 0
transform 1 0 2310 0 1 250
box -6 -8 86 248
use OAI21X1  _9435_
timestamp 0
transform -1 0 2530 0 1 250
box -6 -8 106 248
use NAND2X1  _9436_
timestamp 0
transform 1 0 2430 0 -1 250
box -6 -8 86 248
use NOR2X1  _9437_
timestamp 0
transform 1 0 2550 0 -1 250
box -6 -8 86 248
use AND2X2  _9438_
timestamp 0
transform 1 0 2750 0 1 250
box -6 -8 106 248
use AND2X2  _9439_
timestamp 0
transform -1 0 2250 0 1 250
box -6 -8 106 248
use NAND3X1  _9440_
timestamp 0
transform -1 0 2130 0 -1 250
box -6 -8 106 248
use AOI21X1  _9441_
timestamp 0
transform -1 0 1990 0 -1 250
box -6 -8 106 248
use OAI21X1  _9442_
timestamp 0
transform -1 0 1830 0 -1 250
box -6 -8 106 248
use NOR2X1  _9443_
timestamp 0
transform 1 0 2910 0 1 250
box -6 -8 86 248
use OAI21X1  _9444_
timestamp 0
transform 1 0 3690 0 1 250
box -6 -8 106 248
use NAND2X1  _9445_
timestamp 0
transform -1 0 3790 0 -1 1690
box -6 -8 86 248
use OAI21X1  _9446_
timestamp 0
transform -1 0 5350 0 1 2170
box -6 -8 106 248
use INVX1  _9447_
timestamp 0
transform -1 0 3790 0 -1 250
box -6 -8 66 248
use INVX1  _9448_
timestamp 0
transform 1 0 2690 0 -1 250
box -6 -8 66 248
use NAND2X1  _9449_
timestamp 0
transform 1 0 790 0 1 250
box -6 -8 86 248
use NOR2X1  _9450_
timestamp 0
transform -1 0 510 0 1 1690
box -6 -8 86 248
use INVX1  _9451_
timestamp 0
transform 1 0 470 0 -1 1690
box -6 -8 66 248
use OAI21X1  _9452_
timestamp 0
transform -1 0 850 0 1 1210
box -6 -8 106 248
use NAND3X1  _9453_
timestamp 0
transform -1 0 270 0 -1 250
box -6 -8 106 248
use INVX1  _9454_
timestamp 0
transform -1 0 110 0 -1 250
box -6 -8 66 248
use OAI21X1  _9455_
timestamp 0
transform -1 0 1130 0 -1 250
box -6 -8 106 248
use NAND2X1  _9456_
timestamp 0
transform -1 0 690 0 -1 250
box -6 -8 86 248
use NAND3X1  _9457_
timestamp 0
transform 1 0 470 0 -1 250
box -6 -8 106 248
use NAND3X1  _9458_
timestamp 0
transform 1 0 330 0 -1 250
box -6 -8 106 248
use NAND2X1  _9459_
timestamp 0
transform -1 0 810 0 -1 250
box -6 -8 86 248
use NAND3X1  _9460_
timestamp 0
transform 1 0 870 0 -1 250
box -6 -8 106 248
use NAND2X1  _9461_
timestamp 0
transform -1 0 1250 0 -1 250
box -6 -8 86 248
use OAI21X1  _9462_
timestamp 0
transform 1 0 2810 0 -1 250
box -6 -8 106 248
use NOR2X1  _9463_
timestamp 0
transform 1 0 3050 0 -1 250
box -6 -8 86 248
use INVX1  _9464_
timestamp 0
transform 1 0 2950 0 -1 250
box -6 -8 66 248
use AOI21X1  _9465_
timestamp 0
transform 1 0 3190 0 -1 250
box -6 -8 106 248
use AOI22X1  _9466_
timestamp 0
transform -1 0 3450 0 -1 250
box -6 -8 126 248
use OAI21X1  _9467_
timestamp 0
transform -1 0 1410 0 -1 250
box -6 -8 106 248
use NOR2X1  _9468_
timestamp 0
transform -1 0 1690 0 -1 250
box -6 -8 86 248
use AOI21X1  _9469_
timestamp 0
transform -1 0 1570 0 -1 250
box -6 -8 106 248
use INVX1  _9470_
timestamp 0
transform -1 0 770 0 1 730
box -6 -8 66 248
use NAND3X1  _9471_
timestamp 0
transform -1 0 750 0 1 250
box -6 -8 106 248
use INVX1  _9472_
timestamp 0
transform -1 0 1270 0 1 1210
box -6 -8 66 248
use OAI21X1  _9473_
timestamp 0
transform -1 0 990 0 1 1210
box -6 -8 106 248
use INVX1  _9474_
timestamp 0
transform 1 0 930 0 -1 730
box -6 -8 66 248
use NAND3X1  _9475_
timestamp 0
transform 1 0 770 0 -1 730
box -6 -8 106 248
use OAI21X1  _9476_
timestamp 0
transform -1 0 610 0 1 250
box -6 -8 106 248
use NAND2X1  _9477_
timestamp 0
transform 1 0 650 0 -1 730
box -6 -8 86 248
use AOI21X1  _9478_
timestamp 0
transform 1 0 810 0 1 730
box -6 -8 106 248
use NAND3X1  _9479_
timestamp 0
transform 1 0 370 0 1 250
box -6 -8 106 248
use NAND2X1  _9480_
timestamp 0
transform 1 0 1030 0 -1 730
box -6 -8 86 248
use AOI21X1  _9481_
timestamp 0
transform 1 0 1170 0 -1 730
box -6 -8 106 248
use OAI21X1  _9482_
timestamp 0
transform 1 0 2250 0 -1 730
box -6 -8 106 248
use INVX1  _9483_
timestamp 0
transform 1 0 2530 0 -1 730
box -6 -8 66 248
use OR2X2  _9484_
timestamp 0
transform 1 0 2110 0 -1 730
box -6 -8 106 248
use OAI21X1  _9485_
timestamp 0
transform 1 0 2390 0 -1 730
box -6 -8 106 248
use OAI22X1  _9486_
timestamp 0
transform -1 0 3310 0 -1 730
box -6 -8 126 248
use NAND2X1  _9487_
timestamp 0
transform 1 0 3030 0 1 1210
box -6 -8 86 248
use NOR2X1  _9488_
timestamp 0
transform -1 0 2270 0 1 730
box -6 -8 86 248
use NOR2X1  _9489_
timestamp 0
transform 1 0 2330 0 1 730
box -6 -8 86 248
use OAI21X1  _9490_
timestamp 0
transform -1 0 590 0 1 1210
box -6 -8 106 248
use INVX1  _9491_
timestamp 0
transform -1 0 390 0 1 730
box -6 -8 66 248
use OAI21X1  _9492_
timestamp 0
transform 1 0 490 0 -1 730
box -6 -8 106 248
use NAND2X1  _9493_
timestamp 0
transform -1 0 530 0 1 730
box -6 -8 86 248
use OR2X2  _9494_
timestamp 0
transform 1 0 570 0 1 730
box -6 -8 106 248
use NAND3X1  _9495_
timestamp 0
transform 1 0 550 0 -1 1210
box -6 -8 106 248
use NAND2X1  _9496_
timestamp 0
transform -1 0 510 0 -1 1210
box -6 -8 86 248
use NAND2X1  _9497_
timestamp 0
transform -1 0 770 0 -1 1210
box -6 -8 86 248
use NAND2X1  _9498_
timestamp 0
transform 1 0 1330 0 -1 1210
box -6 -8 86 248
use AND2X2  _9499_
timestamp 0
transform 1 0 2410 0 -1 1210
box -6 -8 106 248
use OAI21X1  _9500_
timestamp 0
transform 1 0 2570 0 -1 1210
box -6 -8 106 248
use OAI21X1  _9501_
timestamp 0
transform 1 0 2650 0 1 1210
box -6 -8 106 248
use INVX1  _9502_
timestamp 0
transform 1 0 5130 0 -1 2650
box -6 -8 66 248
use INVX1  _9503_
timestamp 0
transform 1 0 970 0 -1 1210
box -6 -8 66 248
use AOI21X1  _9504_
timestamp 0
transform 1 0 950 0 1 730
box -6 -8 106 248
use NOR2X1  _9505_
timestamp 0
transform 1 0 1330 0 -1 730
box -6 -8 86 248
use NAND3X1  _9506_
timestamp 0
transform -1 0 1330 0 1 730
box -6 -8 106 248
use OAI21X1  _9507_
timestamp 0
transform -1 0 1190 0 1 730
box -6 -8 106 248
use OAI21X1  _9508_
timestamp 0
transform -1 0 450 0 1 1210
box -6 -8 106 248
use INVX1  _9509_
timestamp 0
transform 1 0 310 0 -1 1210
box -6 -8 66 248
use OR2X2  _9510_
timestamp 0
transform -1 0 310 0 1 250
box -6 -8 106 248
use OAI21X1  _9511_
timestamp 0
transform -1 0 150 0 1 250
box -6 -8 106 248
use NAND2X1  _9512_
timestamp 0
transform 1 0 370 0 -1 730
box -6 -8 86 248
use OR2X2  _9513_
timestamp 0
transform -1 0 150 0 -1 730
box -6 -8 106 248
use NAND3X1  _9514_
timestamp 0
transform -1 0 150 0 1 730
box -6 -8 106 248
use AND2X2  _9515_
timestamp 0
transform 1 0 210 0 -1 730
box -6 -8 106 248
use NOR2X1  _9516_
timestamp 0
transform 1 0 190 0 1 730
box -6 -8 86 248
use OAI21X1  _9517_
timestamp 0
transform 1 0 190 0 1 1210
box -6 -8 106 248
use NAND2X1  _9518_
timestamp 0
transform -1 0 130 0 1 1210
box -6 -8 86 248
use AND2X2  _9519_
timestamp 0
transform -1 0 170 0 -1 1690
box -6 -8 106 248
use NOR2X1  _9520_
timestamp 0
transform 1 0 210 0 -1 1690
box -6 -8 86 248
use NOR2X1  _9521_
timestamp 0
transform 1 0 170 0 1 1690
box -6 -8 86 248
use AOI22X1  _9522_
timestamp 0
transform -1 0 5090 0 -1 2650
box -6 -8 126 248
use NAND2X1  _9523_
timestamp 0
transform -1 0 3290 0 -1 1210
box -6 -8 86 248
use INVX1  _9524_
timestamp 0
transform 1 0 70 0 -1 1210
box -6 -8 66 248
use AOI21X1  _9525_
timestamp 0
transform 1 0 170 0 -1 1210
box -6 -8 106 248
use NAND2X1  _9526_
timestamp 0
transform 1 0 2630 0 -1 730
box -6 -8 86 248
use NOR2X1  _9527_
timestamp 0
transform -1 0 2850 0 -1 730
box -6 -8 86 248
use AOI21X1  _9528_
timestamp 0
transform 1 0 3030 0 -1 730
box -6 -8 106 248
use NOR2X1  _9529_
timestamp 0
transform -1 0 2990 0 -1 730
box -6 -8 86 248
use AND2X2  _9530_
timestamp 0
transform 1 0 2850 0 1 730
box -6 -8 106 248
use OAI21X1  _9531_
timestamp 0
transform 1 0 3010 0 1 730
box -6 -8 106 248
use OAI21X1  _9532_
timestamp 0
transform 1 0 3150 0 1 730
box -6 -8 106 248
use OAI21X1  _9533_
timestamp 0
transform 1 0 770 0 -1 5530
box -6 -8 106 248
use OAI21X1  _9534_
timestamp 0
transform 1 0 1450 0 -1 6010
box -6 -8 106 248
use INVX1  _9535_
timestamp 0
transform 1 0 1590 0 1 6010
box -6 -8 66 248
use NOR2X1  _9536_
timestamp 0
transform 1 0 1310 0 -1 6010
box -6 -8 86 248
use NAND2X1  _9537_
timestamp 0
transform -1 0 1670 0 -1 6010
box -6 -8 86 248
use NAND2X1  _9538_
timestamp 0
transform 1 0 1710 0 -1 6010
box -6 -8 86 248
use NAND2X1  _9539_
timestamp 0
transform 1 0 3650 0 -1 6010
box -6 -8 86 248
use OAI21X1  _9540_
timestamp 0
transform 1 0 3250 0 -1 6010
box -6 -8 106 248
use NAND2X1  _9541_
timestamp 0
transform 1 0 2110 0 -1 6490
box -6 -8 86 248
use INVX1  _9542_
timestamp 0
transform -1 0 1550 0 1 6010
box -6 -8 66 248
use NOR2X1  _9543_
timestamp 0
transform 1 0 1290 0 1 6490
box -6 -8 86 248
use AOI21X1  _9544_
timestamp 0
transform -1 0 1270 0 -1 6490
box -6 -8 106 248
use NOR2X1  _9545_
timestamp 0
transform 1 0 990 0 1 6010
box -6 -8 86 248
use OAI21X1  _9546_
timestamp 0
transform 1 0 850 0 -1 6010
box -6 -8 106 248
use AND2X2  _9547_
timestamp 0
transform -1 0 950 0 1 6010
box -6 -8 106 248
use OR2X2  _9548_
timestamp 0
transform 1 0 890 0 -1 6490
box -6 -8 106 248
use OR2X2  _9549_
timestamp 0
transform -1 0 490 0 1 6490
box -6 -8 106 248
use OAI21X1  _9550_
timestamp 0
transform -1 0 830 0 -1 6490
box -6 -8 106 248
use NAND2X1  _9551_
timestamp 0
transform -1 0 610 0 1 6490
box -6 -8 86 248
use NOR2X1  _9552_
timestamp 0
transform -1 0 1530 0 -1 6490
box -6 -8 86 248
use NAND2X1  _9553_
timestamp 0
transform -1 0 1410 0 -1 6490
box -6 -8 86 248
use NAND2X1  _9554_
timestamp 0
transform -1 0 1650 0 -1 6490
box -6 -8 86 248
use OAI21X1  _9555_
timestamp 0
transform 1 0 1710 0 -1 6490
box -6 -8 106 248
use INVX1  _9556_
timestamp 0
transform 1 0 650 0 1 6490
box -6 -8 66 248
use OAI21X1  _9557_
timestamp 0
transform 1 0 1030 0 -1 6490
box -6 -8 106 248
use OAI21X1  _9558_
timestamp 0
transform 1 0 190 0 -1 5530
box -6 -8 106 248
use OAI21X1  _9559_
timestamp 0
transform 1 0 50 0 1 5530
box -6 -8 106 248
use MUX2X1  _9560_
timestamp 0
transform -1 0 330 0 1 5530
box -6 -8 126 248
use NAND2X1  _9561_
timestamp 0
transform -1 0 290 0 -1 6010
box -6 -8 86 248
use OR2X2  _9562_
timestamp 0
transform -1 0 170 0 -1 6010
box -6 -8 106 248
use NAND2X1  _9563_
timestamp 0
transform -1 0 130 0 1 6010
box -6 -8 86 248
use INVX1  _9564_
timestamp 0
transform -1 0 110 0 -1 6490
box -6 -8 66 248
use NOR2X1  _9565_
timestamp 0
transform 1 0 290 0 -1 6490
box -6 -8 86 248
use NAND2X1  _9566_
timestamp 0
transform -1 0 230 0 -1 6490
box -6 -8 86 248
use NAND2X1  _9567_
timestamp 0
transform -1 0 670 0 -1 6490
box -6 -8 86 248
use OAI22X1  _9568_
timestamp 0
transform -1 0 530 0 -1 6490
box -6 -8 126 248
use NOR2X1  _9569_
timestamp 0
transform -1 0 2170 0 1 6010
box -6 -8 86 248
use NAND2X1  _9570_
timestamp 0
transform -1 0 270 0 1 6010
box -6 -8 86 248
use INVX1  _9571_
timestamp 0
transform 1 0 310 0 1 6010
box -6 -8 66 248
use INVX1  _9572_
timestamp 0
transform -1 0 990 0 1 5530
box -6 -8 66 248
use NOR2X1  _9573_
timestamp 0
transform -1 0 130 0 -1 5530
box -6 -8 86 248
use OAI21X1  _9574_
timestamp 0
transform 1 0 490 0 -1 5530
box -6 -8 106 248
use OAI21X1  _9575_
timestamp 0
transform -1 0 690 0 1 5050
box -6 -8 106 248
use OAI21X1  _9576_
timestamp 0
transform -1 0 730 0 -1 5530
box -6 -8 106 248
use NOR2X1  _9577_
timestamp 0
transform 1 0 670 0 1 5530
box -6 -8 86 248
use NAND2X1  _9578_
timestamp 0
transform 1 0 790 0 1 5530
box -6 -8 86 248
use INVX1  _9579_
timestamp 0
transform -1 0 790 0 -1 6010
box -6 -8 66 248
use NOR2X1  _9580_
timestamp 0
transform -1 0 670 0 -1 6010
box -6 -8 86 248
use OAI21X1  _9581_
timestamp 0
transform -1 0 530 0 1 6010
box -6 -8 106 248
use AOI21X1  _9582_
timestamp 0
transform 1 0 570 0 1 6010
box -6 -8 106 248
use NOR2X1  _9583_
timestamp 0
transform -1 0 2050 0 1 6010
box -6 -8 86 248
use NAND2X1  _9584_
timestamp 0
transform 1 0 4370 0 1 5530
box -6 -8 86 248
use INVX1  _9585_
timestamp 0
transform 1 0 3090 0 1 6010
box -6 -8 66 248
use AOI21X1  _9586_
timestamp 0
transform 1 0 1010 0 -1 6010
box -6 -8 106 248
use OAI21X1  _9587_
timestamp 0
transform -1 0 1250 0 -1 6010
box -6 -8 106 248
use OAI21X1  _9588_
timestamp 0
transform 1 0 1110 0 1 6010
box -6 -8 106 248
use OR2X2  _9589_
timestamp 0
transform 1 0 3210 0 1 6010
box -6 -8 106 248
use NAND2X1  _9590_
timestamp 0
transform 1 0 3350 0 1 6010
box -6 -8 86 248
use NAND2X1  _9591_
timestamp 0
transform 1 0 3490 0 1 6010
box -6 -8 86 248
use AOI21X1  _9592_
timestamp 0
transform 1 0 710 0 1 6010
box -6 -8 106 248
use AND2X2  _9593_
timestamp 0
transform 1 0 3890 0 1 6010
box -6 -8 106 248
use OAI21X1  _9594_
timestamp 0
transform -1 0 3830 0 1 6010
box -6 -8 106 248
use OAI21X1  _9595_
timestamp 0
transform 1 0 3770 0 -1 6010
box -6 -8 106 248
use OAI21X1  _9596_
timestamp 0
transform -1 0 3810 0 -1 6490
box -6 -8 106 248
use INVX1  _9597_
timestamp 0
transform -1 0 2470 0 1 6490
box -6 -8 66 248
use OAI21X1  _9598_
timestamp 0
transform -1 0 1610 0 -1 5050
box -6 -8 106 248
use OAI21X1  _9599_
timestamp 0
transform -1 0 1250 0 -1 5530
box -6 -8 106 248
use OR2X2  _9600_
timestamp 0
transform 1 0 1390 0 -1 5530
box -6 -8 106 248
use NAND2X1  _9601_
timestamp 0
transform 1 0 1550 0 -1 5530
box -6 -8 86 248
use OR2X2  _9602_
timestamp 0
transform 1 0 2890 0 1 6490
box -6 -8 106 248
use NAND2X1  _9603_
timestamp 0
transform -1 0 2850 0 1 6490
box -6 -8 86 248
use NAND2X1  _9604_
timestamp 0
transform -1 0 3110 0 1 6490
box -6 -8 86 248
use INVX1  _9605_
timestamp 0
transform 1 0 3310 0 1 6490
box -6 -8 66 248
use NOR2X1  _9606_
timestamp 0
transform 1 0 3890 0 1 6490
box -6 -8 86 248
use NAND2X1  _9607_
timestamp 0
transform -1 0 3850 0 1 6490
box -6 -8 86 248
use NAND2X1  _9608_
timestamp 0
transform -1 0 4770 0 -1 6490
box -6 -8 86 248
use OAI22X1  _9609_
timestamp 0
transform -1 0 4930 0 -1 6490
box -6 -8 126 248
use NAND2X1  _9610_
timestamp 0
transform -1 0 4570 0 -1 6010
box -6 -8 86 248
use INVX1  _9611_
timestamp 0
transform -1 0 3650 0 -1 6490
box -6 -8 66 248
use NAND2X1  _9612_
timestamp 0
transform -1 0 3950 0 -1 6490
box -6 -8 86 248
use OAI21X1  _9613_
timestamp 0
transform -1 0 3250 0 1 6490
box -6 -8 106 248
use INVX1  _9614_
timestamp 0
transform 1 0 3410 0 1 6490
box -6 -8 66 248
use OAI21X1  _9615_
timestamp 0
transform 1 0 4010 0 -1 6490
box -6 -8 106 248
use OAI21X1  _9616_
timestamp 0
transform 1 0 330 0 -1 5530
box -6 -8 106 248
use NOR2X1  _9617_
timestamp 0
transform 1 0 390 0 1 5530
box -6 -8 86 248
use NAND2X1  _9618_
timestamp 0
transform 1 0 330 0 -1 6010
box -6 -8 86 248
use OAI21X1  _9619_
timestamp 0
transform 1 0 510 0 1 5530
box -6 -8 106 248
use NAND2X1  _9620_
timestamp 0
transform -1 0 550 0 -1 6010
box -6 -8 86 248
use NAND2X1  _9621_
timestamp 0
transform -1 0 2530 0 1 6010
box -6 -8 86 248
use OR2X2  _9622_
timestamp 0
transform 1 0 2490 0 -1 6490
box -6 -8 106 248
use NAND2X1  _9623_
timestamp 0
transform -1 0 2850 0 -1 6490
box -6 -8 86 248
use INVX1  _9624_
timestamp 0
transform 1 0 3030 0 -1 6490
box -6 -8 66 248
use NOR2X1  _9625_
timestamp 0
transform 1 0 4270 0 -1 6490
box -6 -8 86 248
use NAND2X1  _9626_
timestamp 0
transform -1 0 4230 0 -1 6490
box -6 -8 86 248
use NAND2X1  _9627_
timestamp 0
transform -1 0 4630 0 -1 6490
box -6 -8 86 248
use OAI21X1  _9628_
timestamp 0
transform 1 0 4390 0 -1 6490
box -6 -8 106 248
use INVX1  _9629_
timestamp 0
transform -1 0 4690 0 -1 6010
box -6 -8 66 248
use NAND2X1  _9630_
timestamp 0
transform 1 0 4030 0 1 6010
box -6 -8 86 248
use INVX1  _9631_
timestamp 0
transform -1 0 2370 0 1 6490
box -6 -8 66 248
use NAND2X1  _9632_
timestamp 0
transform 1 0 1410 0 1 6490
box -6 -8 86 248
use OR2X2  _9633_
timestamp 0
transform 1 0 1530 0 1 6490
box -6 -8 106 248
use NAND2X1  _9634_
timestamp 0
transform -1 0 1770 0 1 6490
box -6 -8 86 248
use NOR2X1  _9635_
timestamp 0
transform -1 0 2130 0 1 6490
box -6 -8 86 248
use INVX1  _9636_
timestamp 0
transform 1 0 2250 0 -1 6490
box -6 -8 66 248
use NAND2X1  _9637_
timestamp 0
transform -1 0 2250 0 1 6490
box -6 -8 86 248
use NAND2X1  _9638_
timestamp 0
transform 1 0 2350 0 -1 6490
box -6 -8 86 248
use OR2X2  _9639_
timestamp 0
transform 1 0 4170 0 1 6010
box -6 -8 106 248
use AOI21X1  _9640_
timestamp 0
transform 1 0 4150 0 -1 6010
box -6 -8 106 248
use AOI22X1  _9641_
timestamp 0
transform -1 0 4430 0 -1 6010
box -6 -8 126 248
use NAND2X1  _9642_
timestamp 0
transform 1 0 3930 0 -1 5530
box -6 -8 86 248
use NOR2X1  _9643_
timestamp 0
transform -1 0 1450 0 -1 5050
box -6 -8 86 248
use INVX1  _9644_
timestamp 0
transform 1 0 1650 0 1 5050
box -6 -8 66 248
use NAND3X1  _9645_
timestamp 0
transform 1 0 1970 0 -1 5530
box -6 -8 106 248
use INVX1  _9646_
timestamp 0
transform 1 0 2850 0 1 5530
box -6 -8 66 248
use AOI21X1  _9647_
timestamp 0
transform 1 0 1970 0 1 5530
box -6 -8 106 248
use NOR2X1  _9648_
timestamp 0
transform 1 0 2710 0 1 5530
box -6 -8 86 248
use OAI21X1  _9649_
timestamp 0
transform -1 0 2730 0 -1 6490
box -6 -8 106 248
use NOR2X1  _9650_
timestamp 0
transform -1 0 2970 0 -1 6490
box -6 -8 86 248
use AOI21X1  _9651_
timestamp 0
transform 1 0 3150 0 -1 6490
box -6 -8 106 248
use NAND3X1  _9652_
timestamp 0
transform -1 0 3550 0 -1 6490
box -6 -8 106 248
use OAI21X1  _9653_
timestamp 0
transform -1 0 3410 0 -1 6490
box -6 -8 106 248
use NOR2X1  _9654_
timestamp 0
transform -1 0 3390 0 -1 5530
box -6 -8 86 248
use NAND2X1  _9655_
timestamp 0
transform -1 0 3370 0 1 5530
box -6 -8 86 248
use NAND2X1  _9656_
timestamp 0
transform -1 0 3510 0 -1 5530
box -6 -8 86 248
use OAI21X1  _9657_
timestamp 0
transform 1 0 3550 0 -1 5530
box -6 -8 106 248
use AOI21X1  _9658_
timestamp 0
transform -1 0 3070 0 1 5530
box -6 -8 106 248
use OR2X2  _9659_
timestamp 0
transform 1 0 2130 0 1 5050
box -6 -8 106 248
use NAND2X1  _9660_
timestamp 0
transform -1 0 2090 0 1 5050
box -6 -8 86 248
use NAND2X1  _9661_
timestamp 0
transform -1 0 2470 0 1 5050
box -6 -8 86 248
use AND2X2  _9662_
timestamp 0
transform -1 0 2970 0 -1 5530
box -6 -8 106 248
use OAI21X1  _9663_
timestamp 0
transform 1 0 3010 0 -1 5530
box -6 -8 106 248
use OAI22X1  _9664_
timestamp 0
transform -1 0 3270 0 -1 5530
box -6 -8 126 248
use NAND2X1  _9665_
timestamp 0
transform -1 0 3730 0 1 5050
box -6 -8 86 248
use OAI21X1  _9666_
timestamp 0
transform -1 0 2670 0 -1 5530
box -6 -8 106 248
use NAND3X1  _9667_
timestamp 0
transform 1 0 2430 0 -1 5530
box -6 -8 106 248
use INVX1  _9668_
timestamp 0
transform 1 0 2590 0 1 5530
box -6 -8 66 248
use AOI21X1  _9669_
timestamp 0
transform -1 0 2810 0 -1 5530
box -6 -8 106 248
use INVX1  _9670_
timestamp 0
transform 1 0 2710 0 -1 5050
box -6 -8 66 248
use NAND2X1  _9671_
timestamp 0
transform -1 0 2890 0 1 5050
box -6 -8 86 248
use NAND2X1  _9672_
timestamp 0
transform 1 0 2690 0 1 5050
box -6 -8 86 248
use NAND2X1  _9673_
timestamp 0
transform 1 0 2930 0 1 5050
box -6 -8 86 248
use AND2X2  _9674_
timestamp 0
transform 1 0 3210 0 1 5050
box -6 -8 106 248
use OAI21X1  _9675_
timestamp 0
transform 1 0 3350 0 1 5050
box -6 -8 106 248
use OAI21X1  _9676_
timestamp 0
transform 1 0 3490 0 1 5050
box -6 -8 106 248
use NAND2X1  _9677_
timestamp 0
transform -1 0 4270 0 1 5050
box -6 -8 86 248
use OAI21X1  _9678_
timestamp 0
transform -1 0 3150 0 1 5050
box -6 -8 106 248
use OAI21X1  _9679_
timestamp 0
transform 1 0 4030 0 1 5050
box -6 -8 106 248
use NAND2X1  _9680_
timestamp 0
transform -1 0 3090 0 1 4090
box -6 -8 86 248
use NAND2X1  _9681_
timestamp 0
transform -1 0 3690 0 1 4090
box -6 -8 86 248
use NOR2X1  _9682_
timestamp 0
transform -1 0 2970 0 1 4090
box -6 -8 86 248
use NAND2X1  _9683_
timestamp 0
transform -1 0 270 0 -1 3610
box -6 -8 86 248
use OAI21X1  _9684_
timestamp 0
transform -1 0 410 0 -1 3130
box -6 -8 106 248
use NAND2X1  _9685_
timestamp 0
transform -1 0 130 0 1 3130
box -6 -8 86 248
use OAI21X1  _9686_
timestamp 0
transform -1 0 170 0 1 2650
box -6 -8 106 248
use INVX1  _9687_
timestamp 0
transform -1 0 270 0 1 4570
box -6 -8 66 248
use OR2X2  _9688_
timestamp 0
transform -1 0 550 0 1 5050
box -6 -8 106 248
use OAI21X1  _9689_
timestamp 0
transform 1 0 730 0 1 4570
box -6 -8 106 248
use OAI21X1  _9690_
timestamp 0
transform -1 0 970 0 1 4570
box -6 -8 106 248
use INVX1  _9691_
timestamp 0
transform -1 0 130 0 -1 5050
box -6 -8 66 248
use OAI21X1  _9692_
timestamp 0
transform -1 0 550 0 -1 4570
box -6 -8 106 248
use OAI21X1  _9693_
timestamp 0
transform -1 0 430 0 1 4570
box -6 -8 106 248
use NAND2X1  _9694_
timestamp 0
transform 1 0 4370 0 1 4570
box -6 -8 86 248
use NAND2X1  _9695_
timestamp 0
transform -1 0 130 0 -1 4570
box -6 -8 86 248
use OAI21X1  _9696_
timestamp 0
transform -1 0 170 0 1 4570
box -6 -8 106 248
use NAND2X1  _9697_
timestamp 0
transform -1 0 250 0 -1 4570
box -6 -8 86 248
use OAI21X1  _9698_
timestamp 0
transform -1 0 410 0 -1 4570
box -6 -8 106 248
use AND2X2  _9699_
timestamp 0
transform -1 0 3770 0 -1 5050
box -6 -8 106 248
use NAND2X1  _9700_
timestamp 0
transform 1 0 1430 0 -1 3610
box -6 -8 86 248
use OAI21X1  _9701_
timestamp 0
transform 1 0 1290 0 -1 3610
box -6 -8 106 248
use NAND2X1  _9702_
timestamp 0
transform 1 0 1370 0 1 3130
box -6 -8 86 248
use OAI21X1  _9703_
timestamp 0
transform -1 0 1890 0 -1 3130
box -6 -8 106 248
use OAI21X1  _9704_
timestamp 0
transform 1 0 1170 0 1 4570
box -6 -8 106 248
use OAI21X1  _9705_
timestamp 0
transform 1 0 1030 0 1 4570
box -6 -8 106 248
use OAI21X1  _9706_
timestamp 0
transform -1 0 790 0 -1 5050
box -6 -8 106 248
use OAI21X1  _9707_
timestamp 0
transform 1 0 410 0 -1 5050
box -6 -8 106 248
use NAND2X1  _9708_
timestamp 0
transform -1 0 1930 0 -1 4570
box -6 -8 86 248
use OAI21X1  _9709_
timestamp 0
transform -1 0 1790 0 -1 4570
box -6 -8 106 248
use NAND2X1  _9710_
timestamp 0
transform -1 0 1010 0 1 4090
box -6 -8 86 248
use OAI21X1  _9711_
timestamp 0
transform -1 0 1150 0 1 4090
box -6 -8 106 248
use NAND2X1  _9712_
timestamp 0
transform -1 0 2970 0 1 3130
box -6 -8 86 248
use OAI21X1  _9713_
timestamp 0
transform -1 0 3050 0 1 2170
box -6 -8 106 248
use NAND2X1  _9714_
timestamp 0
transform -1 0 370 0 1 3130
box -6 -8 86 248
use OAI21X1  _9715_
timestamp 0
transform -1 0 410 0 1 2170
box -6 -8 106 248
use INVX1  _9716_
timestamp 0
transform -1 0 2410 0 1 4570
box -6 -8 66 248
use OAI21X1  _9717_
timestamp 0
transform 1 0 2050 0 -1 5050
box -6 -8 106 248
use OAI21X1  _9718_
timestamp 0
transform -1 0 1990 0 -1 5050
box -6 -8 106 248
use INVX1  _9719_
timestamp 0
transform -1 0 3430 0 1 4570
box -6 -8 66 248
use OAI21X1  _9720_
timestamp 0
transform 1 0 3630 0 1 4570
box -6 -8 106 248
use OAI21X1  _9721_
timestamp 0
transform 1 0 3470 0 1 4570
box -6 -8 106 248
use NAND2X1  _9722_
timestamp 0
transform 1 0 2370 0 -1 4570
box -6 -8 86 248
use OAI21X1  _9723_
timestamp 0
transform 1 0 2210 0 -1 4570
box -6 -8 106 248
use NAND2X1  _9724_
timestamp 0
transform -1 0 3130 0 -1 4570
box -6 -8 86 248
use OAI21X1  _9725_
timestamp 0
transform -1 0 3270 0 -1 4570
box -6 -8 106 248
use NAND2X1  _9726_
timestamp 0
transform 1 0 3010 0 1 3130
box -6 -8 86 248
use OAI21X1  _9727_
timestamp 0
transform -1 0 3530 0 1 3130
box -6 -8 106 248
use NAND2X1  _9728_
timestamp 0
transform -1 0 2190 0 1 3130
box -6 -8 86 248
use OAI21X1  _9729_
timestamp 0
transform -1 0 2570 0 -1 3130
box -6 -8 106 248
use OAI21X1  _9730_
timestamp 0
transform 1 0 2210 0 1 4570
box -6 -8 106 248
use OAI21X1  _9731_
timestamp 0
transform 1 0 2070 0 1 4570
box -6 -8 106 248
use OAI21X1  _9732_
timestamp 0
transform -1 0 2950 0 1 4570
box -6 -8 106 248
use OAI21X1  _9733_
timestamp 0
transform -1 0 3330 0 1 4570
box -6 -8 106 248
use NAND2X1  _9734_
timestamp 0
transform -1 0 2590 0 -1 4570
box -6 -8 86 248
use OAI21X1  _9735_
timestamp 0
transform 1 0 2630 0 -1 4570
box -6 -8 106 248
use NAND2X1  _9736_
timestamp 0
transform -1 0 930 0 -1 5050
box -6 -8 86 248
use OAI21X1  _9737_
timestamp 0
transform -1 0 1070 0 -1 5050
box -6 -8 106 248
use NAND2X1  _9738_
timestamp 0
transform -1 0 2350 0 1 5050
box -6 -8 86 248
use OAI21X1  _9739_
timestamp 0
transform -1 0 2630 0 1 5050
box -6 -8 106 248
use NAND2X1  _9740_
timestamp 0
transform 1 0 1270 0 1 5050
box -6 -8 86 248
use OAI21X1  _9741_
timestamp 0
transform 1 0 1130 0 1 5050
box -6 -8 106 248
use INVX1  _9742_
timestamp 0
transform -1 0 1890 0 -1 6010
box -6 -8 66 248
use OAI21X1  _9743_
timestamp 0
transform 1 0 1690 0 -1 5530
box -6 -8 106 248
use OAI21X1  _9744_
timestamp 0
transform -1 0 1930 0 -1 5530
box -6 -8 106 248
use INVX1  _9745_
timestamp 0
transform 1 0 1290 0 -1 5530
box -6 -8 66 248
use OAI21X1  _9746_
timestamp 0
transform 1 0 2130 0 -1 5530
box -6 -8 106 248
use OAI21X1  _9747_
timestamp 0
transform -1 0 2370 0 -1 5530
box -6 -8 106 248
use NAND2X1  _9748_
timestamp 0
transform -1 0 2410 0 -1 6010
box -6 -8 86 248
use OAI21X1  _9749_
timestamp 0
transform 1 0 2170 0 -1 6010
box -6 -8 106 248
use NAND2X1  _9750_
timestamp 0
transform 1 0 2610 0 -1 6010
box -6 -8 86 248
use OAI21X1  _9751_
timestamp 0
transform 1 0 2470 0 -1 6010
box -6 -8 106 248
use NAND2X1  _9752_
timestamp 0
transform -1 0 2650 0 1 6010
box -6 -8 86 248
use OAI21X1  _9753_
timestamp 0
transform -1 0 2810 0 1 6010
box -6 -8 106 248
use NAND2X1  _9754_
timestamp 0
transform 1 0 3130 0 -1 6010
box -6 -8 86 248
use OAI21X1  _9755_
timestamp 0
transform 1 0 2990 0 -1 6010
box -6 -8 106 248
use OAI21X1  _9756_
timestamp 0
transform 1 0 1330 0 1 5530
box -6 -8 106 248
use OAI21X1  _9757_
timestamp 0
transform -1 0 1810 0 1 5530
box -6 -8 106 248
use OAI21X1  _9758_
timestamp 0
transform -1 0 1150 0 1 5530
box -6 -8 106 248
use OAI21X1  _9759_
timestamp 0
transform -1 0 1290 0 1 5530
box -6 -8 106 248
use NAND2X1  _9760_
timestamp 0
transform 1 0 1850 0 1 6010
box -6 -8 86 248
use OAI21X1  _9761_
timestamp 0
transform 1 0 1690 0 1 6010
box -6 -8 106 248
use NAND2X1  _9762_
timestamp 0
transform 1 0 1150 0 1 6490
box -6 -8 86 248
use OAI21X1  _9763_
timestamp 0
transform -1 0 1110 0 1 6490
box -6 -8 106 248
use DFFPOSX1  _9764_
timestamp 0
transform 1 0 3650 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _9765_
timestamp 0
transform 1 0 4310 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _9766_
timestamp 0
transform 1 0 7250 0 1 6490
box -6 -8 246 248
use DFFPOSX1  _9767_
timestamp 0
transform 1 0 3690 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _9768_
timestamp 0
transform -1 0 5190 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _9769_
timestamp 0
transform 1 0 5970 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _9770_
timestamp 0
transform 1 0 4710 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _9771_
timestamp 0
transform -1 0 6630 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _9772_
timestamp 0
transform 1 0 4650 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _9773_
timestamp 0
transform 1 0 5270 0 -1 1690
box -6 -8 246 248
use DFFPOSX1  _9774_
timestamp 0
transform -1 0 5370 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _9775_
timestamp 0
transform 1 0 4910 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _9776_
timestamp 0
transform -1 0 6550 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _9777_
timestamp 0
transform 1 0 3310 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _9778_
timestamp 0
transform 1 0 3710 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _9779_
timestamp 0
transform -1 0 4390 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _9780_
timestamp 0
transform 1 0 5690 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _9781_
timestamp 0
transform -1 0 6130 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _9782_
timestamp 0
transform 1 0 3950 0 -1 1690
box -6 -8 246 248
use DFFPOSX1  _9783_
timestamp 0
transform 1 0 5450 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _9784_
timestamp 0
transform 1 0 3450 0 -1 250
box -6 -8 246 248
use DFFPOSX1  _9785_
timestamp 0
transform 1 0 3310 0 -1 730
box -6 -8 246 248
use DFFPOSX1  _9786_
timestamp 0
transform 1 0 2750 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _9787_
timestamp 0
transform -1 0 5430 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _9788_
timestamp 0
transform 1 0 2930 0 -1 1210
box -6 -8 246 248
use DFFPOSX1  _9789_
timestamp 0
transform 1 0 3350 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _9790_
timestamp 0
transform 1 0 1810 0 -1 6490
box -6 -8 246 248
use DFFPOSX1  _9791_
timestamp 0
transform 1 0 10 0 1 6490
box -6 -8 246 248
use DFFPOSX1  _9792_
timestamp 0
transform 1 0 1890 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _9793_
timestamp 0
transform 1 0 3870 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _9794_
timestamp 0
transform 1 0 4630 0 1 6010
box -6 -8 246 248
use DFFPOSX1  _9795_
timestamp 0
transform 1 0 4270 0 1 6010
box -6 -8 246 248
use DFFPOSX1  _9796_
timestamp 0
transform -1 0 4930 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _9797_
timestamp 0
transform 1 0 3650 0 -1 5530
box -6 -8 246 248
use DFFPOSX1  _9798_
timestamp 0
transform 1 0 3370 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _9799_
timestamp 0
transform 1 0 3730 0 1 5050
box -6 -8 246 248
use DFFPOSX1  _9800_
timestamp 0
transform -1 0 4510 0 1 5050
box -6 -8 246 248
use DFFPOSX1  _9801_
timestamp 0
transform 1 0 10 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _9802_
timestamp 0
transform 1 0 10 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _9803_
timestamp 0
transform 1 0 790 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _9804_
timestamp 0
transform -1 0 670 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _9805_
timestamp 0
transform 1 0 10 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _9806_
timestamp 0
transform -1 0 790 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _9807_
timestamp 0
transform -1 0 1230 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _9808_
timestamp 0
transform -1 0 2410 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _9809_
timestamp 0
transform 1 0 1030 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _9810_
timestamp 0
transform 1 0 130 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _9811_
timestamp 0
transform -1 0 1510 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _9812_
timestamp 0
transform 1 0 1170 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _9813_
timestamp 0
transform 1 0 3050 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _9814_
timestamp 0
transform -1 0 250 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _9815_
timestamp 0
transform 1 0 1610 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _9816_
timestamp 0
transform 1 0 3730 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _9817_
timestamp 0
transform 1 0 1930 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _9818_
timestamp 0
transform 1 0 3270 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _9819_
timestamp 0
transform -1 0 3870 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _9820_
timestamp 0
transform 1 0 2570 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _9821_
timestamp 0
transform -1 0 2030 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _9822_
timestamp 0
transform -1 0 3190 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _9823_
timestamp 0
transform -1 0 2790 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _9824_
timestamp 0
transform 1 0 1070 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _9825_
timestamp 0
transform 1 0 2410 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _9826_
timestamp 0
transform -1 0 1070 0 1 5050
box -6 -8 246 248
use DFFPOSX1  _9827_
timestamp 0
transform -1 0 2310 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _9828_
timestamp 0
transform -1 0 2550 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _9829_
timestamp 0
transform 1 0 2170 0 1 6010
box -6 -8 246 248
use DFFPOSX1  _9830_
timestamp 0
transform -1 0 2930 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _9831_
timestamp 0
transform 1 0 2810 0 1 6010
box -6 -8 246 248
use DFFPOSX1  _9832_
timestamp 0
transform -1 0 2710 0 1 6490
box -6 -8 246 248
use DFFPOSX1  _9833_
timestamp 0
transform -1 0 1670 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _9834_
timestamp 0
transform -1 0 1110 0 -1 5530
box -6 -8 246 248
use DFFPOSX1  _9835_
timestamp 0
transform 1 0 1210 0 1 6010
box -6 -8 246 248
use DFFPOSX1  _9836_
timestamp 0
transform -1 0 950 0 1 6490
box -6 -8 246 248
use DFFPOSX1  _9837_
timestamp 0
transform -1 0 5410 0 -1 6490
box -6 -8 246 248
use DFFPOSX1  _9838_
timestamp 0
transform -1 0 4330 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _9839_
timestamp 0
transform 1 0 3390 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _9840_
timestamp 0
transform 1 0 4010 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _9841_
timestamp 0
transform 1 0 4710 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _9842_
timestamp 0
transform -1 0 3570 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _9843_
timestamp 0
transform 1 0 3090 0 1 4090
box -6 -8 246 248
use INVX1  _9844_
timestamp 0
transform 1 0 9490 0 1 5050
box -6 -8 66 248
use INVX2  _9845_
timestamp 0
transform 1 0 9850 0 1 4570
box -6 -8 66 248
use NOR2X1  _9846_
timestamp 0
transform 1 0 11270 0 1 4570
box -6 -8 86 248
use INVX2  _9847_
timestamp 0
transform 1 0 9970 0 1 4570
box -6 -8 66 248
use NOR2X1  _9848_
timestamp 0
transform 1 0 11690 0 -1 6970
box -6 -8 86 248
use INVX4  _9849_
timestamp 0
transform 1 0 11870 0 -1 4090
box -6 -8 86 248
use NOR2X1  _9850_
timestamp 0
transform -1 0 10890 0 -1 4090
box -6 -8 86 248
use OAI21X1  _9851_
timestamp 0
transform -1 0 11090 0 1 6490
box -6 -8 106 248
use INVX2  _9852_
timestamp 0
transform 1 0 10550 0 -1 4090
box -6 -8 66 248
use AND2X2  _9853_
timestamp 0
transform 1 0 10650 0 -1 4090
box -6 -8 106 248
use AOI22X1  _9854_
timestamp 0
transform -1 0 10810 0 1 6490
box -6 -8 126 248
use OAI21X1  _9855_
timestamp 0
transform -1 0 10950 0 1 6490
box -6 -8 106 248
use NOR2X1  _9856_
timestamp 0
transform -1 0 9870 0 -1 4570
box -6 -8 86 248
use AOI22X1  _9857_
timestamp 0
transform 1 0 9890 0 -1 6010
box -6 -8 126 248
use OAI21X1  _9858_
timestamp 0
transform -1 0 9150 0 -1 5530
box -6 -8 106 248
use INVX1  _9859_
timestamp 0
transform 1 0 11710 0 1 7450
box -6 -8 66 248
use OAI21X1  _9860_
timestamp 0
transform -1 0 11910 0 -1 6970
box -6 -8 106 248
use AOI21X1  _9861_
timestamp 0
transform -1 0 11650 0 -1 6970
box -6 -8 106 248
use INVX1  _9862_
timestamp 0
transform -1 0 10530 0 -1 7450
box -6 -8 66 248
use NAND2X1  _9863_
timestamp 0
transform 1 0 9870 0 1 6490
box -6 -8 86 248
use OAI21X1  _9864_
timestamp 0
transform -1 0 10510 0 1 6970
box -6 -8 106 248
use OAI21X1  _9865_
timestamp 0
transform -1 0 10330 0 -1 6970
box -6 -8 106 248
use AOI22X1  _9866_
timestamp 0
transform 1 0 9450 0 1 6010
box -6 -8 126 248
use NAND2X1  _9867_
timestamp 0
transform -1 0 9350 0 -1 6970
box -6 -8 86 248
use INVX1  _9868_
timestamp 0
transform -1 0 14210 0 -1 6490
box -6 -8 66 248
use OAI21X1  _9869_
timestamp 0
transform -1 0 12710 0 1 6490
box -6 -8 106 248
use AOI21X1  _9870_
timestamp 0
transform -1 0 12690 0 -1 6490
box -6 -8 106 248
use INVX1  _9871_
timestamp 0
transform -1 0 13710 0 -1 6490
box -6 -8 66 248
use NAND2X1  _9872_
timestamp 0
transform -1 0 12950 0 -1 6490
box -6 -8 86 248
use OAI21X1  _9873_
timestamp 0
transform 1 0 12730 0 -1 6490
box -6 -8 106 248
use OAI21X1  _9874_
timestamp 0
transform -1 0 12550 0 -1 6490
box -6 -8 106 248
use AOI22X1  _9875_
timestamp 0
transform -1 0 12310 0 1 6010
box -6 -8 126 248
use NAND2X1  _9876_
timestamp 0
transform -1 0 12270 0 -1 6490
box -6 -8 86 248
use INVX1  _9877_
timestamp 0
transform -1 0 13270 0 -1 6970
box -6 -8 66 248
use OAI21X1  _9878_
timestamp 0
transform -1 0 13030 0 -1 6970
box -6 -8 106 248
use AOI21X1  _9879_
timestamp 0
transform -1 0 13170 0 -1 6970
box -6 -8 106 248
use INVX1  _9880_
timestamp 0
transform -1 0 13050 0 -1 6490
box -6 -8 66 248
use NAND2X1  _9881_
timestamp 0
transform -1 0 12990 0 1 6490
box -6 -8 86 248
use OAI21X1  _9882_
timestamp 0
transform 1 0 12750 0 1 6490
box -6 -8 106 248
use OAI21X1  _9883_
timestamp 0
transform -1 0 12870 0 -1 6970
box -6 -8 106 248
use AOI22X1  _9884_
timestamp 0
transform 1 0 12350 0 1 6010
box -6 -8 126 248
use NAND2X1  _9885_
timestamp 0
transform 1 0 12630 0 -1 6970
box -6 -8 86 248
use INVX1  _9886_
timestamp 0
transform 1 0 13590 0 1 2650
box -6 -8 66 248
use OAI21X1  _9887_
timestamp 0
transform -1 0 12330 0 -1 3610
box -6 -8 106 248
use AOI21X1  _9888_
timestamp 0
transform -1 0 12290 0 1 3610
box -6 -8 106 248
use INVX1  _9889_
timestamp 0
transform 1 0 12330 0 1 3130
box -6 -8 66 248
use NAND2X1  _9890_
timestamp 0
transform -1 0 11330 0 -1 4090
box -6 -8 86 248
use OAI21X1  _9891_
timestamp 0
transform -1 0 11470 0 -1 4090
box -6 -8 106 248
use OAI21X1  _9892_
timestamp 0
transform -1 0 11190 0 -1 4090
box -6 -8 106 248
use AOI22X1  _9893_
timestamp 0
transform -1 0 11030 0 -1 4570
box -6 -8 126 248
use NAND2X1  _9894_
timestamp 0
transform -1 0 10850 0 -1 4570
box -6 -8 86 248
use INVX1  _9895_
timestamp 0
transform 1 0 11910 0 1 3610
box -6 -8 66 248
use NOR2X1  _9896_
timestamp 0
transform -1 0 11670 0 -1 3610
box -6 -8 86 248
use OAI21X1  _9897_
timestamp 0
transform -1 0 11830 0 -1 3610
box -6 -8 106 248
use AOI22X1  _9898_
timestamp 0
transform 1 0 11290 0 -1 3610
box -6 -8 126 248
use OAI21X1  _9899_
timestamp 0
transform -1 0 11550 0 -1 3610
box -6 -8 106 248
use AOI22X1  _9900_
timestamp 0
transform 1 0 10470 0 -1 4570
box -6 -8 126 248
use OAI21X1  _9901_
timestamp 0
transform -1 0 10410 0 -1 4570
box -6 -8 106 248
use INVX1  _9902_
timestamp 0
transform -1 0 12590 0 1 6010
box -6 -8 66 248
use INVX1  _9903_
timestamp 0
transform 1 0 12950 0 1 5530
box -6 -8 66 248
use INVX8  _9904_
timestamp 0
transform 1 0 15030 0 1 4570
box -6 -8 126 248
use INVX8  _9905_
timestamp 0
transform 1 0 15550 0 1 4090
box -6 -8 126 248
use INVX1  _9906_
timestamp 0
transform 1 0 15030 0 -1 3130
box -6 -8 66 248
use NAND2X1  _9907_
timestamp 0
transform -1 0 14850 0 -1 3130
box -6 -8 86 248
use OAI21X1  _9908_
timestamp 0
transform -1 0 14990 0 -1 3130
box -6 -8 106 248
use INVX1  _9909_
timestamp 0
transform -1 0 13430 0 -1 3610
box -6 -8 66 248
use NAND2X1  _9910_
timestamp 0
transform -1 0 14230 0 1 3610
box -6 -8 86 248
use OAI21X1  _9911_
timestamp 0
transform 1 0 14010 0 1 3610
box -6 -8 106 248
use MUX2X1  _9912_
timestamp 0
transform -1 0 14110 0 -1 4090
box -6 -8 126 248
use INVX1  _9913_
timestamp 0
transform -1 0 13450 0 1 4570
box -6 -8 66 248
use NAND2X1  _9914_
timestamp 0
transform -1 0 13210 0 1 4570
box -6 -8 86 248
use OAI21X1  _9915_
timestamp 0
transform -1 0 13350 0 1 4570
box -6 -8 106 248
use INVX1  _9916_
timestamp 0
transform -1 0 12650 0 1 4570
box -6 -8 66 248
use NAND2X1  _9917_
timestamp 0
transform 1 0 13810 0 1 4570
box -6 -8 86 248
use OAI21X1  _9918_
timestamp 0
transform 1 0 13670 0 1 4570
box -6 -8 106 248
use MUX2X1  _9919_
timestamp 0
transform 1 0 13510 0 1 4570
box -6 -8 126 248
use MUX2X1  _9920_
timestamp 0
transform -1 0 13610 0 -1 5050
box -6 -8 126 248
use NOR2X1  _9921_
timestamp 0
transform 1 0 12590 0 1 5530
box -6 -8 86 248
use NAND2X1  _9922_
timestamp 0
transform 1 0 13050 0 1 5530
box -6 -8 86 248
use INVX1  _9923_
timestamp 0
transform -1 0 12910 0 1 5530
box -6 -8 66 248
use NAND2X1  _9924_
timestamp 0
transform 1 0 12670 0 -1 5530
box -6 -8 86 248
use OAI21X1  _9925_
timestamp 0
transform -1 0 12430 0 1 3610
box -6 -8 106 248
use INVX2  _9926_
timestamp 0
transform -1 0 12450 0 -1 3610
box -6 -8 66 248
use OAI21X1  _9927_
timestamp 0
transform 1 0 12710 0 1 5530
box -6 -8 106 248
use OAI21X1  _9928_
timestamp 0
transform 1 0 12730 0 -1 6010
box -6 -8 106 248
use INVX8  _9929_
timestamp 0
transform -1 0 11050 0 -1 4090
box -6 -8 126 248
use NAND2X1  _9930_
timestamp 0
transform -1 0 12290 0 -1 6010
box -6 -8 86 248
use NOR2X1  _9931_
timestamp 0
transform -1 0 14010 0 1 5050
box -6 -8 86 248
use MUX2X1  _9932_
timestamp 0
transform 1 0 14330 0 1 4090
box -6 -8 126 248
use MUX2X1  _9933_
timestamp 0
transform 1 0 13730 0 1 4090
box -6 -8 126 248
use MUX2X1  _9934_
timestamp 0
transform -1 0 14530 0 1 4570
box -6 -8 126 248
use INVX2  _9935_
timestamp 0
transform -1 0 11670 0 -1 5530
box -6 -8 66 248
use NAND2X1  _9936_
timestamp 0
transform -1 0 12870 0 -1 5050
box -6 -8 86 248
use AOI21X1  _9937_
timestamp 0
transform 1 0 13070 0 -1 5050
box -6 -8 106 248
use NAND3X1  _9938_
timestamp 0
transform 1 0 12650 0 -1 5050
box -6 -8 106 248
use NAND3X1  _9939_
timestamp 0
transform -1 0 14030 0 1 4570
box -6 -8 106 248
use NAND3X1  _9940_
timestamp 0
transform -1 0 13030 0 -1 5050
box -6 -8 106 248
use OAI22X1  _9941_
timestamp 0
transform 1 0 13210 0 -1 5050
box -6 -8 126 248
use INVX1  _9942_
timestamp 0
transform 1 0 13810 0 1 5050
box -6 -8 66 248
use INVX8  _9943_
timestamp 0
transform 1 0 14870 0 1 4570
box -6 -8 126 248
use INVX1  _9944_
timestamp 0
transform 1 0 15810 0 -1 2170
box -6 -8 66 248
use NAND2X1  _9945_
timestamp 0
transform -1 0 16030 0 1 2170
box -6 -8 86 248
use OAI21X1  _9946_
timestamp 0
transform 1 0 15790 0 1 2170
box -6 -8 106 248
use INVX1  _9947_
timestamp 0
transform -1 0 13830 0 -1 3610
box -6 -8 66 248
use NAND2X1  _9948_
timestamp 0
transform 1 0 14470 0 -1 4090
box -6 -8 86 248
use OAI21X1  _9949_
timestamp 0
transform 1 0 14330 0 -1 4090
box -6 -8 106 248
use MUX2X1  _9950_
timestamp 0
transform -1 0 14290 0 -1 4090
box -6 -8 126 248
use INVX1  _9951_
timestamp 0
transform -1 0 13650 0 -1 4090
box -6 -8 66 248
use NAND2X1  _9952_
timestamp 0
transform 1 0 13850 0 -1 4090
box -6 -8 86 248
use OAI21X1  _9953_
timestamp 0
transform 1 0 13690 0 -1 4090
box -6 -8 106 248
use INVX1  _9954_
timestamp 0
transform -1 0 13750 0 -1 4570
box -6 -8 66 248
use NAND2X1  _9955_
timestamp 0
transform -1 0 13190 0 1 4090
box -6 -8 86 248
use OAI21X1  _9956_
timestamp 0
transform -1 0 13330 0 1 4090
box -6 -8 106 248
use MUX2X1  _9957_
timestamp 0
transform -1 0 13670 0 1 4090
box -6 -8 126 248
use MUX2X1  _9958_
timestamp 0
transform -1 0 13490 0 1 4090
box -6 -8 126 248
use NAND3X1  _9959_
timestamp 0
transform 1 0 13250 0 -1 5530
box -6 -8 106 248
use MUX2X1  _9960_
timestamp 0
transform 1 0 14490 0 1 4090
box -6 -8 126 248
use MUX2X1  _9961_
timestamp 0
transform 1 0 13890 0 1 4090
box -6 -8 126 248
use MUX2X1  _9962_
timestamp 0
transform -1 0 14790 0 1 4090
box -6 -8 126 248
use MUX2X1  _9963_
timestamp 0
transform 1 0 14330 0 -1 4570
box -6 -8 126 248
use MUX2X1  _9964_
timestamp 0
transform 1 0 14170 0 -1 4570
box -6 -8 126 248
use MUX2X1  _9965_
timestamp 0
transform 1 0 14490 0 -1 4570
box -6 -8 126 248
use MUX2X1  _9966_
timestamp 0
transform 1 0 14670 0 -1 4570
box -6 -8 126 248
use OAI21X1  _9967_
timestamp 0
transform 1 0 13830 0 -1 5530
box -6 -8 106 248
use AOI21X1  _9968_
timestamp 0
transform 1 0 13690 0 -1 5530
box -6 -8 106 248
use INVX1  _9969_
timestamp 0
transform -1 0 13690 0 1 5530
box -6 -8 66 248
use NAND3X1  _9970_
timestamp 0
transform 1 0 13550 0 -1 5530
box -6 -8 106 248
use AND2X2  _9971_
timestamp 0
transform -1 0 13570 0 1 5530
box -6 -8 106 248
use OAI21X1  _9972_
timestamp 0
transform 1 0 13170 0 1 5530
box -6 -8 106 248
use OR2X2  _9973_
timestamp 0
transform -1 0 13410 0 1 5530
box -6 -8 106 248
use AOI21X1  _9974_
timestamp 0
transform 1 0 13330 0 -1 6010
box -6 -8 106 248
use OAI21X1  _9975_
timestamp 0
transform 1 0 12330 0 -1 6010
box -6 -8 106 248
use INVX1  _9976_
timestamp 0
transform 1 0 7750 0 1 11290
box -6 -8 66 248
use NAND2X1  _9977_
timestamp 0
transform -1 0 8290 0 1 7930
box -6 -8 86 248
use OAI21X1  _9978_
timestamp 0
transform 1 0 7710 0 -1 11290
box -6 -8 106 248
use NAND2X1  _9979_
timestamp 0
transform 1 0 12870 0 1 6010
box -6 -8 86 248
use AOI21X1  _9980_
timestamp 0
transform 1 0 13730 0 1 5530
box -6 -8 106 248
use MUX2X1  _9981_
timestamp 0
transform -1 0 15490 0 1 4090
box -6 -8 126 248
use MUX2X1  _9982_
timestamp 0
transform 1 0 15190 0 1 4570
box -6 -8 126 248
use MUX2X1  _9983_
timestamp 0
transform 1 0 14250 0 1 4570
box -6 -8 126 248
use NAND2X1  _9984_
timestamp 0
transform -1 0 13990 0 -1 5050
box -6 -8 86 248
use OAI22X1  _9985_
timestamp 0
transform 1 0 14070 0 1 4570
box -6 -8 126 248
use AOI21X1  _9986_
timestamp 0
transform -1 0 14690 0 1 4570
box -6 -8 106 248
use AOI21X1  _9987_
timestamp 0
transform -1 0 14290 0 -1 5530
box -6 -8 106 248
use NAND2X1  _9988_
timestamp 0
transform 1 0 14190 0 1 5530
box -6 -8 86 248
use INVX1  _9989_
timestamp 0
transform -1 0 14150 0 -1 5530
box -6 -8 66 248
use OAI21X1  _9990_
timestamp 0
transform 1 0 13410 0 -1 5530
box -6 -8 106 248
use NAND2X1  _9991_
timestamp 0
transform -1 0 14050 0 -1 5530
box -6 -8 86 248
use AOI21X1  _9992_
timestamp 0
transform -1 0 13970 0 1 5530
box -6 -8 106 248
use NAND3X1  _9993_
timestamp 0
transform 1 0 14030 0 1 5530
box -6 -8 106 248
use INVX1  _9994_
timestamp 0
transform 1 0 14610 0 -1 6010
box -6 -8 66 248
use OR2X2  _9995_
timestamp 0
transform -1 0 14270 0 -1 6010
box -6 -8 106 248
use NOR2X1  _9996_
timestamp 0
transform 1 0 14030 0 -1 6010
box -6 -8 86 248
use INVX1  _9997_
timestamp 0
transform -1 0 13990 0 -1 6010
box -6 -8 66 248
use OAI21X1  _9998_
timestamp 0
transform -1 0 14410 0 -1 6010
box -6 -8 106 248
use AOI21X1  _9999_
timestamp 0
transform -1 0 13870 0 -1 6010
box -6 -8 106 248
use INVX2  _10000_
timestamp 0
transform 1 0 13310 0 1 5050
box -6 -8 66 248
use OAI21X1  _10001_
timestamp 0
transform -1 0 13730 0 -1 6010
box -6 -8 106 248
use OAI21X1  _10002_
timestamp 0
transform -1 0 13570 0 -1 6010
box -6 -8 106 248
use INVX1  _10003_
timestamp 0
transform -1 0 13310 0 1 6010
box -6 -8 66 248
use INVX2  _10004_
timestamp 0
transform 1 0 13750 0 1 6010
box -6 -8 66 248
use OAI21X1  _10005_
timestamp 0
transform 1 0 14470 0 -1 6010
box -6 -8 106 248
use INVX1  _10006_
timestamp 0
transform -1 0 14210 0 1 6010
box -6 -8 66 248
use INVX1  _10007_
timestamp 0
transform -1 0 14670 0 1 5050
box -6 -8 66 248
use NAND3X1  _10008_
timestamp 0
transform 1 0 14350 0 -1 5530
box -6 -8 106 248
use INVX1  _10009_
timestamp 0
transform 1 0 16210 0 -1 2650
box -6 -8 66 248
use NAND2X1  _10010_
timestamp 0
transform 1 0 16470 0 -1 2650
box -6 -8 86 248
use OAI21X1  _10011_
timestamp 0
transform 1 0 16310 0 -1 2650
box -6 -8 106 248
use NAND2X1  _10012_
timestamp 0
transform -1 0 15310 0 1 4090
box -6 -8 86 248
use OAI21X1  _10013_
timestamp 0
transform -1 0 15830 0 1 4090
box -6 -8 106 248
use NOR2X1  _10014_
timestamp 0
transform -1 0 14810 0 -1 4090
box -6 -8 86 248
use NOR2X1  _10015_
timestamp 0
transform 1 0 14490 0 1 5050
box -6 -8 86 248
use AOI22X1  _10016_
timestamp 0
transform 1 0 14170 0 1 4090
box -6 -8 126 248
use OAI21X1  _10017_
timestamp 0
transform -1 0 15630 0 -1 4570
box -6 -8 106 248
use NAND3X1  _10018_
timestamp 0
transform 1 0 14830 0 1 5530
box -6 -8 106 248
use INVX1  _10019_
timestamp 0
transform -1 0 14370 0 1 5530
box -6 -8 66 248
use INVX1  _10020_
timestamp 0
transform -1 0 14790 0 1 5530
box -6 -8 66 248
use OAI21X1  _10021_
timestamp 0
transform 1 0 14410 0 1 5530
box -6 -8 106 248
use NAND3X1  _10022_
timestamp 0
transform -1 0 14830 0 -1 6010
box -6 -8 106 248
use AOI21X1  _10023_
timestamp 0
transform 1 0 14870 0 -1 6010
box -6 -8 106 248
use INVX1  _10024_
timestamp 0
transform -1 0 14450 0 1 6010
box -6 -8 66 248
use NAND2X1  _10025_
timestamp 0
transform -1 0 14350 0 1 6010
box -6 -8 86 248
use AOI21X1  _10026_
timestamp 0
transform -1 0 14110 0 1 6010
box -6 -8 106 248
use OAI21X1  _10027_
timestamp 0
transform -1 0 13970 0 1 6010
box -6 -8 106 248
use AOI22X1  _10028_
timestamp 0
transform 1 0 13590 0 1 6010
box -6 -8 126 248
use AOI21X1  _10029_
timestamp 0
transform 1 0 14510 0 1 6010
box -6 -8 106 248
use INVX1  _10030_
timestamp 0
transform 1 0 14970 0 -1 5050
box -6 -8 66 248
use INVX1  _10031_
timestamp 0
transform 1 0 16810 0 1 2650
box -6 -8 66 248
use NAND2X1  _10032_
timestamp 0
transform -1 0 15270 0 -1 17050
box -6 -8 86 248
use OAI21X1  _10033_
timestamp 0
transform 1 0 16890 0 1 3130
box -6 -8 106 248
use NAND2X1  _10034_
timestamp 0
transform -1 0 16130 0 -1 4570
box -6 -8 86 248
use OAI21X1  _10035_
timestamp 0
transform -1 0 16270 0 -1 4570
box -6 -8 106 248
use NAND2X1  _10036_
timestamp 0
transform -1 0 14790 0 -1 5050
box -6 -8 86 248
use OAI21X1  _10037_
timestamp 0
transform -1 0 14930 0 -1 5050
box -6 -8 106 248
use INVX2  _10038_
timestamp 0
transform 1 0 15230 0 -1 5530
box -6 -8 66 248
use OAI21X1  _10039_
timestamp 0
transform -1 0 15050 0 -1 5530
box -6 -8 106 248
use OR2X2  _10040_
timestamp 0
transform 1 0 15090 0 -1 5530
box -6 -8 106 248
use NOR2X1  _10041_
timestamp 0
transform 1 0 15130 0 1 5530
box -6 -8 86 248
use OAI21X1  _10042_
timestamp 0
transform 1 0 14970 0 1 5530
box -6 -8 106 248
use NAND3X1  _10043_
timestamp 0
transform -1 0 15110 0 -1 6010
box -6 -8 106 248
use NOR2X1  _10044_
timestamp 0
transform -1 0 14730 0 -1 5530
box -6 -8 86 248
use AND2X2  _10045_
timestamp 0
transform -1 0 14590 0 -1 5530
box -6 -8 106 248
use OAI21X1  _10046_
timestamp 0
transform 1 0 14790 0 -1 5530
box -6 -8 106 248
use NAND2X1  _10047_
timestamp 0
transform -1 0 14730 0 1 6010
box -6 -8 86 248
use AOI21X1  _10048_
timestamp 0
transform -1 0 14930 0 -1 6490
box -6 -8 106 248
use OAI21X1  _10049_
timestamp 0
transform -1 0 14770 0 -1 6490
box -6 -8 106 248
use AOI22X1  _10050_
timestamp 0
transform 1 0 13990 0 -1 6490
box -6 -8 126 248
use OAI21X1  _10051_
timestamp 0
transform 1 0 14990 0 -1 6490
box -6 -8 106 248
use INVX1  _10052_
timestamp 0
transform 1 0 15570 0 -1 5050
box -6 -8 66 248
use NAND3X1  _10053_
timestamp 0
transform 1 0 14570 0 1 5530
box -6 -8 106 248
use NAND2X1  _10054_
timestamp 0
transform 1 0 16390 0 -1 4090
box -6 -8 86 248
use INVX1  _10055_
timestamp 0
transform -1 0 16370 0 1 4090
box -6 -8 66 248
use AOI21X1  _10056_
timestamp 0
transform 1 0 16030 0 1 4090
box -6 -8 106 248
use NAND2X1  _10057_
timestamp 0
transform -1 0 15870 0 -1 4570
box -6 -8 86 248
use OAI21X1  _10058_
timestamp 0
transform -1 0 15910 0 1 4570
box -6 -8 106 248
use NAND3X1  _10059_
timestamp 0
transform -1 0 15490 0 1 5530
box -6 -8 106 248
use NOR3X1  _10060_
timestamp 0
transform 1 0 15350 0 -1 5530
box -6 -8 186 248
use INVX1  _10061_
timestamp 0
transform 1 0 15710 0 -1 5530
box -6 -8 66 248
use OAI21X1  _10062_
timestamp 0
transform -1 0 15670 0 -1 5530
box -6 -8 106 248
use NAND3X1  _10063_
timestamp 0
transform -1 0 15550 0 -1 6010
box -6 -8 106 248
use AOI21X1  _10064_
timestamp 0
transform -1 0 15390 0 -1 6010
box -6 -8 106 248
use INVX1  _10065_
timestamp 0
transform 1 0 15350 0 1 6010
box -6 -8 66 248
use NAND2X1  _10066_
timestamp 0
transform 1 0 15270 0 -1 6490
box -6 -8 86 248
use AND2X2  _10067_
timestamp 0
transform -1 0 14990 0 -1 6970
box -6 -8 106 248
use OAI21X1  _10068_
timestamp 0
transform 1 0 14990 0 1 6490
box -6 -8 106 248
use OAI21X1  _10069_
timestamp 0
transform -1 0 14950 0 1 6490
box -6 -8 106 248
use OAI21X1  _10070_
timestamp 0
transform 1 0 13050 0 1 6490
box -6 -8 106 248
use INVX1  _10071_
timestamp 0
transform 1 0 14450 0 1 6490
box -6 -8 66 248
use INVX1  _10072_
timestamp 0
transform -1 0 15670 0 -1 6010
box -6 -8 66 248
use NAND3X1  _10073_
timestamp 0
transform 1 0 15250 0 1 5530
box -6 -8 106 248
use AOI21X1  _10074_
timestamp 0
transform -1 0 16270 0 1 4090
box -6 -8 106 248
use NAND2X1  _10075_
timestamp 0
transform -1 0 16050 0 1 4570
box -6 -8 86 248
use OAI21X1  _10076_
timestamp 0
transform -1 0 16190 0 1 4570
box -6 -8 106 248
use NAND3X1  _10077_
timestamp 0
transform 1 0 15710 0 1 5530
box -6 -8 106 248
use INVX1  _10078_
timestamp 0
transform 1 0 15970 0 1 5530
box -6 -8 66 248
use OAI21X1  _10079_
timestamp 0
transform 1 0 15550 0 1 5530
box -6 -8 106 248
use NAND2X1  _10080_
timestamp 0
transform 1 0 15850 0 1 5530
box -6 -8 86 248
use NAND3X1  _10081_
timestamp 0
transform -1 0 15810 0 -1 6010
box -6 -8 106 248
use NAND3X1  _10082_
timestamp 0
transform 1 0 16090 0 1 5530
box -6 -8 106 248
use NAND2X1  _10083_
timestamp 0
transform -1 0 16090 0 -1 6010
box -6 -8 86 248
use NAND3X1  _10084_
timestamp 0
transform 1 0 16150 0 -1 6010
box -6 -8 106 248
use NAND2X1  _10085_
timestamp 0
transform -1 0 15710 0 -1 6490
box -6 -8 86 248
use AOI21X1  _10086_
timestamp 0
transform 1 0 15150 0 -1 6010
box -6 -8 106 248
use NOR2X1  _10087_
timestamp 0
transform -1 0 15150 0 1 6010
box -6 -8 86 248
use OAI21X1  _10088_
timestamp 0
transform 1 0 14910 0 1 6010
box -6 -8 106 248
use NAND2X1  _10089_
timestamp 0
transform -1 0 15230 0 -1 6490
box -6 -8 86 248
use AOI21X1  _10090_
timestamp 0
transform -1 0 15390 0 1 6490
box -6 -8 106 248
use OAI21X1  _10091_
timestamp 0
transform -1 0 15250 0 1 6490
box -6 -8 106 248
use AOI22X1  _10092_
timestamp 0
transform 1 0 14550 0 1 6490
box -6 -8 126 248
use INVX1  _10093_
timestamp 0
transform -1 0 13250 0 1 6490
box -6 -8 66 248
use AOI21X1  _10094_
timestamp 0
transform 1 0 15870 0 -1 6010
box -6 -8 106 248
use AND2X2  _10095_
timestamp 0
transform 1 0 14770 0 1 6010
box -6 -8 106 248
use NAND3X1  _10096_
timestamp 0
transform 1 0 15470 0 1 6010
box -6 -8 106 248
use AOI21X1  _10097_
timestamp 0
transform 1 0 15190 0 1 6010
box -6 -8 106 248
use OAI21X1  _10098_
timestamp 0
transform 1 0 15630 0 1 6010
box -6 -8 106 248
use AOI21X1  _10099_
timestamp 0
transform -1 0 15870 0 1 6010
box -6 -8 106 248
use INVX1  _10100_
timestamp 0
transform 1 0 15910 0 1 5050
box -6 -8 66 248
use NAND3X1  _10101_
timestamp 0
transform 1 0 15830 0 -1 5530
box -6 -8 106 248
use INVX1  _10102_
timestamp 0
transform 1 0 16510 0 -1 4090
box -6 -8 66 248
use NOR2X1  _10103_
timestamp 0
transform 1 0 16530 0 1 4570
box -6 -8 86 248
use INVX1  _10104_
timestamp 0
transform 1 0 16650 0 1 4570
box -6 -8 66 248
use OAI21X1  _10105_
timestamp 0
transform 1 0 16230 0 1 4570
box -6 -8 106 248
use NAND3X1  _10106_
timestamp 0
transform -1 0 16410 0 1 5050
box -6 -8 106 248
use INVX1  _10107_
timestamp 0
transform -1 0 16150 0 -1 5050
box -6 -8 66 248
use OAI21X1  _10108_
timestamp 0
transform 1 0 16250 0 1 5530
box -6 -8 106 248
use NAND2X1  _10109_
timestamp 0
transform 1 0 16170 0 1 5050
box -6 -8 86 248
use NAND3X1  _10110_
timestamp 0
transform -1 0 16130 0 1 5050
box -6 -8 106 248
use NAND3X1  _10111_
timestamp 0
transform -1 0 16230 0 -1 5530
box -6 -8 106 248
use NAND2X1  _10112_
timestamp 0
transform 1 0 16270 0 -1 5530
box -6 -8 86 248
use NAND3X1  _10113_
timestamp 0
transform 1 0 15990 0 -1 5530
box -6 -8 106 248
use NAND2X1  _10114_
timestamp 0
transform 1 0 15890 0 -1 6490
box -6 -8 86 248
use INVX1  _10115_
timestamp 0
transform -1 0 15590 0 -1 6490
box -6 -8 66 248
use NOR2X1  _10116_
timestamp 0
transform 1 0 15390 0 -1 6490
box -6 -8 86 248
use OAI21X1  _10117_
timestamp 0
transform 1 0 15590 0 1 6490
box -6 -8 106 248
use OAI21X1  _10118_
timestamp 0
transform -1 0 15530 0 1 6490
box -6 -8 106 248
use OAI21X1  _10119_
timestamp 0
transform 1 0 13490 0 -1 6490
box -6 -8 106 248
use INVX1  _10120_
timestamp 0
transform 1 0 13710 0 1 6490
box -6 -8 66 248
use OAI21X1  _10121_
timestamp 0
transform -1 0 14810 0 1 6490
box -6 -8 106 248
use OAI21X1  _10122_
timestamp 0
transform 1 0 13550 0 1 6490
box -6 -8 106 248
use INVX1  _10123_
timestamp 0
transform 1 0 13910 0 -1 6970
box -6 -8 66 248
use OAI21X1  _10124_
timestamp 0
transform 1 0 16010 0 1 6490
box -6 -8 106 248
use NOR2X1  _10125_
timestamp 0
transform 1 0 15750 0 1 6490
box -6 -8 86 248
use AOI21X1  _10126_
timestamp 0
transform 1 0 15870 0 1 6490
box -6 -8 106 248
use INVX1  _10127_
timestamp 0
transform 1 0 16530 0 1 5530
box -6 -8 66 248
use OR2X2  _10128_
timestamp 0
transform 1 0 16390 0 -1 5530
box -6 -8 106 248
use OAI21X1  _10129_
timestamp 0
transform 1 0 16490 0 -1 5050
box -6 -8 106 248
use NAND3X1  _10130_
timestamp 0
transform -1 0 16890 0 1 5530
box -6 -8 106 248
use NOR2X1  _10131_
timestamp 0
transform -1 0 16610 0 -1 5530
box -6 -8 86 248
use INVX1  _10132_
timestamp 0
transform -1 0 17010 0 -1 5530
box -6 -8 66 248
use OAI21X1  _10133_
timestamp 0
transform 1 0 16790 0 -1 5530
box -6 -8 106 248
use NAND3X1  _10134_
timestamp 0
transform 1 0 16650 0 1 5530
box -6 -8 106 248
use NAND3X1  _10135_
timestamp 0
transform 1 0 16930 0 1 5530
box -6 -8 106 248
use OAI21X1  _10136_
timestamp 0
transform -1 0 16750 0 -1 5530
box -6 -8 106 248
use NAND3X1  _10137_
timestamp 0
transform -1 0 16970 0 -1 6010
box -6 -8 106 248
use AND2X2  _10138_
timestamp 0
transform 1 0 16630 0 1 6010
box -6 -8 106 248
use INVX1  _10139_
timestamp 0
transform -1 0 16530 0 1 6490
box -6 -8 66 248
use AOI21X1  _10140_
timestamp 0
transform -1 0 16250 0 1 6490
box -6 -8 106 248
use OAI21X1  _10141_
timestamp 0
transform -1 0 16410 0 1 6490
box -6 -8 106 248
use AOI22X1  _10142_
timestamp 0
transform 1 0 14050 0 1 6490
box -6 -8 126 248
use NAND2X1  _10143_
timestamp 0
transform -1 0 15990 0 1 6010
box -6 -8 86 248
use AND2X2  _10144_
timestamp 0
transform -1 0 16150 0 1 6010
box -6 -8 106 248
use AND2X2  _10145_
timestamp 0
transform 1 0 15750 0 -1 6490
box -6 -8 106 248
use NAND3X1  _10146_
timestamp 0
transform 1 0 16030 0 -1 6490
box -6 -8 106 248
use OAI21X1  _10147_
timestamp 0
transform 1 0 16170 0 -1 6490
box -6 -8 106 248
use INVX1  _10148_
timestamp 0
transform 1 0 16610 0 -1 6010
box -6 -8 66 248
use AOI21X1  _10149_
timestamp 0
transform -1 0 16550 0 -1 6010
box -6 -8 106 248
use INVX1  _10150_
timestamp 0
transform -1 0 16530 0 -1 6970
box -6 -8 66 248
use NOR3X1  _10151_
timestamp 0
transform 1 0 16470 0 1 5050
box -6 -8 186 248
use INVX1  _10152_
timestamp 0
transform 1 0 17050 0 -1 5050
box -6 -8 66 248
use OAI21X1  _10153_
timestamp 0
transform 1 0 16650 0 -1 5050
box -6 -8 106 248
use NAND3X1  _10154_
timestamp 0
transform 1 0 16990 0 1 5050
box -6 -8 106 248
use INVX1  _10155_
timestamp 0
transform 1 0 16950 0 -1 5050
box -6 -8 66 248
use OAI21X1  _10156_
timestamp 0
transform 1 0 16810 0 -1 5050
box -6 -8 106 248
use NAND3X1  _10157_
timestamp 0
transform 1 0 17070 0 1 5530
box -6 -8 106 248
use NAND3X1  _10158_
timestamp 0
transform 1 0 16270 0 -1 17050
box -6 -8 106 248
use OAI21X1  _10159_
timestamp 0
transform 1 0 16690 0 1 5050
box -6 -8 106 248
use NAND3X1  _10160_
timestamp 0
transform 1 0 16850 0 1 5050
box -6 -8 106 248
use AND2X2  _10161_
timestamp 0
transform -1 0 16810 0 -1 6010
box -6 -8 106 248
use AND2X2  _10162_
timestamp 0
transform -1 0 16430 0 1 6010
box -6 -8 106 248
use OAI21X1  _10163_
timestamp 0
transform -1 0 16410 0 -1 6010
box -6 -8 106 248
use OAI21X1  _10164_
timestamp 0
transform -1 0 16290 0 1 6010
box -6 -8 106 248
use OAI21X1  _10165_
timestamp 0
transform 1 0 13350 0 -1 6490
box -6 -8 106 248
use INVX1  _10166_
timestamp 0
transform 1 0 16830 0 1 4090
box -6 -8 66 248
use OAI21X1  _10167_
timestamp 0
transform 1 0 16370 0 1 4570
box -6 -8 106 248
use INVX1  _10168_
timestamp 0
transform -1 0 17130 0 1 4570
box -6 -8 66 248
use AOI21X1  _10169_
timestamp 0
transform 1 0 15730 0 -1 17050
box -6 -8 106 248
use NAND3X1  _10170_
timestamp 0
transform -1 0 17010 0 1 4570
box -6 -8 106 248
use NAND2X1  _10171_
timestamp 0
transform -1 0 17010 0 1 4090
box -6 -8 86 248
use NAND2X1  _10172_
timestamp 0
transform 1 0 16770 0 1 4570
box -6 -8 86 248
use OAI21X1  _10173_
timestamp 0
transform -1 0 16210 0 -1 17050
box -6 -8 106 248
use NAND2X1  _10174_
timestamp 0
transform 1 0 17030 0 1 250
box -6 -8 86 248
use INVX1  _10175_
timestamp 0
transform -1 0 17170 0 1 2170
box -6 -8 66 248
use AND2X2  _10176_
timestamp 0
transform -1 0 17150 0 1 4090
box -6 -8 106 248
use NAND2X1  _10177_
timestamp 0
transform 1 0 16990 0 -1 4570
box -6 -8 86 248
use NAND3X1  _10178_
timestamp 0
transform -1 0 16930 0 -1 4570
box -6 -8 106 248
use NAND2X1  _10179_
timestamp 0
transform 1 0 17070 0 1 6010
box -6 -8 86 248
use AOI21X1  _10180_
timestamp 0
transform -1 0 17150 0 -1 5530
box -6 -8 106 248
use AOI21X1  _10181_
timestamp 0
transform 1 0 17010 0 -1 6010
box -6 -8 106 248
use NAND3X1  _10182_
timestamp 0
transform 1 0 16490 0 1 6010
box -6 -8 106 248
use AOI21X1  _10183_
timestamp 0
transform -1 0 17010 0 1 6010
box -6 -8 106 248
use AND2X2  _10184_
timestamp 0
transform -1 0 17130 0 -1 6490
box -6 -8 106 248
use NAND3X1  _10185_
timestamp 0
transform -1 0 16870 0 1 6010
box -6 -8 106 248
use OAI21X1  _10186_
timestamp 0
transform 1 0 16610 0 -1 6490
box -6 -8 106 248
use OAI21X1  _10187_
timestamp 0
transform -1 0 16570 0 -1 6490
box -6 -8 106 248
use OR2X2  _10188_
timestamp 0
transform -1 0 16410 0 -1 6490
box -6 -8 106 248
use AOI22X1  _10189_
timestamp 0
transform 1 0 14510 0 -1 6490
box -6 -8 126 248
use NAND2X1  _10190_
timestamp 0
transform -1 0 12190 0 1 6490
box -6 -8 86 248
use INVX1  _10191_
timestamp 0
transform -1 0 16970 0 -1 6490
box -6 -8 66 248
use NAND2X1  _10192_
timestamp 0
transform 1 0 17070 0 1 3610
box -6 -8 86 248
use INVX1  _10193_
timestamp 0
transform 1 0 16830 0 -1 3610
box -6 -8 66 248
use NAND2X1  _10194_
timestamp 0
transform -1 0 17030 0 -1 3610
box -6 -8 86 248
use NAND2X1  _10195_
timestamp 0
transform 1 0 17070 0 -1 3610
box -6 -8 86 248
use INVX1  _10196_
timestamp 0
transform 1 0 16770 0 -1 4090
box -6 -8 66 248
use NAND2X1  _10197_
timestamp 0
transform 1 0 15310 0 -1 17050
box -6 -8 86 248
use NAND2X1  _10198_
timestamp 0
transform -1 0 16950 0 -1 4090
box -6 -8 86 248
use NAND2X1  _10199_
timestamp 0
transform 1 0 17010 0 -1 4090
box -6 -8 86 248
use INVX1  _10200_
timestamp 0
transform 1 0 17110 0 1 6490
box -6 -8 66 248
use NOR3X1  _10201_
timestamp 0
transform -1 0 17070 0 1 6490
box -6 -8 186 248
use AOI21X1  _10202_
timestamp 0
transform 1 0 16750 0 -1 6490
box -6 -8 106 248
use OAI21X1  _10203_
timestamp 0
transform -1 0 16830 0 1 6490
box -6 -8 106 248
use OAI21X1  _10204_
timestamp 0
transform -1 0 16670 0 1 6490
box -6 -8 106 248
use NAND2X1  _10205_
timestamp 0
transform 1 0 12470 0 1 6490
box -6 -8 86 248
use NAND2X1  _10206_
timestamp 0
transform -1 0 11670 0 -1 4570
box -6 -8 86 248
use INVX1  _10207_
timestamp 0
transform 1 0 14310 0 -1 5050
box -6 -8 66 248
use NAND2X1  _10208_
timestamp 0
transform 1 0 14570 0 -1 5050
box -6 -8 86 248
use OAI21X1  _10209_
timestamp 0
transform 1 0 14410 0 -1 5050
box -6 -8 106 248
use NAND2X1  _10210_
timestamp 0
transform 1 0 14190 0 -1 5050
box -6 -8 86 248
use NOR2X1  _10211_
timestamp 0
transform -1 0 12870 0 -1 5530
box -6 -8 86 248
use NOR2X1  _10212_
timestamp 0
transform -1 0 12610 0 -1 5530
box -6 -8 86 248
use AOI22X1  _10213_
timestamp 0
transform -1 0 13190 0 -1 5530
box -6 -8 126 248
use NAND3X1  _10214_
timestamp 0
transform -1 0 14130 0 -1 5050
box -6 -8 106 248
use NAND2X1  _10215_
timestamp 0
transform 1 0 15790 0 1 5050
box -6 -8 86 248
use OAI21X1  _10216_
timestamp 0
transform 1 0 15670 0 -1 5050
box -6 -8 106 248
use NAND2X1  _10217_
timestamp 0
transform 1 0 15510 0 1 4570
box -6 -8 86 248
use OAI21X1  _10218_
timestamp 0
transform 1 0 15370 0 1 4570
box -6 -8 106 248
use MUX2X1  _10219_
timestamp 0
transform 1 0 15390 0 -1 4090
box -6 -8 126 248
use NAND2X1  _10220_
timestamp 0
transform 1 0 15410 0 1 3610
box -6 -8 86 248
use AND2X2  _10221_
timestamp 0
transform 1 0 14950 0 1 3610
box -6 -8 106 248
use NOR2X1  _10222_
timestamp 0
transform 1 0 13010 0 -1 4570
box -6 -8 86 248
use NAND2X1  _10223_
timestamp 0
transform -1 0 15330 0 -1 4570
box -6 -8 86 248
use NAND2X1  _10224_
timestamp 0
transform 1 0 15670 0 -1 4570
box -6 -8 86 248
use NAND2X1  _10225_
timestamp 0
transform 1 0 15390 0 -1 4570
box -6 -8 86 248
use OAI21X1  _10226_
timestamp 0
transform -1 0 15210 0 -1 4570
box -6 -8 106 248
use OAI21X1  _10227_
timestamp 0
transform 1 0 13270 0 -1 4570
box -6 -8 106 248
use OAI21X1  _10228_
timestamp 0
transform -1 0 12050 0 -1 4570
box -6 -8 106 248
use NAND2X1  _10229_
timestamp 0
transform 1 0 10850 0 1 4570
box -6 -8 86 248
use NOR2X1  _10230_
timestamp 0
transform 1 0 13130 0 -1 4570
box -6 -8 86 248
use NAND2X1  _10231_
timestamp 0
transform -1 0 14950 0 1 5050
box -6 -8 86 248
use OAI21X1  _10232_
timestamp 0
transform 1 0 14730 0 1 5050
box -6 -8 106 248
use NAND2X1  _10233_
timestamp 0
transform -1 0 14270 0 1 5050
box -6 -8 86 248
use OAI21X1  _10234_
timestamp 0
transform -1 0 14430 0 1 5050
box -6 -8 106 248
use MUX2X1  _10235_
timestamp 0
transform 1 0 14950 0 -1 4570
box -6 -8 126 248
use NAND2X1  _10236_
timestamp 0
transform -1 0 15610 0 1 3610
box -6 -8 86 248
use NAND2X1  _10237_
timestamp 0
transform -1 0 15910 0 -1 5050
box -6 -8 86 248
use OAI21X1  _10238_
timestamp 0
transform -1 0 16050 0 -1 5050
box -6 -8 106 248
use INVX1  _10239_
timestamp 0
transform 1 0 15970 0 1 3610
box -6 -8 66 248
use NAND2X1  _10240_
timestamp 0
transform -1 0 15730 0 1 5050
box -6 -8 86 248
use OAI21X1  _10241_
timestamp 0
transform 1 0 15650 0 1 4570
box -6 -8 106 248
use NAND2X1  _10242_
timestamp 0
transform -1 0 15810 0 -1 4090
box -6 -8 86 248
use OAI21X1  _10243_
timestamp 0
transform -1 0 15910 0 1 3610
box -6 -8 106 248
use OAI21X1  _10244_
timestamp 0
transform -1 0 15770 0 1 3610
box -6 -8 106 248
use NAND3X1  _10245_
timestamp 0
transform -1 0 14370 0 1 3610
box -6 -8 106 248
use MUX2X1  _10246_
timestamp 0
transform -1 0 15690 0 -1 4090
box -6 -8 126 248
use MUX2X1  _10247_
timestamp 0
transform 1 0 15110 0 -1 4090
box -6 -8 126 248
use OAI21X1  _10248_
timestamp 0
transform 1 0 14590 0 -1 4090
box -6 -8 106 248
use AOI21X1  _10249_
timestamp 0
transform -1 0 12890 0 1 4090
box -6 -8 106 248
use INVX1  _10250_
timestamp 0
transform -1 0 12430 0 1 4090
box -6 -8 66 248
use NAND3X1  _10251_
timestamp 0
transform -1 0 13050 0 1 4090
box -6 -8 106 248
use AND2X2  _10252_
timestamp 0
transform 1 0 12470 0 1 4090
box -6 -8 106 248
use NAND2X1  _10253_
timestamp 0
transform 1 0 12710 0 1 4570
box -6 -8 86 248
use OR2X2  _10254_
timestamp 0
transform 1 0 12830 0 1 4570
box -6 -8 106 248
use AOI21X1  _10255_
timestamp 0
transform 1 0 12970 0 1 4570
box -6 -8 106 248
use OAI21X1  _10256_
timestamp 0
transform -1 0 11090 0 1 4570
box -6 -8 106 248
use NAND2X1  _10257_
timestamp 0
transform -1 0 11150 0 -1 4570
box -6 -8 86 248
use AOI21X1  _10258_
timestamp 0
transform 1 0 12630 0 1 4090
box -6 -8 106 248
use NAND2X1  _10259_
timestamp 0
transform 1 0 14550 0 1 3610
box -6 -8 86 248
use NAND2X1  _10260_
timestamp 0
transform 1 0 16350 0 -1 5050
box -6 -8 86 248
use OAI21X1  _10261_
timestamp 0
transform 1 0 16190 0 -1 5050
box -6 -8 106 248
use NAND2X1  _10262_
timestamp 0
transform -1 0 16190 0 -1 4090
box -6 -8 86 248
use OAI21X1  _10263_
timestamp 0
transform 1 0 16250 0 -1 4090
box -6 -8 106 248
use NAND2X1  _10264_
timestamp 0
transform -1 0 14810 0 1 4570
box -6 -8 86 248
use NAND2X1  _10265_
timestamp 0
transform -1 0 15050 0 1 4090
box -6 -8 86 248
use NAND2X1  _10266_
timestamp 0
transform 1 0 14830 0 1 4090
box -6 -8 86 248
use AOI21X1  _10267_
timestamp 0
transform -1 0 15350 0 1 3610
box -6 -8 106 248
use INVX1  _10268_
timestamp 0
transform -1 0 14610 0 -1 3610
box -6 -8 66 248
use NAND3X1  _10269_
timestamp 0
transform 1 0 14410 0 1 3610
box -6 -8 106 248
use AOI21X1  _10270_
timestamp 0
transform 1 0 15110 0 1 3610
box -6 -8 106 248
use OAI21X1  _10271_
timestamp 0
transform -1 0 14770 0 1 3610
box -6 -8 106 248
use NAND3X1  _10272_
timestamp 0
transform -1 0 13550 0 -1 4090
box -6 -8 106 248
use INVX1  _10273_
timestamp 0
transform 1 0 13190 0 -1 4090
box -6 -8 66 248
use AOI21X1  _10274_
timestamp 0
transform -1 0 13390 0 -1 4090
box -6 -8 106 248
use NOR2X1  _10275_
timestamp 0
transform 1 0 13070 0 -1 4090
box -6 -8 86 248
use AND2X2  _10276_
timestamp 0
transform -1 0 12330 0 -1 4090
box -6 -8 106 248
use NOR2X1  _10277_
timestamp 0
transform 1 0 12250 0 1 4090
box -6 -8 86 248
use OAI21X1  _10278_
timestamp 0
transform -1 0 12190 0 1 4090
box -6 -8 106 248
use OAI21X1  _10279_
timestamp 0
transform -1 0 11530 0 -1 4570
box -6 -8 106 248
use OAI21X1  _10280_
timestamp 0
transform 1 0 12910 0 -1 4090
box -6 -8 106 248
use INVX1  _10281_
timestamp 0
transform -1 0 12930 0 1 3610
box -6 -8 66 248
use NAND2X1  _10282_
timestamp 0
transform 1 0 16710 0 1 4090
box -6 -8 86 248
use OAI21X1  _10283_
timestamp 0
transform 1 0 16550 0 1 4090
box -6 -8 106 248
use MUX2X1  _10284_
timestamp 0
transform 1 0 16090 0 1 3610
box -6 -8 126 248
use NOR2X1  _10285_
timestamp 0
transform 1 0 15750 0 -1 3610
box -6 -8 86 248
use NAND2X1  _10286_
timestamp 0
transform 1 0 14830 0 -1 4570
box -6 -8 86 248
use NAND2X1  _10287_
timestamp 0
transform -1 0 15070 0 -1 4090
box -6 -8 86 248
use NAND2X1  _10288_
timestamp 0
transform 1 0 14850 0 -1 4090
box -6 -8 86 248
use OR2X2  _10289_
timestamp 0
transform 1 0 14810 0 -1 3610
box -6 -8 106 248
use OAI21X1  _10290_
timestamp 0
transform -1 0 14490 0 -1 3610
box -6 -8 106 248
use OR2X2  _10291_
timestamp 0
transform -1 0 14230 0 -1 3610
box -6 -8 106 248
use OAI21X1  _10292_
timestamp 0
transform -1 0 14750 0 -1 3610
box -6 -8 106 248
use AOI21X1  _10293_
timestamp 0
transform -1 0 13570 0 -1 3610
box -6 -8 106 248
use INVX1  _10294_
timestamp 0
transform -1 0 12870 0 -1 3610
box -6 -8 66 248
use NAND3X1  _10295_
timestamp 0
transform 1 0 13610 0 -1 3610
box -6 -8 106 248
use NAND2X1  _10296_
timestamp 0
transform -1 0 12750 0 -1 3610
box -6 -8 86 248
use OR2X2  _10297_
timestamp 0
transform -1 0 12710 0 1 3610
box -6 -8 106 248
use NAND2X1  _10298_
timestamp 0
transform -1 0 12830 0 1 3610
box -6 -8 86 248
use NAND2X1  _10299_
timestamp 0
transform -1 0 12570 0 1 3610
box -6 -8 86 248
use AOI22X1  _10300_
timestamp 0
transform 1 0 12010 0 1 3610
box -6 -8 126 248
use AOI21X1  _10301_
timestamp 0
transform 1 0 12930 0 -1 3610
box -6 -8 106 248
use NAND2X1  _10302_
timestamp 0
transform -1 0 17030 0 1 3610
box -6 -8 86 248
use OAI21X1  _10303_
timestamp 0
transform 1 0 16810 0 1 3610
box -6 -8 106 248
use NAND2X1  _10304_
timestamp 0
transform 1 0 16390 0 1 3610
box -6 -8 86 248
use OAI21X1  _10305_
timestamp 0
transform 1 0 16250 0 1 3610
box -6 -8 106 248
use NAND2X1  _10306_
timestamp 0
transform 1 0 15510 0 -1 3610
box -6 -8 86 248
use OAI21X1  _10307_
timestamp 0
transform 1 0 15350 0 -1 3610
box -6 -8 106 248
use INVX1  _10308_
timestamp 0
transform -1 0 15430 0 1 3130
box -6 -8 66 248
use NAND3X1  _10309_
timestamp 0
transform 1 0 14810 0 1 3610
box -6 -8 106 248
use OAI21X1  _10310_
timestamp 0
transform -1 0 14930 0 1 3130
box -6 -8 106 248
use OR2X2  _10311_
timestamp 0
transform -1 0 14630 0 1 3130
box -6 -8 106 248
use NOR2X1  _10312_
timestamp 0
transform 1 0 14970 0 1 3130
box -6 -8 86 248
use OAI21X1  _10313_
timestamp 0
transform 1 0 15430 0 -1 3130
box -6 -8 106 248
use NAND3X1  _10314_
timestamp 0
transform -1 0 14470 0 1 3130
box -6 -8 106 248
use OR2X2  _10315_
timestamp 0
transform -1 0 14790 0 1 3130
box -6 -8 106 248
use OAI21X1  _10316_
timestamp 0
transform 1 0 15090 0 1 3130
box -6 -8 106 248
use NAND3X1  _10317_
timestamp 0
transform -1 0 13910 0 1 3130
box -6 -8 106 248
use NAND2X1  _10318_
timestamp 0
transform -1 0 13610 0 1 3130
box -6 -8 86 248
use OR2X2  _10319_
timestamp 0
transform -1 0 13330 0 1 3130
box -6 -8 106 248
use NAND2X1  _10320_
timestamp 0
transform -1 0 13470 0 1 3130
box -6 -8 86 248
use NAND2X1  _10321_
timestamp 0
transform -1 0 13190 0 1 3130
box -6 -8 86 248
use AOI22X1  _10322_
timestamp 0
transform 1 0 12450 0 1 3130
box -6 -8 126 248
use INVX1  _10323_
timestamp 0
transform 1 0 12230 0 -1 3130
box -6 -8 66 248
use OAI21X1  _10324_
timestamp 0
transform 1 0 13790 0 -1 3130
box -6 -8 106 248
use NAND2X1  _10325_
timestamp 0
transform 1 0 15850 0 -1 3130
box -6 -8 86 248
use NOR2X1  _10326_
timestamp 0
transform -1 0 16110 0 -1 3610
box -6 -8 86 248
use AOI21X1  _10327_
timestamp 0
transform 1 0 16170 0 -1 3610
box -6 -8 106 248
use NAND2X1  _10328_
timestamp 0
transform 1 0 15850 0 1 3130
box -6 -8 86 248
use OAI21X1  _10329_
timestamp 0
transform -1 0 16070 0 1 3130
box -6 -8 106 248
use INVX1  _10330_
timestamp 0
transform -1 0 16190 0 -1 3130
box -6 -8 66 248
use NAND3X1  _10331_
timestamp 0
transform -1 0 16070 0 -1 3130
box -6 -8 106 248
use NOR2X1  _10332_
timestamp 0
transform 1 0 14970 0 -1 3610
box -6 -8 86 248
use NAND3X1  _10333_
timestamp 0
transform 1 0 15090 0 -1 3610
box -6 -8 106 248
use OAI21X1  _10334_
timestamp 0
transform 1 0 15710 0 1 3130
box -6 -8 106 248
use NAND2X1  _10335_
timestamp 0
transform 1 0 15570 0 -1 3130
box -6 -8 86 248
use AOI21X1  _10336_
timestamp 0
transform -1 0 15230 0 -1 3130
box -6 -8 106 248
use INVX1  _10337_
timestamp 0
transform -1 0 14710 0 -1 3130
box -6 -8 66 248
use NAND3X1  _10338_
timestamp 0
transform 1 0 15270 0 -1 3130
box -6 -8 106 248
use NAND2X1  _10339_
timestamp 0
transform -1 0 14030 0 -1 3130
box -6 -8 86 248
use NOR2X1  _10340_
timestamp 0
transform 1 0 13670 0 -1 3130
box -6 -8 86 248
use AND2X2  _10341_
timestamp 0
transform -1 0 13630 0 -1 3130
box -6 -8 106 248
use OAI21X1  _10342_
timestamp 0
transform -1 0 13470 0 -1 3130
box -6 -8 106 248
use OAI21X1  _10343_
timestamp 0
transform 1 0 12330 0 -1 3130
box -6 -8 106 248
use INVX1  _10344_
timestamp 0
transform 1 0 11390 0 1 3610
box -6 -8 66 248
use NAND3X1  _10345_
timestamp 0
transform -1 0 15790 0 -1 3130
box -6 -8 106 248
use AOI21X1  _10346_
timestamp 0
transform 1 0 16330 0 -1 3610
box -6 -8 106 248
use NAND2X1  _10347_
timestamp 0
transform 1 0 16510 0 -1 3130
box -6 -8 86 248
use OAI21X1  _10348_
timestamp 0
transform 1 0 16370 0 -1 3130
box -6 -8 106 248
use NAND3X1  _10349_
timestamp 0
transform 1 0 15190 0 1 2650
box -6 -8 106 248
use NOR3X1  _10350_
timestamp 0
transform -1 0 15650 0 1 3130
box -6 -8 186 248
use INVX1  _10351_
timestamp 0
transform 1 0 15630 0 1 2650
box -6 -8 66 248
use OAI21X1  _10352_
timestamp 0
transform 1 0 15330 0 1 2650
box -6 -8 106 248
use NAND2X1  _10353_
timestamp 0
transform 1 0 15050 0 1 2650
box -6 -8 86 248
use NAND2X1  _10354_
timestamp 0
transform 1 0 14770 0 1 2650
box -6 -8 86 248
use NAND3X1  _10355_
timestamp 0
transform -1 0 14990 0 1 2650
box -6 -8 106 248
use NAND2X1  _10356_
timestamp 0
transform -1 0 14590 0 1 2650
box -6 -8 86 248
use AOI21X1  _10357_
timestamp 0
transform 1 0 13950 0 1 3130
box -6 -8 106 248
use NOR2X1  _10358_
timestamp 0
transform 1 0 14250 0 1 3130
box -6 -8 86 248
use OAI21X1  _10359_
timestamp 0
transform 1 0 14090 0 1 3130
box -6 -8 106 248
use NAND2X1  _10360_
timestamp 0
transform -1 0 14290 0 -1 3130
box -6 -8 86 248
use NOR2X1  _10361_
timestamp 0
transform -1 0 14330 0 1 2650
box -6 -8 86 248
use AND2X2  _10362_
timestamp 0
transform -1 0 14730 0 1 2650
box -6 -8 106 248
use AND2X2  _10363_
timestamp 0
transform -1 0 13770 0 1 3130
box -6 -8 106 248
use NAND3X1  _10364_
timestamp 0
transform 1 0 14070 0 -1 3130
box -6 -8 106 248
use AOI21X1  _10365_
timestamp 0
transform 1 0 14490 0 -1 3130
box -6 -8 106 248
use OAI21X1  _10366_
timestamp 0
transform 1 0 14330 0 -1 3130
box -6 -8 106 248
use NOR2X1  _10367_
timestamp 0
transform -1 0 14450 0 1 2650
box -6 -8 86 248
use OAI21X1  _10368_
timestamp 0
transform -1 0 13970 0 1 2650
box -6 -8 106 248
use NAND2X1  _10369_
timestamp 0
transform 1 0 12930 0 1 2650
box -6 -8 86 248
use OAI21X1  _10370_
timestamp 0
transform 1 0 11510 0 1 3610
box -6 -8 106 248
use INVX1  _10371_
timestamp 0
transform 1 0 12830 0 -1 3130
box -6 -8 66 248
use INVX1  _10372_
timestamp 0
transform -1 0 14090 0 1 2650
box -6 -8 66 248
use NAND2X1  _10373_
timestamp 0
transform 1 0 15250 0 -1 2650
box -6 -8 86 248
use NOR2X1  _10374_
timestamp 0
transform 1 0 16350 0 1 3130
box -6 -8 86 248
use INVX1  _10375_
timestamp 0
transform 1 0 16490 0 1 3130
box -6 -8 66 248
use OAI21X1  _10376_
timestamp 0
transform 1 0 16230 0 -1 3130
box -6 -8 106 248
use NAND3X1  _10377_
timestamp 0
transform -1 0 14970 0 -1 2650
box -6 -8 106 248
use INVX1  _10378_
timestamp 0
transform -1 0 15210 0 -1 2650
box -6 -8 66 248
use OAI21X1  _10379_
timestamp 0
transform 1 0 15470 0 1 2650
box -6 -8 106 248
use NAND2X1  _10380_
timestamp 0
transform -1 0 15110 0 -1 2650
box -6 -8 86 248
use NAND3X1  _10381_
timestamp 0
transform -1 0 14810 0 -1 2650
box -6 -8 106 248
use NAND3X1  _10382_
timestamp 0
transform 1 0 15530 0 -1 2650
box -6 -8 106 248
use NAND2X1  _10383_
timestamp 0
transform 1 0 15510 0 1 2170
box -6 -8 86 248
use NAND3X1  _10384_
timestamp 0
transform -1 0 15750 0 1 2170
box -6 -8 106 248
use NAND2X1  _10385_
timestamp 0
transform 1 0 15230 0 1 2170
box -6 -8 86 248
use OAI21X1  _10386_
timestamp 0
transform 1 0 13450 0 1 2650
box -6 -8 106 248
use NOR2X1  _10387_
timestamp 0
transform -1 0 13410 0 1 2650
box -6 -8 86 248
use INVX1  _10388_
timestamp 0
transform -1 0 13270 0 1 2650
box -6 -8 66 248
use AOI21X1  _10389_
timestamp 0
transform -1 0 13170 0 1 2650
box -6 -8 106 248
use AOI22X1  _10390_
timestamp 0
transform 1 0 12930 0 -1 3130
box -6 -8 126 248
use OAI21X1  _10391_
timestamp 0
transform 1 0 14570 0 -1 2650
box -6 -8 106 248
use NOR2X1  _10392_
timestamp 0
transform -1 0 14390 0 -1 2650
box -6 -8 86 248
use AOI21X1  _10393_
timestamp 0
transform 1 0 14430 0 -1 2650
box -6 -8 106 248
use INVX1  _10394_
timestamp 0
transform 1 0 16170 0 -1 2170
box -6 -8 66 248
use NAND3X1  _10395_
timestamp 0
transform -1 0 15470 0 -1 2650
box -6 -8 106 248
use INVX1  _10396_
timestamp 0
transform -1 0 16310 0 1 3130
box -6 -8 66 248
use OAI21X1  _10397_
timestamp 0
transform 1 0 16290 0 1 2650
box -6 -8 106 248
use INVX1  _10398_
timestamp 0
transform 1 0 16610 0 1 2170
box -6 -8 66 248
use NAND3X1  _10399_
timestamp 0
transform -1 0 16670 0 -1 2170
box -6 -8 106 248
use OAI21X1  _10400_
timestamp 0
transform 1 0 15670 0 -1 2650
box -6 -8 106 248
use NAND2X1  _10401_
timestamp 0
transform -1 0 16370 0 -1 2170
box -6 -8 86 248
use AOI21X1  _10402_
timestamp 0
transform 1 0 16410 0 -1 2170
box -6 -8 106 248
use NAND3X1  _10403_
timestamp 0
transform -1 0 16830 0 -1 2170
box -6 -8 106 248
use NAND2X1  _10404_
timestamp 0
transform 1 0 16210 0 1 2170
box -6 -8 86 248
use AOI21X1  _10405_
timestamp 0
transform -1 0 16170 0 1 2170
box -6 -8 106 248
use OAI21X1  _10406_
timestamp 0
transform -1 0 14250 0 -1 2650
box -6 -8 106 248
use INVX1  _10407_
timestamp 0
transform -1 0 14190 0 1 2650
box -6 -8 66 248
use OR2X2  _10408_
timestamp 0
transform -1 0 15470 0 1 2170
box -6 -8 106 248
use OAI21X1  _10409_
timestamp 0
transform -1 0 13830 0 -1 2650
box -6 -8 106 248
use OAI22X1  _10410_
timestamp 0
transform 1 0 13690 0 1 2650
box -6 -8 126 248
use NAND2X1  _10411_
timestamp 0
transform 1 0 12810 0 1 2650
box -6 -8 86 248
use NOR2X1  _10412_
timestamp 0
transform -1 0 13950 0 -1 2650
box -6 -8 86 248
use NOR2X1  _10413_
timestamp 0
transform -1 0 14090 0 -1 2650
box -6 -8 86 248
use OAI21X1  _10414_
timestamp 0
transform 1 0 16990 0 -1 3130
box -6 -8 106 248
use INVX1  _10415_
timestamp 0
transform 1 0 16950 0 -1 250
box -6 -8 66 248
use OAI21X1  _10416_
timestamp 0
transform -1 0 16970 0 -1 2170
box -6 -8 106 248
use NAND2X1  _10417_
timestamp 0
transform 1 0 17010 0 -1 2170
box -6 -8 86 248
use OR2X2  _10418_
timestamp 0
transform 1 0 15450 0 -1 17050
box -6 -8 106 248
use NAND3X1  _10419_
timestamp 0
transform 1 0 16950 0 1 2170
box -6 -8 106 248
use NAND2X1  _10420_
timestamp 0
transform 1 0 16970 0 -1 12250
box -6 -8 86 248
use NAND2X1  _10421_
timestamp 0
transform 1 0 16710 0 1 2170
box -6 -8 86 248
use NAND2X1  _10422_
timestamp 0
transform -1 0 16170 0 -1 2650
box -6 -8 86 248
use AND2X2  _10423_
timestamp 0
transform -1 0 13450 0 -1 2650
box -6 -8 106 248
use OAI21X1  _10424_
timestamp 0
transform -1 0 13290 0 -1 2650
box -6 -8 106 248
use OAI21X1  _10425_
timestamp 0
transform -1 0 13150 0 -1 2650
box -6 -8 106 248
use INVX1  _10426_
timestamp 0
transform 1 0 13090 0 -1 3130
box -6 -8 66 248
use INVX1  _10427_
timestamp 0
transform 1 0 16850 0 1 2170
box -6 -8 66 248
use AOI21X1  _10428_
timestamp 0
transform -1 0 16050 0 -1 2650
box -6 -8 106 248
use NOR2X1  _10429_
timestamp 0
transform -1 0 16410 0 1 2170
box -6 -8 86 248
use NAND3X1  _10430_
timestamp 0
transform -1 0 16570 0 1 2170
box -6 -8 106 248
use OAI21X1  _10431_
timestamp 0
transform 1 0 15810 0 -1 2650
box -6 -8 106 248
use OAI21X1  _10432_
timestamp 0
transform -1 0 16450 0 -1 250
box -6 -8 106 248
use INVX1  _10433_
timestamp 0
transform 1 0 16410 0 -1 17050
box -6 -8 66 248
use OR2X2  _10434_
timestamp 0
transform 1 0 16610 0 -1 2650
box -6 -8 106 248
use OAI21X1  _10435_
timestamp 0
transform -1 0 17010 0 -1 2650
box -6 -8 106 248
use NAND2X1  _10436_
timestamp 0
transform 1 0 16870 0 -1 3130
box -6 -8 86 248
use OR2X2  _10437_
timestamp 0
transform -1 0 16870 0 -1 2650
box -6 -8 106 248
use NAND3X1  _10438_
timestamp 0
transform -1 0 16770 0 1 2650
box -6 -8 106 248
use AND2X2  _10439_
timestamp 0
transform 1 0 17070 0 1 2650
box -6 -8 106 248
use NOR2X1  _10440_
timestamp 0
transform -1 0 17130 0 -1 2650
box -6 -8 86 248
use OAI21X1  _10441_
timestamp 0
transform -1 0 17010 0 1 2650
box -6 -8 106 248
use NAND2X1  _10442_
timestamp 0
transform 1 0 16550 0 1 2650
box -6 -8 86 248
use AND2X2  _10443_
timestamp 0
transform 1 0 15990 0 1 2650
box -6 -8 106 248
use NOR2X1  _10444_
timestamp 0
transform -1 0 15950 0 1 2650
box -6 -8 86 248
use NOR2X1  _10445_
timestamp 0
transform -1 0 15810 0 1 2650
box -6 -8 86 248
use AOI22X1  _10446_
timestamp 0
transform 1 0 13210 0 -1 3130
box -6 -8 126 248
use NAND2X1  _10447_
timestamp 0
transform 1 0 12110 0 -1 3610
box -6 -8 86 248
use INVX1  _10448_
timestamp 0
transform 1 0 16430 0 1 2650
box -6 -8 66 248
use AOI21X1  _10449_
timestamp 0
transform 1 0 16150 0 1 2650
box -6 -8 106 248
use NAND2X1  _10450_
timestamp 0
transform 1 0 16710 0 -1 3610
box -6 -8 86 248
use NOR2X1  _10451_
timestamp 0
transform 1 0 16670 0 1 3610
box -6 -8 86 248
use AOI21X1  _10452_
timestamp 0
transform 1 0 16610 0 -1 4090
box -6 -8 106 248
use NOR2X1  _10453_
timestamp 0
transform 1 0 16530 0 1 3610
box -6 -8 86 248
use AND2X2  _10454_
timestamp 0
transform -1 0 13310 0 -1 3610
box -6 -8 106 248
use OAI21X1  _10455_
timestamp 0
transform -1 0 13170 0 -1 3610
box -6 -8 106 248
use OAI21X1  _10456_
timestamp 0
transform -1 0 12610 0 -1 3610
box -6 -8 106 248
use OAI21X1  _10457_
timestamp 0
transform 1 0 11190 0 1 5530
box -6 -8 106 248
use OAI21X1  _10458_
timestamp 0
transform -1 0 9530 0 1 5530
box -6 -8 106 248
use INVX1  _10459_
timestamp 0
transform -1 0 9370 0 1 5530
box -6 -8 66 248
use NOR2X1  _10460_
timestamp 0
transform 1 0 9710 0 1 5530
box -6 -8 86 248
use NAND2X1  _10461_
timestamp 0
transform 1 0 9590 0 1 5530
box -6 -8 86 248
use NAND2X1  _10462_
timestamp 0
transform 1 0 9750 0 -1 6010
box -6 -8 86 248
use NAND2X1  _10463_
timestamp 0
transform 1 0 10010 0 1 6010
box -6 -8 86 248
use OAI21X1  _10464_
timestamp 0
transform 1 0 9850 0 1 6010
box -6 -8 106 248
use NAND2X1  _10465_
timestamp 0
transform 1 0 9310 0 1 6010
box -6 -8 86 248
use INVX1  _10466_
timestamp 0
transform -1 0 9190 0 -1 6010
box -6 -8 66 248
use NOR2X1  _10467_
timestamp 0
transform 1 0 10610 0 1 5530
box -6 -8 86 248
use AOI21X1  _10468_
timestamp 0
transform -1 0 10090 0 -1 5530
box -6 -8 106 248
use NOR2X1  _10469_
timestamp 0
transform -1 0 9930 0 -1 5530
box -6 -8 86 248
use OAI21X1  _10470_
timestamp 0
transform 1 0 9990 0 1 5530
box -6 -8 106 248
use AND2X2  _10471_
timestamp 0
transform -1 0 9930 0 1 5530
box -6 -8 106 248
use OR2X2  _10472_
timestamp 0
transform -1 0 9010 0 -1 5530
box -6 -8 106 248
use OR2X2  _10473_
timestamp 0
transform -1 0 8770 0 1 5530
box -6 -8 106 248
use OAI21X1  _10474_
timestamp 0
transform -1 0 8870 0 -1 5530
box -6 -8 106 248
use NAND2X1  _10475_
timestamp 0
transform -1 0 8730 0 -1 5530
box -6 -8 86 248
use NOR2X1  _10476_
timestamp 0
transform -1 0 8870 0 1 6010
box -6 -8 86 248
use NAND2X1  _10477_
timestamp 0
transform -1 0 8970 0 -1 6010
box -6 -8 86 248
use NAND2X1  _10478_
timestamp 0
transform -1 0 9090 0 -1 6010
box -6 -8 86 248
use OAI21X1  _10479_
timestamp 0
transform 1 0 8910 0 1 6010
box -6 -8 106 248
use INVX1  _10480_
timestamp 0
transform 1 0 8830 0 1 5530
box -6 -8 66 248
use OAI21X1  _10481_
timestamp 0
transform 1 0 8930 0 1 5530
box -6 -8 106 248
use OAI21X1  _10482_
timestamp 0
transform -1 0 11230 0 -1 5050
box -6 -8 106 248
use OAI21X1  _10483_
timestamp 0
transform -1 0 10350 0 -1 5050
box -6 -8 106 248
use MUX2X1  _10484_
timestamp 0
transform -1 0 10530 0 -1 5050
box -6 -8 126 248
use NAND2X1  _10485_
timestamp 0
transform 1 0 9370 0 -1 5050
box -6 -8 86 248
use OR2X2  _10486_
timestamp 0
transform -1 0 9330 0 -1 5050
box -6 -8 106 248
use NAND2X1  _10487_
timestamp 0
transform 1 0 9110 0 -1 5050
box -6 -8 86 248
use INVX1  _10488_
timestamp 0
transform -1 0 9050 0 -1 5050
box -6 -8 66 248
use NOR2X1  _10489_
timestamp 0
transform -1 0 8830 0 -1 5050
box -6 -8 86 248
use NAND2X1  _10490_
timestamp 0
transform -1 0 8950 0 -1 5050
box -6 -8 86 248
use NAND2X1  _10491_
timestamp 0
transform 1 0 9770 0 1 5050
box -6 -8 86 248
use OAI22X1  _10492_
timestamp 0
transform 1 0 9610 0 1 5050
box -6 -8 126 248
use NOR2X1  _10493_
timestamp 0
transform -1 0 9590 0 -1 6010
box -6 -8 86 248
use NAND2X1  _10494_
timestamp 0
transform 1 0 9910 0 1 5050
box -6 -8 86 248
use INVX1  _10495_
timestamp 0
transform 1 0 10030 0 1 5050
box -6 -8 66 248
use INVX1  _10496_
timestamp 0
transform 1 0 10290 0 1 5050
box -6 -8 66 248
use NOR2X1  _10497_
timestamp 0
transform 1 0 11330 0 -1 5530
box -6 -8 86 248
use OAI21X1  _10498_
timestamp 0
transform -1 0 11290 0 -1 5530
box -6 -8 106 248
use OAI21X1  _10499_
timestamp 0
transform 1 0 11050 0 1 5530
box -6 -8 106 248
use OAI21X1  _10500_
timestamp 0
transform -1 0 11150 0 -1 5530
box -6 -8 106 248
use NOR2X1  _10501_
timestamp 0
transform 1 0 10530 0 1 5050
box -6 -8 86 248
use NAND2X1  _10502_
timestamp 0
transform 1 0 10390 0 1 5050
box -6 -8 86 248
use INVX1  _10503_
timestamp 0
transform -1 0 9690 0 -1 5530
box -6 -8 66 248
use NOR2X1  _10504_
timestamp 0
transform -1 0 9590 0 -1 5530
box -6 -8 86 248
use OAI21X1  _10505_
timestamp 0
transform -1 0 9290 0 -1 5530
box -6 -8 106 248
use AOI21X1  _10506_
timestamp 0
transform 1 0 9350 0 -1 5530
box -6 -8 106 248
use NOR2X1  _10507_
timestamp 0
transform 1 0 9630 0 -1 6010
box -6 -8 86 248
use NAND2X1  _10508_
timestamp 0
transform 1 0 11030 0 -1 6970
box -6 -8 86 248
use INVX1  _10509_
timestamp 0
transform -1 0 10650 0 1 6010
box -6 -8 66 248
use AOI21X1  _10510_
timestamp 0
transform -1 0 10990 0 1 5530
box -6 -8 106 248
use OAI21X1  _10511_
timestamp 0
transform 1 0 10750 0 1 5530
box -6 -8 106 248
use OAI21X1  _10512_
timestamp 0
transform 1 0 10130 0 1 5530
box -6 -8 106 248
use OR2X2  _10513_
timestamp 0
transform 1 0 10530 0 -1 6490
box -6 -8 106 248
use NAND2X1  _10514_
timestamp 0
transform -1 0 10470 0 -1 6490
box -6 -8 86 248
use NAND2X1  _10515_
timestamp 0
transform 1 0 10490 0 -1 6970
box -6 -8 86 248
use AOI21X1  _10516_
timestamp 0
transform 1 0 10130 0 1 5050
box -6 -8 106 248
use AND2X2  _10517_
timestamp 0
transform 1 0 10730 0 -1 6970
box -6 -8 106 248
use OAI21X1  _10518_
timestamp 0
transform 1 0 11010 0 1 6970
box -6 -8 106 248
use OAI21X1  _10519_
timestamp 0
transform -1 0 10970 0 -1 6970
box -6 -8 106 248
use OAI21X1  _10520_
timestamp 0
transform -1 0 10950 0 1 6970
box -6 -8 106 248
use INVX1  _10521_
timestamp 0
transform -1 0 11250 0 1 6010
box -6 -8 66 248
use OAI21X1  _10522_
timestamp 0
transform -1 0 13010 0 -1 5530
box -6 -8 106 248
use OAI21X1  _10523_
timestamp 0
transform 1 0 13170 0 -1 6010
box -6 -8 106 248
use OR2X2  _10524_
timestamp 0
transform -1 0 13110 0 -1 6010
box -6 -8 106 248
use NAND2X1  _10525_
timestamp 0
transform -1 0 12970 0 -1 6010
box -6 -8 86 248
use OR2X2  _10526_
timestamp 0
transform -1 0 11050 0 -1 6490
box -6 -8 106 248
use NAND2X1  _10527_
timestamp 0
transform -1 0 11190 0 -1 6490
box -6 -8 86 248
use NAND2X1  _10528_
timestamp 0
transform -1 0 10910 0 -1 6490
box -6 -8 86 248
use INVX1  _10529_
timestamp 0
transform -1 0 10630 0 1 6490
box -6 -8 66 248
use NOR2X1  _10530_
timestamp 0
transform 1 0 11010 0 -1 7450
box -6 -8 86 248
use NAND2X1  _10531_
timestamp 0
transform 1 0 10870 0 -1 7450
box -6 -8 86 248
use NAND2X1  _10532_
timestamp 0
transform 1 0 10750 0 -1 7450
box -6 -8 86 248
use OAI22X1  _10533_
timestamp 0
transform 1 0 10570 0 -1 7450
box -6 -8 126 248
use NAND2X1  _10534_
timestamp 0
transform -1 0 9550 0 1 6490
box -6 -8 86 248
use INVX1  _10535_
timestamp 0
transform 1 0 10630 0 -1 6970
box -6 -8 66 248
use NAND2X1  _10536_
timestamp 0
transform -1 0 10790 0 1 6970
box -6 -8 86 248
use OAI21X1  _10537_
timestamp 0
transform 1 0 10690 0 -1 6490
box -6 -8 106 248
use INVX1  _10538_
timestamp 0
transform 1 0 10370 0 -1 6970
box -6 -8 66 248
use OAI21X1  _10539_
timestamp 0
transform -1 0 10670 0 1 6970
box -6 -8 106 248
use OAI21X1  _10540_
timestamp 0
transform -1 0 11550 0 -1 5530
box -6 -8 106 248
use NOR2X1  _10541_
timestamp 0
transform 1 0 10930 0 -1 5530
box -6 -8 86 248
use NAND2X1  _10542_
timestamp 0
transform -1 0 10610 0 -1 5530
box -6 -8 86 248
use OAI21X1  _10543_
timestamp 0
transform -1 0 10890 0 -1 5530
box -6 -8 106 248
use NAND2X1  _10544_
timestamp 0
transform -1 0 10750 0 -1 5530
box -6 -8 86 248
use NAND2X1  _10545_
timestamp 0
transform 1 0 10870 0 -1 6010
box -6 -8 86 248
use OR2X2  _10546_
timestamp 0
transform 1 0 11010 0 -1 6010
box -6 -8 106 248
use NAND2X1  _10547_
timestamp 0
transform 1 0 10470 0 1 6010
box -6 -8 86 248
use INVX1  _10548_
timestamp 0
transform -1 0 10190 0 -1 6970
box -6 -8 66 248
use NOR2X1  _10549_
timestamp 0
transform -1 0 9970 0 -1 6970
box -6 -8 86 248
use NAND2X1  _10550_
timestamp 0
transform -1 0 10090 0 -1 6970
box -6 -8 86 248
use NAND2X1  _10551_
timestamp 0
transform 1 0 9750 0 1 6490
box -6 -8 86 248
use OAI21X1  _10552_
timestamp 0
transform -1 0 9690 0 1 6490
box -6 -8 106 248
use INVX1  _10553_
timestamp 0
transform -1 0 9330 0 -1 6490
box -6 -8 66 248
use NAND2X1  _10554_
timestamp 0
transform -1 0 9930 0 -1 6490
box -6 -8 86 248
use INVX1  _10555_
timestamp 0
transform 1 0 10270 0 1 5530
box -6 -8 66 248
use NAND2X1  _10556_
timestamp 0
transform 1 0 10750 0 -1 6010
box -6 -8 86 248
use OR2X2  _10557_
timestamp 0
transform -1 0 10690 0 -1 6010
box -6 -8 106 248
use NAND2X1  _10558_
timestamp 0
transform -1 0 10550 0 -1 6010
box -6 -8 86 248
use NOR2X1  _10559_
timestamp 0
transform -1 0 10270 0 -1 6010
box -6 -8 86 248
use INVX1  _10560_
timestamp 0
transform -1 0 10190 0 1 6010
box -6 -8 66 248
use NAND2X1  _10561_
timestamp 0
transform 1 0 10330 0 -1 6010
box -6 -8 86 248
use NAND2X1  _10562_
timestamp 0
transform -1 0 10350 0 -1 6490
box -6 -8 86 248
use OR2X2  _10563_
timestamp 0
transform -1 0 9650 0 -1 6490
box -6 -8 106 248
use AOI21X1  _10564_
timestamp 0
transform -1 0 9790 0 -1 6490
box -6 -8 106 248
use AOI22X1  _10565_
timestamp 0
transform 1 0 9370 0 -1 6490
box -6 -8 126 248
use NAND2X1  _10566_
timestamp 0
transform 1 0 11170 0 1 6970
box -6 -8 86 248
use NOR2X1  _10567_
timestamp 0
transform -1 0 11410 0 1 5530
box -6 -8 86 248
use INVX1  _10568_
timestamp 0
transform 1 0 11470 0 1 5530
box -6 -8 66 248
use NAND3X1  _10569_
timestamp 0
transform -1 0 11530 0 -1 6010
box -6 -8 106 248
use INVX1  _10570_
timestamp 0
transform -1 0 11210 0 1 6490
box -6 -8 66 248
use AOI21X1  _10571_
timestamp 0
transform 1 0 11570 0 -1 6010
box -6 -8 106 248
use NOR2X1  _10572_
timestamp 0
transform -1 0 11310 0 -1 6490
box -6 -8 86 248
use OAI21X1  _10573_
timestamp 0
transform 1 0 10130 0 -1 6490
box -6 -8 106 248
use NOR2X1  _10574_
timestamp 0
transform 1 0 9990 0 1 6490
box -6 -8 86 248
use AOI21X1  _10575_
timestamp 0
transform 1 0 10130 0 1 6490
box -6 -8 106 248
use NAND3X1  _10576_
timestamp 0
transform -1 0 10530 0 1 6490
box -6 -8 106 248
use OAI21X1  _10577_
timestamp 0
transform -1 0 10390 0 1 6490
box -6 -8 106 248
use NOR2X1  _10578_
timestamp 0
transform 1 0 11430 0 1 6970
box -6 -8 86 248
use NAND2X1  _10579_
timestamp 0
transform 1 0 11550 0 1 6970
box -6 -8 86 248
use NAND2X1  _10580_
timestamp 0
transform 1 0 11690 0 1 6970
box -6 -8 86 248
use OAI21X1  _10581_
timestamp 0
transform -1 0 11390 0 1 6970
box -6 -8 106 248
use AOI21X1  _10582_
timestamp 0
transform 1 0 11410 0 -1 6970
box -6 -8 106 248
use OR2X2  _10583_
timestamp 0
transform 1 0 11530 0 1 6010
box -6 -8 106 248
use NAND2X1  _10584_
timestamp 0
transform 1 0 11670 0 1 6010
box -6 -8 86 248
use NAND2X1  _10585_
timestamp 0
transform -1 0 11730 0 -1 6490
box -6 -8 86 248
use AND2X2  _10586_
timestamp 0
transform -1 0 11470 0 -1 7450
box -6 -8 106 248
use OAI21X1  _10587_
timestamp 0
transform 1 0 11690 0 -1 7450
box -6 -8 106 248
use OAI22X1  _10588_
timestamp 0
transform -1 0 11630 0 -1 7450
box -6 -8 126 248
use NAND2X1  _10589_
timestamp 0
transform -1 0 11910 0 1 6970
box -6 -8 86 248
use OAI21X1  _10590_
timestamp 0
transform -1 0 11450 0 -1 6490
box -6 -8 106 248
use NAND3X1  _10591_
timestamp 0
transform -1 0 11590 0 -1 6490
box -6 -8 106 248
use INVX1  _10592_
timestamp 0
transform -1 0 11330 0 1 6490
box -6 -8 66 248
use AOI21X1  _10593_
timestamp 0
transform 1 0 11370 0 1 6490
box -6 -8 106 248
use INVX1  _10594_
timestamp 0
transform -1 0 11950 0 1 6490
box -6 -8 66 248
use NAND2X1  _10595_
timestamp 0
transform -1 0 12130 0 -1 6490
box -6 -8 86 248
use NAND2X1  _10596_
timestamp 0
transform 1 0 11930 0 -1 6490
box -6 -8 86 248
use NAND2X1  _10597_
timestamp 0
transform -1 0 12070 0 1 6490
box -6 -8 86 248
use AND2X2  _10598_
timestamp 0
transform 1 0 12490 0 1 6970
box -6 -8 106 248
use OAI21X1  _10599_
timestamp 0
transform -1 0 12450 0 1 6970
box -6 -8 106 248
use OAI21X1  _10600_
timestamp 0
transform -1 0 12290 0 1 6970
box -6 -8 106 248
use NAND2X1  _10601_
timestamp 0
transform -1 0 12050 0 -1 6970
box -6 -8 86 248
use OAI21X1  _10602_
timestamp 0
transform -1 0 12330 0 -1 6970
box -6 -8 106 248
use OAI21X1  _10603_
timestamp 0
transform -1 0 12190 0 -1 6970
box -6 -8 106 248
use NAND2X1  _10604_
timestamp 0
transform 1 0 10490 0 1 4090
box -6 -8 86 248
use NAND2X1  _10605_
timestamp 0
transform -1 0 11350 0 -1 5050
box -6 -8 86 248
use NOR2X1  _10606_
timestamp 0
transform 1 0 10630 0 1 4090
box -6 -8 86 248
use NAND2X1  _10607_
timestamp 0
transform 1 0 15230 0 1 3130
box -6 -8 86 248
use OAI21X1  _10608_
timestamp 0
transform -1 0 16710 0 1 3130
box -6 -8 106 248
use NAND2X1  _10609_
timestamp 0
transform -1 0 16190 0 1 3130
box -6 -8 86 248
use OAI21X1  _10610_
timestamp 0
transform 1 0 16750 0 1 3130
box -6 -8 106 248
use INVX1  _10611_
timestamp 0
transform 1 0 11610 0 1 4090
box -6 -8 66 248
use OR2X2  _10612_
timestamp 0
transform 1 0 10750 0 1 4090
box -6 -8 106 248
use OAI21X1  _10613_
timestamp 0
transform 1 0 11310 0 1 4090
box -6 -8 106 248
use OAI21X1  _10614_
timestamp 0
transform -1 0 11550 0 1 4090
box -6 -8 106 248
use INVX1  _10615_
timestamp 0
transform -1 0 11250 0 1 4090
box -6 -8 66 248
use OAI21X1  _10616_
timestamp 0
transform 1 0 10910 0 1 4090
box -6 -8 106 248
use OAI21X1  _10617_
timestamp 0
transform -1 0 11150 0 1 4090
box -6 -8 106 248
use NAND2X1  _10618_
timestamp 0
transform -1 0 10730 0 -1 4570
box -6 -8 86 248
use NAND2X1  _10619_
timestamp 0
transform -1 0 12850 0 -1 4090
box -6 -8 86 248
use OAI21X1  _10620_
timestamp 0
transform 1 0 12630 0 -1 4090
box -6 -8 106 248
use NAND2X1  _10621_
timestamp 0
transform 1 0 11990 0 -1 4090
box -6 -8 86 248
use OAI21X1  _10622_
timestamp 0
transform 1 0 11950 0 1 4090
box -6 -8 106 248
use AND2X2  _10623_
timestamp 0
transform 1 0 10170 0 -1 4570
box -6 -8 106 248
use NAND2X1  _10624_
timestamp 0
transform 1 0 13610 0 1 3610
box -6 -8 86 248
use OAI21X1  _10625_
timestamp 0
transform 1 0 13470 0 1 3610
box -6 -8 106 248
use NAND2X1  _10626_
timestamp 0
transform -1 0 13810 0 1 3610
box -6 -8 86 248
use OAI21X1  _10627_
timestamp 0
transform -1 0 13970 0 1 3610
box -6 -8 106 248
use OAI21X1  _10628_
timestamp 0
transform 1 0 12430 0 1 4570
box -6 -8 106 248
use OAI21X1  _10629_
timestamp 0
transform 1 0 12090 0 -1 4570
box -6 -8 106 248
use OAI21X1  _10630_
timestamp 0
transform -1 0 12390 0 1 4570
box -6 -8 106 248
use OAI21X1  _10631_
timestamp 0
transform 1 0 11890 0 1 4570
box -6 -8 106 248
use NAND2X1  _10632_
timestamp 0
transform 1 0 12490 0 -1 4570
box -6 -8 86 248
use OAI21X1  _10633_
timestamp 0
transform -1 0 12710 0 -1 4570
box -6 -8 106 248
use NAND2X1  _10634_
timestamp 0
transform -1 0 13490 0 -1 4570
box -6 -8 86 248
use OAI21X1  _10635_
timestamp 0
transform 1 0 13550 0 -1 4570
box -6 -8 106 248
use NAND2X1  _10636_
timestamp 0
transform 1 0 16310 0 -1 4570
box -6 -8 86 248
use OAI21X1  _10637_
timestamp 0
transform -1 0 16550 0 -1 4570
box -6 -8 106 248
use NAND2X1  _10638_
timestamp 0
transform 1 0 15230 0 -1 3610
box -6 -8 86 248
use OAI21X1  _10639_
timestamp 0
transform -1 0 15990 0 -1 3610
box -6 -8 106 248
use INVX1  _10640_
timestamp 0
transform -1 0 11910 0 1 5050
box -6 -8 66 248
use OAI21X1  _10641_
timestamp 0
transform -1 0 12210 0 1 5050
box -6 -8 106 248
use OAI21X1  _10642_
timestamp 0
transform 1 0 11970 0 1 5050
box -6 -8 106 248
use INVX1  _10643_
timestamp 0
transform -1 0 12050 0 -1 5050
box -6 -8 66 248
use OAI21X1  _10644_
timestamp 0
transform 1 0 12410 0 1 5050
box -6 -8 106 248
use OAI21X1  _10645_
timestamp 0
transform 1 0 12250 0 1 5050
box -6 -8 106 248
use NAND2X1  _10646_
timestamp 0
transform -1 0 12490 0 -1 5530
box -6 -8 86 248
use OAI21X1  _10647_
timestamp 0
transform 1 0 12030 0 -1 5530
box -6 -8 106 248
use NAND2X1  _10648_
timestamp 0
transform -1 0 13030 0 1 5050
box -6 -8 86 248
use OAI21X1  _10649_
timestamp 0
transform 1 0 12810 0 1 5050
box -6 -8 106 248
use NAND2X1  _10650_
timestamp 0
transform 1 0 15390 0 1 5050
box -6 -8 86 248
use OAI21X1  _10651_
timestamp 0
transform 1 0 15250 0 1 5050
box -6 -8 106 248
use NAND2X1  _10652_
timestamp 0
transform -1 0 15150 0 -1 5050
box -6 -8 86 248
use OAI21X1  _10653_
timestamp 0
transform -1 0 15290 0 -1 5050
box -6 -8 106 248
use OAI21X1  _10654_
timestamp 0
transform -1 0 11830 0 -1 5530
box -6 -8 106 248
use OAI21X1  _10655_
timestamp 0
transform -1 0 11810 0 1 5050
box -6 -8 106 248
use OAI21X1  _10656_
timestamp 0
transform 1 0 12250 0 -1 5050
box -6 -8 106 248
use OAI21X1  _10657_
timestamp 0
transform 1 0 12090 0 -1 5050
box -6 -8 106 248
use NAND2X1  _10658_
timestamp 0
transform -1 0 11970 0 -1 5530
box -6 -8 86 248
use OAI21X1  _10659_
timestamp 0
transform -1 0 12290 0 1 5530
box -6 -8 106 248
use NAND2X1  _10660_
timestamp 0
transform -1 0 13450 0 -1 5050
box -6 -8 86 248
use OAI21X1  _10661_
timestamp 0
transform -1 0 13530 0 1 5050
box -6 -8 106 248
use NAND2X1  _10662_
timestamp 0
transform 1 0 11790 0 1 6010
box -6 -8 86 248
use OAI21X1  _10663_
timestamp 0
transform -1 0 12030 0 1 6010
box -6 -8 106 248
use NAND2X1  _10664_
timestamp 0
transform 1 0 11710 0 -1 6010
box -6 -8 86 248
use OAI21X1  _10665_
timestamp 0
transform -1 0 11930 0 -1 6010
box -6 -8 106 248
use INVX1  _10666_
timestamp 0
transform -1 0 9810 0 -1 5530
box -6 -8 66 248
use OAI21X1  _10667_
timestamp 0
transform -1 0 11670 0 1 5050
box -6 -8 106 248
use OAI21X1  _10668_
timestamp 0
transform 1 0 11190 0 1 5050
box -6 -8 106 248
use INVX1  _10669_
timestamp 0
transform -1 0 10190 0 -1 5530
box -6 -8 66 248
use OAI21X1  _10670_
timestamp 0
transform -1 0 11070 0 -1 5050
box -6 -8 106 248
use OAI21X1  _10671_
timestamp 0
transform 1 0 10810 0 -1 5050
box -6 -8 106 248
use NAND2X1  _10672_
timestamp 0
transform -1 0 10730 0 1 5050
box -6 -8 86 248
use OAI21X1  _10673_
timestamp 0
transform -1 0 10890 0 1 5050
box -6 -8 106 248
use NAND2X1  _10674_
timestamp 0
transform -1 0 10310 0 -1 5530
box -6 -8 86 248
use OAI21X1  _10675_
timestamp 0
transform -1 0 10470 0 -1 5530
box -6 -8 106 248
use NAND2X1  _10676_
timestamp 0
transform 1 0 11070 0 1 6010
box -6 -8 86 248
use OAI21X1  _10677_
timestamp 0
transform 1 0 10930 0 1 6010
box -6 -8 106 248
use NAND2X1  _10678_
timestamp 0
transform 1 0 11170 0 -1 6010
box -6 -8 86 248
use OAI21X1  _10679_
timestamp 0
transform 1 0 11290 0 -1 6010
box -6 -8 106 248
use OAI21X1  _10680_
timestamp 0
transform -1 0 9790 0 1 4570
box -6 -8 106 248
use OAI21X1  _10681_
timestamp 0
transform -1 0 9830 0 -1 5050
box -6 -8 106 248
use OAI21X1  _10682_
timestamp 0
transform -1 0 10190 0 1 4570
box -6 -8 106 248
use OAI21X1  _10683_
timestamp 0
transform -1 0 10210 0 -1 5050
box -6 -8 106 248
use NAND2X1  _10684_
timestamp 0
transform 1 0 9390 0 -1 6010
box -6 -8 86 248
use OAI21X1  _10685_
timestamp 0
transform 1 0 9250 0 -1 6010
box -6 -8 106 248
use NAND2X1  _10686_
timestamp 0
transform -1 0 8670 0 -1 6010
box -6 -8 86 248
use OAI21X1  _10687_
timestamp 0
transform -1 0 8830 0 -1 6010
box -6 -8 106 248
use DFFPOSX1  _10688_
timestamp 0
transform -1 0 12830 0 1 6010
box -6 -8 246 248
use DFFPOSX1  _10689_
timestamp 0
transform -1 0 12670 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _10690_
timestamp 0
transform 1 0 7410 0 -1 11290
box -6 -8 246 248
use DFFPOSX1  _10691_
timestamp 0
transform -1 0 13190 0 1 6010
box -6 -8 246 248
use DFFPOSX1  _10692_
timestamp 0
transform -1 0 13550 0 1 6010
box -6 -8 246 248
use DFFPOSX1  _10693_
timestamp 0
transform -1 0 13950 0 -1 6490
box -6 -8 246 248
use DFFPOSX1  _10694_
timestamp 0
transform -1 0 13290 0 -1 6490
box -6 -8 246 248
use DFFPOSX1  _10695_
timestamp 0
transform -1 0 14410 0 1 6490
box -6 -8 246 248
use DFFPOSX1  _10696_
timestamp 0
transform -1 0 13490 0 1 6490
box -6 -8 246 248
use DFFPOSX1  _10697_
timestamp 0
transform -1 0 14010 0 1 6490
box -6 -8 246 248
use DFFPOSX1  _10698_
timestamp 0
transform -1 0 13510 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _10699_
timestamp 0
transform -1 0 14450 0 -1 6490
box -6 -8 246 248
use DFFPOSX1  _10700_
timestamp 0
transform -1 0 12430 0 1 6490
box -6 -8 246 248
use DFFPOSX1  _10701_
timestamp 0
transform -1 0 11910 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _10702_
timestamp 0
transform -1 0 10790 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _10703_
timestamp 0
transform -1 0 11390 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _10704_
timestamp 0
transform 1 0 11610 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _10705_
timestamp 0
transform 1 0 12050 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _10706_
timestamp 0
transform -1 0 12050 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _10707_
timestamp 0
transform 1 0 11090 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _10708_
timestamp 0
transform -1 0 12790 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _10709_
timestamp 0
transform -1 0 13690 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _10710_
timestamp 0
transform -1 0 12990 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _10711_
timestamp 0
transform -1 0 13070 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _10712_
timestamp 0
transform -1 0 12070 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _10713_
timestamp 0
transform -1 0 10430 0 1 6010
box -6 -8 246 248
use DFFPOSX1  _10714_
timestamp 0
transform 1 0 9010 0 1 6010
box -6 -8 246 248
use DFFPOSX1  _10715_
timestamp 0
transform 1 0 9210 0 1 5050
box -6 -8 246 248
use DFFPOSX1  _10716_
timestamp 0
transform -1 0 9810 0 1 6010
box -6 -8 246 248
use DFFPOSX1  _10717_
timestamp 0
transform -1 0 11350 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _10718_
timestamp 0
transform -1 0 10750 0 1 7450
box -6 -8 246 248
use DFFPOSX1  _10719_
timestamp 0
transform 1 0 9350 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _10720_
timestamp 0
transform 1 0 9190 0 1 6490
box -6 -8 246 248
use DFFPOSX1  _10721_
timestamp 0
transform -1 0 11330 0 -1 7450
box -6 -8 246 248
use DFFPOSX1  _10722_
timestamp 0
transform 1 0 11410 0 1 7450
box -6 -8 246 248
use DFFPOSX1  _10723_
timestamp 0
transform -1 0 12150 0 1 6970
box -6 -8 246 248
use DFFPOSX1  _10724_
timestamp 0
transform -1 0 12570 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _10725_
timestamp 0
transform 1 0 16590 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _10726_
timestamp 0
transform -1 0 16070 0 -1 17050
box -6 -8 246 248
use DFFPOSX1  _10727_
timestamp 0
transform 1 0 11470 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _10728_
timestamp 0
transform 1 0 12330 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _10729_
timestamp 0
transform 1 0 12930 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _10730_
timestamp 0
transform 1 0 11670 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _10731_
timestamp 0
transform 1 0 13170 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _10732_
timestamp 0
transform 1 0 13830 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _10733_
timestamp 0
transform 1 0 12190 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _10734_
timestamp 0
transform 1 0 11990 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _10735_
timestamp 0
transform 1 0 12710 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _10736_
timestamp 0
transform 1 0 13750 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _10737_
timestamp 0
transform 1 0 16550 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _10738_
timestamp 0
transform 1 0 16430 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _10739_
timestamp 0
transform 1 0 11710 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _10740_
timestamp 0
transform 1 0 12510 0 1 5050
box -6 -8 246 248
use DFFPOSX1  _10741_
timestamp 0
transform 1 0 12130 0 -1 5530
box -6 -8 246 248
use DFFPOSX1  _10742_
timestamp 0
transform 1 0 13030 0 1 5050
box -6 -8 246 248
use DFFPOSX1  _10743_
timestamp 0
transform -1 0 15190 0 1 5050
box -6 -8 246 248
use DFFPOSX1  _10744_
timestamp 0
transform 1 0 15290 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _10745_
timestamp 0
transform 1 0 11470 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _10746_
timestamp 0
transform 1 0 12350 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _10747_
timestamp 0
transform 1 0 12290 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _10748_
timestamp 0
transform 1 0 13530 0 1 5050
box -6 -8 246 248
use DFFPOSX1  _10749_
timestamp 0
transform 1 0 11590 0 1 6490
box -6 -8 246 248
use DFFPOSX1  _10750_
timestamp 0
transform 1 0 11930 0 -1 6010
box -6 -8 246 248
use DFFPOSX1  _10751_
timestamp 0
transform 1 0 11290 0 1 5050
box -6 -8 246 248
use DFFPOSX1  _10752_
timestamp 0
transform 1 0 10530 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _10753_
timestamp 0
transform -1 0 11130 0 1 5050
box -6 -8 246 248
use DFFPOSX1  _10754_
timestamp 0
transform -1 0 10570 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _10755_
timestamp 0
transform -1 0 10890 0 1 6010
box -6 -8 246 248
use DFFPOSX1  _10756_
timestamp 0
transform -1 0 11490 0 1 6010
box -6 -8 246 248
use DFFPOSX1  _10757_
timestamp 0
transform -1 0 9690 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _10758_
timestamp 0
transform 1 0 9830 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _10759_
timestamp 0
transform 1 0 9030 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _10760_
timestamp 0
transform 1 0 8370 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _10761_
timestamp 0
transform 1 0 7690 0 1 6010
box -6 -8 246 248
use DFFPOSX1  _10762_
timestamp 0
transform -1 0 9750 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _10763_
timestamp 0
transform 1 0 9230 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _10764_
timestamp 0
transform 1 0 9470 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _10765_
timestamp 0
transform 1 0 9710 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _10766_
timestamp 0
transform 1 0 9950 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _10767_
timestamp 0
transform 1 0 10190 0 1 4090
box -6 -8 246 248
use INVX1  _10768_
timestamp 0
transform -1 0 5730 0 1 11290
box -6 -8 66 248
use INVX2  _10769_
timestamp 0
transform -1 0 4930 0 -1 13210
box -6 -8 66 248
use NOR2X1  _10770_
timestamp 0
transform -1 0 4830 0 -1 13690
box -6 -8 86 248
use INVX2  _10771_
timestamp 0
transform -1 0 5590 0 -1 13690
box -6 -8 66 248
use NOR2X1  _10772_
timestamp 0
transform 1 0 5670 0 -1 12250
box -6 -8 86 248
use INVX4  _10773_
timestamp 0
transform -1 0 4450 0 -1 13690
box -6 -8 86 248
use NOR2X1  _10774_
timestamp 0
transform 1 0 5590 0 1 13210
box -6 -8 86 248
use OAI21X1  _10775_
timestamp 0
transform 1 0 5590 0 1 12250
box -6 -8 106 248
use INVX2  _10776_
timestamp 0
transform -1 0 2750 0 -1 12250
box -6 -8 66 248
use AND2X2  _10777_
timestamp 0
transform 1 0 5470 0 -1 13210
box -6 -8 106 248
use AOI22X1  _10778_
timestamp 0
transform 1 0 5950 0 -1 12250
box -6 -8 126 248
use OAI21X1  _10779_
timestamp 0
transform 1 0 5810 0 -1 12250
box -6 -8 106 248
use NOR2X1  _10780_
timestamp 0
transform -1 0 4630 0 -1 12730
box -6 -8 86 248
use AOI22X1  _10781_
timestamp 0
transform -1 0 5950 0 1 11770
box -6 -8 126 248
use OAI21X1  _10782_
timestamp 0
transform 1 0 5470 0 -1 11770
box -6 -8 106 248
use INVX1  _10783_
timestamp 0
transform 1 0 5130 0 -1 12250
box -6 -8 66 248
use OAI21X1  _10784_
timestamp 0
transform 1 0 5370 0 -1 12250
box -6 -8 106 248
use AOI21X1  _10785_
timestamp 0
transform 1 0 5510 0 -1 12250
box -6 -8 106 248
use INVX1  _10786_
timestamp 0
transform -1 0 6830 0 1 11290
box -6 -8 66 248
use NAND2X1  _10787_
timestamp 0
transform -1 0 5690 0 -1 13210
box -6 -8 86 248
use OAI21X1  _10788_
timestamp 0
transform -1 0 6230 0 -1 12250
box -6 -8 106 248
use OAI21X1  _10789_
timestamp 0
transform 1 0 6270 0 -1 12250
box -6 -8 106 248
use AOI22X1  _10790_
timestamp 0
transform 1 0 6490 0 1 11770
box -6 -8 126 248
use NAND2X1  _10791_
timestamp 0
transform 1 0 6670 0 1 11770
box -6 -8 86 248
use INVX1  _10792_
timestamp 0
transform -1 0 5970 0 1 14170
box -6 -8 66 248
use OAI21X1  _10793_
timestamp 0
transform -1 0 5430 0 1 13690
box -6 -8 106 248
use AOI21X1  _10794_
timestamp 0
transform 1 0 5470 0 1 13690
box -6 -8 106 248
use INVX1  _10795_
timestamp 0
transform 1 0 5850 0 -1 14650
box -6 -8 66 248
use NAND2X1  _10796_
timestamp 0
transform 1 0 6190 0 -1 14170
box -6 -8 86 248
use OAI21X1  _10797_
timestamp 0
transform 1 0 6030 0 -1 14170
box -6 -8 106 248
use OAI21X1  _10798_
timestamp 0
transform 1 0 5630 0 1 13690
box -6 -8 106 248
use AOI22X1  _10799_
timestamp 0
transform 1 0 5150 0 1 13690
box -6 -8 126 248
use NAND2X1  _10800_
timestamp 0
transform 1 0 6350 0 -1 13690
box -6 -8 86 248
use INVX1  _10801_
timestamp 0
transform -1 0 5690 0 -1 15610
box -6 -8 66 248
use OAI21X1  _10802_
timestamp 0
transform -1 0 5730 0 -1 13690
box -6 -8 106 248
use AOI21X1  _10803_
timestamp 0
transform 1 0 5790 0 -1 13690
box -6 -8 106 248
use INVX1  _10804_
timestamp 0
transform -1 0 5410 0 -1 16090
box -6 -8 66 248
use NAND2X1  _10805_
timestamp 0
transform 1 0 5790 0 1 13690
box -6 -8 86 248
use OAI21X1  _10806_
timestamp 0
transform 1 0 5910 0 1 13690
box -6 -8 106 248
use OAI21X1  _10807_
timestamp 0
transform 1 0 5930 0 -1 13690
box -6 -8 106 248
use AOI22X1  _10808_
timestamp 0
transform 1 0 5130 0 -1 13690
box -6 -8 126 248
use NAND2X1  _10809_
timestamp 0
transform 1 0 6210 0 -1 13690
box -6 -8 86 248
use INVX1  _10810_
timestamp 0
transform 1 0 1130 0 -1 12250
box -6 -8 66 248
use OAI21X1  _10811_
timestamp 0
transform 1 0 1950 0 -1 12730
box -6 -8 106 248
use AOI21X1  _10812_
timestamp 0
transform 1 0 1270 0 1 12250
box -6 -8 106 248
use INVX1  _10813_
timestamp 0
transform 1 0 1570 0 1 12730
box -6 -8 66 248
use NAND2X1  _10814_
timestamp 0
transform 1 0 1570 0 1 12250
box -6 -8 86 248
use OAI21X1  _10815_
timestamp 0
transform -1 0 1530 0 1 12250
box -6 -8 106 248
use OAI21X1  _10816_
timestamp 0
transform 1 0 1690 0 1 12250
box -6 -8 106 248
use AOI22X1  _10817_
timestamp 0
transform 1 0 2810 0 -1 13210
box -6 -8 126 248
use NAND2X1  _10818_
timestamp 0
transform -1 0 2370 0 1 12250
box -6 -8 86 248
use INVX1  _10819_
timestamp 0
transform 1 0 2770 0 -1 12730
box -6 -8 66 248
use NOR2X1  _10820_
timestamp 0
transform -1 0 2110 0 -1 12250
box -6 -8 86 248
use OAI21X1  _10821_
timestamp 0
transform -1 0 2250 0 1 12250
box -6 -8 106 248
use AOI22X1  _10822_
timestamp 0
transform -1 0 1990 0 -1 12250
box -6 -8 126 248
use OAI21X1  _10823_
timestamp 0
transform 1 0 2150 0 -1 12250
box -6 -8 106 248
use AOI22X1  _10824_
timestamp 0
transform -1 0 2930 0 -1 12250
box -6 -8 126 248
use OAI21X1  _10825_
timestamp 0
transform -1 0 3070 0 -1 12250
box -6 -8 106 248
use INVX1  _10826_
timestamp 0
transform -1 0 5110 0 1 13690
box -6 -8 66 248
use INVX1  _10827_
timestamp 0
transform -1 0 5070 0 1 14170
box -6 -8 66 248
use INVX8  _10828_
timestamp 0
transform -1 0 770 0 1 15610
box -6 -8 126 248
use INVX8  _10829_
timestamp 0
transform -1 0 590 0 -1 17050
box -6 -8 126 248
use INVX1  _10830_
timestamp 0
transform -1 0 1330 0 1 13690
box -6 -8 66 248
use NAND2X1  _10831_
timestamp 0
transform 1 0 1530 0 1 13690
box -6 -8 86 248
use OAI21X1  _10832_
timestamp 0
transform 1 0 1370 0 1 13690
box -6 -8 106 248
use INVX1  _10833_
timestamp 0
transform -1 0 110 0 1 13690
box -6 -8 66 248
use NAND2X1  _10834_
timestamp 0
transform 1 0 2290 0 1 14170
box -6 -8 86 248
use OAI21X1  _10835_
timestamp 0
transform 1 0 2130 0 1 14170
box -6 -8 106 248
use MUX2X1  _10836_
timestamp 0
transform 1 0 1910 0 -1 14170
box -6 -8 126 248
use INVX1  _10837_
timestamp 0
transform 1 0 2970 0 -1 14170
box -6 -8 66 248
use NAND2X1  _10838_
timestamp 0
transform 1 0 3390 0 -1 14170
box -6 -8 86 248
use OAI21X1  _10839_
timestamp 0
transform 1 0 3090 0 -1 14170
box -6 -8 106 248
use INVX1  _10840_
timestamp 0
transform -1 0 1950 0 1 13210
box -6 -8 66 248
use NAND2X1  _10841_
timestamp 0
transform 1 0 3050 0 1 14170
box -6 -8 86 248
use OAI21X1  _10842_
timestamp 0
transform 1 0 2650 0 -1 14170
box -6 -8 106 248
use MUX2X1  _10843_
timestamp 0
transform -1 0 2930 0 -1 14170
box -6 -8 126 248
use MUX2X1  _10844_
timestamp 0
transform -1 0 3350 0 -1 14170
box -6 -8 126 248
use NOR2X1  _10845_
timestamp 0
transform -1 0 4810 0 -1 14170
box -6 -8 86 248
use NAND2X1  _10846_
timestamp 0
transform 1 0 4870 0 -1 14170
box -6 -8 86 248
use INVX1  _10847_
timestamp 0
transform -1 0 4630 0 1 13690
box -6 -8 66 248
use NAND2X1  _10848_
timestamp 0
transform -1 0 3270 0 1 14170
box -6 -8 86 248
use OAI21X1  _10849_
timestamp 0
transform -1 0 1550 0 -1 12730
box -6 -8 106 248
use INVX2  _10850_
timestamp 0
transform -1 0 1410 0 -1 12730
box -6 -8 66 248
use OAI21X1  _10851_
timestamp 0
transform -1 0 4530 0 1 13690
box -6 -8 106 248
use OAI21X1  _10852_
timestamp 0
transform -1 0 5010 0 1 13690
box -6 -8 106 248
use INVX8  _10853_
timestamp 0
transform 1 0 1850 0 1 12250
box -6 -8 126 248
use NAND2X1  _10854_
timestamp 0
transform -1 0 4570 0 -1 13690
box -6 -8 86 248
use NOR2X1  _10855_
timestamp 0
transform 1 0 3910 0 1 14170
box -6 -8 86 248
use MUX2X1  _10856_
timestamp 0
transform 1 0 2670 0 -1 14650
box -6 -8 126 248
use MUX2X1  _10857_
timestamp 0
transform 1 0 3110 0 -1 14650
box -6 -8 126 248
use MUX2X1  _10858_
timestamp 0
transform 1 0 3430 0 -1 14650
box -6 -8 126 248
use INVX2  _10859_
timestamp 0
transform -1 0 3030 0 1 12730
box -6 -8 66 248
use NAND2X1  _10860_
timestamp 0
transform 1 0 3610 0 -1 13690
box -6 -8 86 248
use AOI21X1  _10861_
timestamp 0
transform 1 0 3510 0 -1 14170
box -6 -8 106 248
use NAND3X1  _10862_
timestamp 0
transform 1 0 2910 0 -1 13690
box -6 -8 106 248
use NAND3X1  _10863_
timestamp 0
transform 1 0 3310 0 1 14170
box -6 -8 106 248
use NAND3X1  _10864_
timestamp 0
transform 1 0 3450 0 1 14170
box -6 -8 106 248
use OAI22X1  _10865_
timestamp 0
transform 1 0 3610 0 1 14170
box -6 -8 126 248
use INVX1  _10866_
timestamp 0
transform 1 0 4430 0 1 14170
box -6 -8 66 248
use INVX8  _10867_
timestamp 0
transform 1 0 770 0 1 15130
box -6 -8 126 248
use INVX1  _10868_
timestamp 0
transform 1 0 1750 0 1 14170
box -6 -8 66 248
use NAND2X1  _10869_
timestamp 0
transform 1 0 2010 0 1 14170
box -6 -8 86 248
use OAI21X1  _10870_
timestamp 0
transform 1 0 1870 0 1 14170
box -6 -8 106 248
use INVX1  _10871_
timestamp 0
transform -1 0 2470 0 1 14170
box -6 -8 66 248
use NAND2X1  _10872_
timestamp 0
transform -1 0 2150 0 -1 14650
box -6 -8 86 248
use OAI21X1  _10873_
timestamp 0
transform -1 0 2290 0 -1 14650
box -6 -8 106 248
use MUX2X1  _10874_
timestamp 0
transform -1 0 2410 0 1 14650
box -6 -8 126 248
use INVX1  _10875_
timestamp 0
transform -1 0 2710 0 1 15130
box -6 -8 66 248
use NAND2X1  _10876_
timestamp 0
transform 1 0 2450 0 -1 15130
box -6 -8 86 248
use OAI21X1  _10877_
timestamp 0
transform 1 0 2230 0 1 15130
box -6 -8 106 248
use INVX1  _10878_
timestamp 0
transform -1 0 3090 0 1 14650
box -6 -8 66 248
use NAND2X1  _10879_
timestamp 0
transform -1 0 2030 0 1 15130
box -6 -8 86 248
use OAI21X1  _10880_
timestamp 0
transform -1 0 2170 0 1 15130
box -6 -8 106 248
use MUX2X1  _10881_
timestamp 0
transform -1 0 2250 0 -1 15130
box -6 -8 126 248
use MUX2X1  _10882_
timestamp 0
transform -1 0 2410 0 -1 15130
box -6 -8 126 248
use NAND3X1  _10883_
timestamp 0
transform 1 0 3890 0 -1 14650
box -6 -8 106 248
use MUX2X1  _10884_
timestamp 0
transform -1 0 2470 0 -1 14650
box -6 -8 126 248
use MUX2X1  _10885_
timestamp 0
transform -1 0 2630 0 -1 14650
box -6 -8 126 248
use MUX2X1  _10886_
timestamp 0
transform 1 0 2470 0 1 14650
box -6 -8 126 248
use MUX2X1  _10887_
timestamp 0
transform -1 0 3250 0 1 14650
box -6 -8 126 248
use MUX2X1  _10888_
timestamp 0
transform 1 0 3630 0 1 14650
box -6 -8 126 248
use MUX2X1  _10889_
timestamp 0
transform 1 0 3310 0 1 14650
box -6 -8 126 248
use MUX2X1  _10890_
timestamp 0
transform 1 0 3470 0 1 14650
box -6 -8 126 248
use OAI21X1  _10891_
timestamp 0
transform -1 0 4610 0 1 14650
box -6 -8 106 248
use AOI21X1  _10892_
timestamp 0
transform 1 0 4310 0 -1 14650
box -6 -8 106 248
use INVX1  _10893_
timestamp 0
transform -1 0 4530 0 -1 14650
box -6 -8 66 248
use NAND3X1  _10894_
timestamp 0
transform 1 0 4170 0 -1 14650
box -6 -8 106 248
use AND2X2  _10895_
timestamp 0
transform 1 0 4570 0 -1 14650
box -6 -8 106 248
use OAI21X1  _10896_
timestamp 0
transform 1 0 4550 0 1 14170
box -6 -8 106 248
use OR2X2  _10897_
timestamp 0
transform 1 0 4850 0 1 14170
box -6 -8 106 248
use AOI21X1  _10898_
timestamp 0
transform -1 0 4810 0 1 14170
box -6 -8 106 248
use OAI21X1  _10899_
timestamp 0
transform -1 0 4710 0 -1 13690
box -6 -8 106 248
use INVX1  _10900_
timestamp 0
transform -1 0 8430 0 1 11290
box -6 -8 66 248
use NAND2X1  _10901_
timestamp 0
transform -1 0 7930 0 1 11290
box -6 -8 86 248
use OAI21X1  _10902_
timestamp 0
transform -1 0 8070 0 1 11290
box -6 -8 106 248
use NAND2X1  _10903_
timestamp 0
transform 1 0 5530 0 -1 14170
box -6 -8 86 248
use AOI21X1  _10904_
timestamp 0
transform 1 0 4710 0 -1 14650
box -6 -8 106 248
use MUX2X1  _10905_
timestamp 0
transform -1 0 2610 0 -1 14170
box -6 -8 126 248
use MUX2X1  _10906_
timestamp 0
transform -1 0 2750 0 1 14650
box -6 -8 126 248
use MUX2X1  _10907_
timestamp 0
transform -1 0 3910 0 1 14650
box -6 -8 126 248
use NAND2X1  _10908_
timestamp 0
transform -1 0 3690 0 -1 14650
box -6 -8 86 248
use OAI22X1  _10909_
timestamp 0
transform 1 0 3730 0 -1 14650
box -6 -8 126 248
use AOI21X1  _10910_
timestamp 0
transform 1 0 3970 0 1 14650
box -6 -8 106 248
use AOI21X1  _10911_
timestamp 0
transform 1 0 4650 0 1 14650
box -6 -8 106 248
use NAND2X1  _10912_
timestamp 0
transform 1 0 4810 0 1 14650
box -6 -8 86 248
use INVX1  _10913_
timestamp 0
transform -1 0 4310 0 1 14650
box -6 -8 66 248
use OAI21X1  _10914_
timestamp 0
transform 1 0 4030 0 -1 14650
box -6 -8 106 248
use NAND2X1  _10915_
timestamp 0
transform -1 0 4210 0 1 14650
box -6 -8 86 248
use AOI21X1  _10916_
timestamp 0
transform 1 0 4930 0 1 14650
box -6 -8 106 248
use NAND3X1  _10917_
timestamp 0
transform 1 0 5090 0 1 14650
box -6 -8 106 248
use INVX1  _10918_
timestamp 0
transform 1 0 5550 0 1 14650
box -6 -8 66 248
use OR2X2  _10919_
timestamp 0
transform -1 0 5190 0 -1 14650
box -6 -8 106 248
use NOR2X1  _10920_
timestamp 0
transform 1 0 4870 0 -1 14650
box -6 -8 86 248
use INVX1  _10921_
timestamp 0
transform 1 0 4990 0 -1 14650
box -6 -8 66 248
use OAI21X1  _10922_
timestamp 0
transform -1 0 5350 0 1 14650
box -6 -8 106 248
use AOI21X1  _10923_
timestamp 0
transform 1 0 5230 0 -1 14650
box -6 -8 106 248
use INVX2  _10924_
timestamp 0
transform -1 0 1110 0 -1 16570
box -6 -8 66 248
use OAI21X1  _10925_
timestamp 0
transform 1 0 5350 0 1 14170
box -6 -8 106 248
use OAI21X1  _10926_
timestamp 0
transform 1 0 5490 0 1 14170
box -6 -8 106 248
use INVX1  _10927_
timestamp 0
transform 1 0 5670 0 1 14650
box -6 -8 66 248
use INVX2  _10928_
timestamp 0
transform 1 0 5630 0 1 14170
box -6 -8 66 248
use OAI21X1  _10929_
timestamp 0
transform 1 0 5410 0 1 14650
box -6 -8 106 248
use INVX1  _10930_
timestamp 0
transform 1 0 5370 0 -1 15610
box -6 -8 66 248
use INVX1  _10931_
timestamp 0
transform 1 0 3690 0 1 15130
box -6 -8 66 248
use NAND3X1  _10932_
timestamp 0
transform -1 0 4450 0 1 14650
box -6 -8 106 248
use INVX1  _10933_
timestamp 0
transform 1 0 1270 0 -1 13690
box -6 -8 66 248
use NAND2X1  _10934_
timestamp 0
transform 1 0 1650 0 -1 14170
box -6 -8 86 248
use OAI21X1  _10935_
timestamp 0
transform 1 0 1490 0 -1 14170
box -6 -8 106 248
use NAND2X1  _10936_
timestamp 0
transform 1 0 1790 0 1 16090
box -6 -8 86 248
use OAI21X1  _10937_
timestamp 0
transform 1 0 1490 0 1 16090
box -6 -8 106 248
use NOR2X1  _10938_
timestamp 0
transform 1 0 1230 0 1 16090
box -6 -8 86 248
use NOR2X1  _10939_
timestamp 0
transform -1 0 3930 0 -1 15130
box -6 -8 86 248
use AOI22X1  _10940_
timestamp 0
transform -1 0 2170 0 -1 15610
box -6 -8 126 248
use OAI21X1  _10941_
timestamp 0
transform 1 0 1870 0 -1 16090
box -6 -8 106 248
use NAND3X1  _10942_
timestamp 0
transform 1 0 3390 0 -1 16090
box -6 -8 106 248
use INVX1  _10943_
timestamp 0
transform 1 0 3690 0 1 15610
box -6 -8 66 248
use INVX1  _10944_
timestamp 0
transform 1 0 3530 0 -1 16090
box -6 -8 66 248
use OAI21X1  _10945_
timestamp 0
transform -1 0 3890 0 1 15610
box -6 -8 106 248
use NAND3X1  _10946_
timestamp 0
transform 1 0 4090 0 1 15610
box -6 -8 106 248
use AOI21X1  _10947_
timestamp 0
transform 1 0 3930 0 1 15610
box -6 -8 106 248
use INVX1  _10948_
timestamp 0
transform -1 0 4610 0 1 15610
box -6 -8 66 248
use NAND2X1  _10949_
timestamp 0
transform -1 0 4730 0 1 15610
box -6 -8 86 248
use AOI21X1  _10950_
timestamp 0
transform -1 0 5170 0 -1 15610
box -6 -8 106 248
use OAI21X1  _10951_
timestamp 0
transform -1 0 5330 0 -1 15610
box -6 -8 106 248
use AOI22X1  _10952_
timestamp 0
transform -1 0 5510 0 -1 15130
box -6 -8 126 248
use AOI21X1  _10953_
timestamp 0
transform -1 0 4890 0 1 15610
box -6 -8 106 248
use INVX1  _10954_
timestamp 0
transform -1 0 4590 0 -1 15130
box -6 -8 66 248
use INVX1  _10955_
timestamp 0
transform -1 0 1850 0 -1 14170
box -6 -8 66 248
use NAND2X1  _10956_
timestamp 0
transform -1 0 1530 0 -1 16090
box -6 -8 86 248
use OAI21X1  _10957_
timestamp 0
transform -1 0 1670 0 -1 16090
box -6 -8 106 248
use NAND2X1  _10958_
timestamp 0
transform 1 0 1730 0 -1 16090
box -6 -8 86 248
use OAI21X1  _10959_
timestamp 0
transform 1 0 1630 0 1 16090
box -6 -8 106 248
use NAND2X1  _10960_
timestamp 0
transform 1 0 3330 0 -1 15130
box -6 -8 86 248
use OAI21X1  _10961_
timestamp 0
transform 1 0 2410 0 -1 16090
box -6 -8 106 248
use INVX2  _10962_
timestamp 0
transform 1 0 2790 0 -1 16570
box -6 -8 66 248
use OAI21X1  _10963_
timestamp 0
transform 1 0 3670 0 1 16090
box -6 -8 106 248
use OR2X2  _10964_
timestamp 0
transform 1 0 3970 0 1 16090
box -6 -8 106 248
use NOR2X1  _10965_
timestamp 0
transform -1 0 3490 0 -1 16570
box -6 -8 86 248
use OAI21X1  _10966_
timestamp 0
transform 1 0 3530 0 -1 16570
box -6 -8 106 248
use NAND3X1  _10967_
timestamp 0
transform 1 0 4450 0 1 16090
box -6 -8 106 248
use NOR2X1  _10968_
timestamp 0
transform 1 0 3770 0 -1 16090
box -6 -8 86 248
use AND2X2  _10969_
timestamp 0
transform -1 0 3730 0 -1 16090
box -6 -8 106 248
use OAI21X1  _10970_
timestamp 0
transform 1 0 3910 0 -1 16090
box -6 -8 106 248
use NAND2X1  _10971_
timestamp 0
transform -1 0 4830 0 1 16090
box -6 -8 86 248
use AOI21X1  _10972_
timestamp 0
transform 1 0 4930 0 -1 16090
box -6 -8 106 248
use OAI21X1  _10973_
timestamp 0
transform 1 0 5070 0 -1 16090
box -6 -8 106 248
use AOI22X1  _10974_
timestamp 0
transform -1 0 5910 0 1 14650
box -6 -8 126 248
use OAI21X1  _10975_
timestamp 0
transform -1 0 5110 0 1 16090
box -6 -8 106 248
use INVX1  _10976_
timestamp 0
transform -1 0 4190 0 1 15130
box -6 -8 66 248
use NAND3X1  _10977_
timestamp 0
transform 1 0 3830 0 1 16090
box -6 -8 106 248
use NAND2X1  _10978_
timestamp 0
transform 1 0 1150 0 -1 16570
box -6 -8 86 248
use INVX1  _10979_
timestamp 0
transform 1 0 1310 0 1 16570
box -6 -8 66 248
use AOI21X1  _10980_
timestamp 0
transform -1 0 1450 0 1 16090
box -6 -8 106 248
use NAND2X1  _10981_
timestamp 0
transform 1 0 2550 0 -1 16090
box -6 -8 86 248
use OAI21X1  _10982_
timestamp 0
transform 1 0 2490 0 1 16090
box -6 -8 106 248
use NAND3X1  _10983_
timestamp 0
transform 1 0 3830 0 -1 16570
box -6 -8 106 248
use NOR3X1  _10984_
timestamp 0
transform 1 0 2910 0 -1 16570
box -6 -8 186 248
use INVX1  _10985_
timestamp 0
transform -1 0 3190 0 -1 16570
box -6 -8 66 248
use OAI21X1  _10986_
timestamp 0
transform 1 0 3250 0 -1 16570
box -6 -8 106 248
use NAND3X1  _10987_
timestamp 0
transform 1 0 4110 0 -1 16570
box -6 -8 106 248
use AOI21X1  _10988_
timestamp 0
transform 1 0 4250 0 -1 16570
box -6 -8 106 248
use INVX1  _10989_
timestamp 0
transform 1 0 4890 0 1 16570
box -6 -8 66 248
use NAND2X1  _10990_
timestamp 0
transform 1 0 5090 0 -1 16570
box -6 -8 86 248
use AND2X2  _10991_
timestamp 0
transform 1 0 5170 0 1 16090
box -6 -8 106 248
use OAI21X1  _10992_
timestamp 0
transform 1 0 5310 0 1 16090
box -6 -8 106 248
use OAI21X1  _10993_
timestamp 0
transform 1 0 5470 0 1 16090
box -6 -8 106 248
use OAI21X1  _10994_
timestamp 0
transform 1 0 5450 0 -1 16090
box -6 -8 106 248
use INVX1  _10995_
timestamp 0
transform -1 0 6010 0 -1 15130
box -6 -8 66 248
use INVX1  _10996_
timestamp 0
transform 1 0 1990 0 1 16570
box -6 -8 66 248
use NAND3X1  _10997_
timestamp 0
transform -1 0 3290 0 1 16570
box -6 -8 106 248
use AOI21X1  _10998_
timestamp 0
transform -1 0 1390 0 -1 16570
box -6 -8 106 248
use NAND2X1  _10999_
timestamp 0
transform -1 0 3030 0 -1 15130
box -6 -8 86 248
use OAI21X1  _11000_
timestamp 0
transform -1 0 2330 0 -1 16570
box -6 -8 106 248
use NAND3X1  _11001_
timestamp 0
transform 1 0 2530 0 -1 17050
box -6 -8 106 248
use INVX1  _11002_
timestamp 0
transform 1 0 2670 0 -1 17050
box -6 -8 66 248
use OAI21X1  _11003_
timestamp 0
transform -1 0 3790 0 -1 16570
box -6 -8 106 248
use NAND2X1  _11004_
timestamp 0
transform 1 0 3210 0 -1 17050
box -6 -8 86 248
use NAND3X1  _11005_
timestamp 0
transform 1 0 2930 0 -1 17050
box -6 -8 106 248
use NAND3X1  _11006_
timestamp 0
transform 1 0 2770 0 -1 17050
box -6 -8 106 248
use NAND2X1  _11007_
timestamp 0
transform 1 0 3330 0 1 16570
box -6 -8 86 248
use NAND3X1  _11008_
timestamp 0
transform 1 0 3470 0 1 16570
box -6 -8 106 248
use NAND2X1  _11009_
timestamp 0
transform 1 0 3910 0 -1 17050
box -6 -8 86 248
use AOI21X1  _11010_
timestamp 0
transform 1 0 4290 0 1 16090
box -6 -8 106 248
use NOR2X1  _11011_
timestamp 0
transform -1 0 4470 0 -1 16570
box -6 -8 86 248
use OAI21X1  _11012_
timestamp 0
transform -1 0 4710 0 1 16090
box -6 -8 106 248
use NAND2X1  _11013_
timestamp 0
transform -1 0 4730 0 -1 16570
box -6 -8 86 248
use AOI21X1  _11014_
timestamp 0
transform 1 0 5210 0 -1 16570
box -6 -8 106 248
use OAI21X1  _11015_
timestamp 0
transform 1 0 5370 0 -1 16570
box -6 -8 106 248
use AOI22X1  _11016_
timestamp 0
transform -1 0 5910 0 -1 15130
box -6 -8 126 248
use INVX1  _11017_
timestamp 0
transform 1 0 5770 0 1 15610
box -6 -8 66 248
use AOI21X1  _11018_
timestamp 0
transform 1 0 3070 0 -1 17050
box -6 -8 106 248
use AND2X2  _11019_
timestamp 0
transform 1 0 4870 0 1 16090
box -6 -8 106 248
use NAND3X1  _11020_
timestamp 0
transform -1 0 5050 0 -1 16570
box -6 -8 106 248
use AOI21X1  _11021_
timestamp 0
transform 1 0 4510 0 -1 16570
box -6 -8 106 248
use OAI21X1  _11022_
timestamp 0
transform -1 0 4890 0 -1 16570
box -6 -8 106 248
use AOI21X1  _11023_
timestamp 0
transform -1 0 3870 0 -1 17050
box -6 -8 106 248
use INVX1  _11024_
timestamp 0
transform -1 0 1370 0 -1 17050
box -6 -8 66 248
use NAND3X1  _11025_
timestamp 0
transform -1 0 3150 0 1 16570
box -6 -8 106 248
use INVX1  _11026_
timestamp 0
transform -1 0 2170 0 1 15610
box -6 -8 66 248
use NOR2X1  _11027_
timestamp 0
transform -1 0 2250 0 -1 16090
box -6 -8 86 248
use INVX1  _11028_
timestamp 0
transform -1 0 2110 0 1 16090
box -6 -8 66 248
use OAI21X1  _11029_
timestamp 0
transform -1 0 1550 0 -1 16570
box -6 -8 106 248
use NAND3X1  _11030_
timestamp 0
transform -1 0 1670 0 -1 17050
box -6 -8 106 248
use INVX1  _11031_
timestamp 0
transform 1 0 1710 0 -1 17050
box -6 -8 66 248
use OAI21X1  _11032_
timestamp 0
transform -1 0 2470 0 -1 17050
box -6 -8 106 248
use NAND2X1  _11033_
timestamp 0
transform 1 0 1810 0 -1 17050
box -6 -8 86 248
use NAND3X1  _11034_
timestamp 0
transform 1 0 1430 0 -1 17050
box -6 -8 106 248
use NAND3X1  _11035_
timestamp 0
transform 1 0 1930 0 -1 17050
box -6 -8 106 248
use NAND2X1  _11036_
timestamp 0
transform 1 0 2230 0 -1 17050
box -6 -8 86 248
use NAND3X1  _11037_
timestamp 0
transform 1 0 2070 0 -1 17050
box -6 -8 106 248
use NAND2X1  _11038_
timestamp 0
transform 1 0 4030 0 -1 17050
box -6 -8 86 248
use INVX1  _11039_
timestamp 0
transform 1 0 4290 0 -1 17050
box -6 -8 66 248
use NOR2X1  _11040_
timestamp 0
transform -1 0 4230 0 -1 17050
box -6 -8 86 248
use OAI21X1  _11041_
timestamp 0
transform -1 0 4690 0 1 16570
box -6 -8 106 248
use OAI21X1  _11042_
timestamp 0
transform 1 0 4730 0 1 16570
box -6 -8 106 248
use OAI21X1  _11043_
timestamp 0
transform 1 0 5270 0 1 15130
box -6 -8 106 248
use INVX1  _11044_
timestamp 0
transform 1 0 5410 0 1 15130
box -6 -8 66 248
use OAI21X1  _11045_
timestamp 0
transform 1 0 5210 0 -1 16090
box -6 -8 106 248
use OAI21X1  _11046_
timestamp 0
transform -1 0 5470 0 1 15610
box -6 -8 106 248
use INVX1  _11047_
timestamp 0
transform -1 0 5730 0 1 15130
box -6 -8 66 248
use OAI21X1  _11048_
timestamp 0
transform -1 0 4270 0 1 16570
box -6 -8 106 248
use NOR2X1  _11049_
timestamp 0
transform 1 0 4450 0 1 16570
box -6 -8 86 248
use AOI21X1  _11050_
timestamp 0
transform -1 0 4410 0 1 16570
box -6 -8 106 248
use INVX1  _11051_
timestamp 0
transform -1 0 2870 0 1 16570
box -6 -8 66 248
use OR2X2  _11052_
timestamp 0
transform 1 0 2210 0 1 16570
box -6 -8 106 248
use OAI21X1  _11053_
timestamp 0
transform -1 0 1710 0 -1 16570
box -6 -8 106 248
use NAND3X1  _11054_
timestamp 0
transform 1 0 2350 0 1 16570
box -6 -8 106 248
use NOR2X1  _11055_
timestamp 0
transform -1 0 2070 0 -1 16570
box -6 -8 86 248
use INVX1  _11056_
timestamp 0
transform 1 0 2370 0 -1 16570
box -6 -8 66 248
use OAI21X1  _11057_
timestamp 0
transform 1 0 2630 0 -1 16570
box -6 -8 106 248
use NAND3X1  _11058_
timestamp 0
transform -1 0 2750 0 1 16570
box -6 -8 106 248
use NAND3X1  _11059_
timestamp 0
transform 1 0 2490 0 1 16570
box -6 -8 106 248
use OAI21X1  _11060_
timestamp 0
transform -1 0 2590 0 -1 16570
box -6 -8 106 248
use NAND3X1  _11061_
timestamp 0
transform 1 0 2910 0 1 16570
box -6 -8 106 248
use AND2X2  _11062_
timestamp 0
transform -1 0 3990 0 1 16570
box -6 -8 106 248
use INVX1  _11063_
timestamp 0
transform 1 0 4950 0 1 15610
box -6 -8 66 248
use AOI21X1  _11064_
timestamp 0
transform 1 0 5050 0 1 15610
box -6 -8 106 248
use OAI21X1  _11065_
timestamp 0
transform 1 0 5210 0 1 15610
box -6 -8 106 248
use AOI22X1  _11066_
timestamp 0
transform -1 0 5630 0 1 15130
box -6 -8 126 248
use NAND2X1  _11067_
timestamp 0
transform -1 0 3430 0 -1 17050
box -6 -8 86 248
use AND2X2  _11068_
timestamp 0
transform 1 0 3610 0 1 16570
box -6 -8 106 248
use AND2X2  _11069_
timestamp 0
transform -1 0 3570 0 -1 17050
box -6 -8 106 248
use NAND3X1  _11070_
timestamp 0
transform 1 0 3630 0 -1 17050
box -6 -8 106 248
use OAI21X1  _11071_
timestamp 0
transform -1 0 3850 0 1 16570
box -6 -8 106 248
use INVX1  _11072_
timestamp 0
transform -1 0 4110 0 1 16570
box -6 -8 66 248
use AOI21X1  _11073_
timestamp 0
transform 1 0 3970 0 -1 16570
box -6 -8 106 248
use INVX1  _11074_
timestamp 0
transform 1 0 3290 0 1 16090
box -6 -8 66 248
use NOR3X1  _11075_
timestamp 0
transform 1 0 1750 0 -1 16570
box -6 -8 186 248
use INVX1  _11076_
timestamp 0
transform 1 0 2970 0 -1 16090
box -6 -8 66 248
use OAI21X1  _11077_
timestamp 0
transform -1 0 2430 0 1 16090
box -6 -8 106 248
use NAND3X1  _11078_
timestamp 0
transform 1 0 3130 0 1 16090
box -6 -8 106 248
use INVX1  _11079_
timestamp 0
transform 1 0 2650 0 1 16090
box -6 -8 66 248
use OAI21X1  _11080_
timestamp 0
transform 1 0 2850 0 1 16090
box -6 -8 106 248
use NAND3X1  _11081_
timestamp 0
transform 1 0 3530 0 1 16090
box -6 -8 106 248
use NAND3X1  _11082_
timestamp 0
transform 1 0 3090 0 -1 16090
box -6 -8 106 248
use OAI21X1  _11083_
timestamp 0
transform 1 0 2990 0 1 16090
box -6 -8 106 248
use NAND3X1  _11084_
timestamp 0
transform 1 0 3250 0 -1 16090
box -6 -8 106 248
use AND2X2  _11085_
timestamp 0
transform 1 0 4050 0 -1 16090
box -6 -8 106 248
use AND2X2  _11086_
timestamp 0
transform 1 0 4490 0 -1 16090
box -6 -8 106 248
use OAI21X1  _11087_
timestamp 0
transform 1 0 4630 0 -1 16090
box -6 -8 106 248
use OAI21X1  _11088_
timestamp 0
transform 1 0 4770 0 -1 16090
box -6 -8 106 248
use OAI21X1  _11089_
timestamp 0
transform -1 0 5590 0 -1 15610
box -6 -8 106 248
use INVX1  _11090_
timestamp 0
transform -1 0 3850 0 1 15130
box -6 -8 66 248
use OAI21X1  _11091_
timestamp 0
transform 1 0 2170 0 1 16090
box -6 -8 106 248
use INVX1  _11092_
timestamp 0
transform 1 0 2750 0 1 16090
box -6 -8 66 248
use AOI21X1  _11093_
timestamp 0
transform 1 0 2670 0 -1 16090
box -6 -8 106 248
use NAND3X1  _11094_
timestamp 0
transform 1 0 2830 0 -1 16090
box -6 -8 106 248
use NAND2X1  _11095_
timestamp 0
transform -1 0 3070 0 1 15610
box -6 -8 86 248
use NAND2X1  _11096_
timestamp 0
transform -1 0 3630 0 1 15610
box -6 -8 86 248
use OAI21X1  _11097_
timestamp 0
transform 1 0 3670 0 -1 15610
box -6 -8 106 248
use NAND2X1  _11098_
timestamp 0
transform -1 0 4050 0 -1 15610
box -6 -8 86 248
use INVX1  _11099_
timestamp 0
transform 1 0 3570 0 -1 15610
box -6 -8 66 248
use AND2X2  _11100_
timestamp 0
transform 1 0 3110 0 1 15610
box -6 -8 106 248
use NAND2X1  _11101_
timestamp 0
transform -1 0 3530 0 -1 15610
box -6 -8 86 248
use NAND3X1  _11102_
timestamp 0
transform 1 0 3810 0 -1 15610
box -6 -8 106 248
use NAND2X1  _11103_
timestamp 0
transform -1 0 4470 0 -1 15610
box -6 -8 86 248
use AOI21X1  _11104_
timestamp 0
transform 1 0 3390 0 1 16090
box -6 -8 106 248
use AOI21X1  _11105_
timestamp 0
transform 1 0 4130 0 1 16090
box -6 -8 106 248
use NAND3X1  _11106_
timestamp 0
transform 1 0 4330 0 -1 16090
box -6 -8 106 248
use AOI21X1  _11107_
timestamp 0
transform 1 0 4390 0 1 15610
box -6 -8 106 248
use AND2X2  _11108_
timestamp 0
transform 1 0 4530 0 -1 15610
box -6 -8 106 248
use NAND3X1  _11109_
timestamp 0
transform 1 0 4190 0 -1 16090
box -6 -8 106 248
use OAI21X1  _11110_
timestamp 0
transform 1 0 4250 0 1 15610
box -6 -8 106 248
use OAI21X1  _11111_
timestamp 0
transform 1 0 4930 0 -1 15610
box -6 -8 106 248
use OR2X2  _11112_
timestamp 0
transform 1 0 5110 0 1 15130
box -6 -8 106 248
use AOI22X1  _11113_
timestamp 0
transform -1 0 5870 0 1 14170
box -6 -8 126 248
use NAND2X1  _11114_
timestamp 0
transform -1 0 6170 0 1 14650
box -6 -8 86 248
use INVX1  _11115_
timestamp 0
transform 1 0 4690 0 -1 15610
box -6 -8 66 248
use NAND2X1  _11116_
timestamp 0
transform -1 0 2690 0 -1 15610
box -6 -8 86 248
use INVX1  _11117_
timestamp 0
transform -1 0 2530 0 1 15610
box -6 -8 66 248
use NAND2X1  _11118_
timestamp 0
transform -1 0 2070 0 1 15610
box -6 -8 86 248
use NAND2X1  _11119_
timestamp 0
transform -1 0 2570 0 -1 15610
box -6 -8 86 248
use INVX1  _11120_
timestamp 0
transform -1 0 3110 0 1 15130
box -6 -8 66 248
use NAND2X1  _11121_
timestamp 0
transform 1 0 3150 0 1 15130
box -6 -8 86 248
use NAND2X1  _11122_
timestamp 0
transform 1 0 3310 0 -1 15610
box -6 -8 86 248
use NAND2X1  _11123_
timestamp 0
transform 1 0 3270 0 1 15130
box -6 -8 86 248
use INVX1  _11124_
timestamp 0
transform 1 0 4470 0 1 15130
box -6 -8 66 248
use NOR3X1  _11125_
timestamp 0
transform 1 0 4590 0 1 15130
box -6 -8 186 248
use AOI21X1  _11126_
timestamp 0
transform -1 0 4890 0 -1 15610
box -6 -8 106 248
use OAI21X1  _11127_
timestamp 0
transform 1 0 4830 0 1 15130
box -6 -8 106 248
use OAI21X1  _11128_
timestamp 0
transform 1 0 4970 0 1 15130
box -6 -8 106 248
use NAND2X1  _11129_
timestamp 0
transform -1 0 6050 0 1 14650
box -6 -8 86 248
use NAND2X1  _11130_
timestamp 0
transform 1 0 2010 0 -1 13690
box -6 -8 86 248
use INVX1  _11131_
timestamp 0
transform -1 0 3510 0 -1 15130
box -6 -8 66 248
use NAND2X1  _11132_
timestamp 0
transform 1 0 3550 0 1 15130
box -6 -8 86 248
use OAI21X1  _11133_
timestamp 0
transform -1 0 3490 0 1 15130
box -6 -8 106 248
use NAND2X1  _11134_
timestamp 0
transform 1 0 2370 0 -1 15610
box -6 -8 86 248
use NOR2X1  _11135_
timestamp 0
transform -1 0 4170 0 -1 14170
box -6 -8 86 248
use NOR2X1  _11136_
timestamp 0
transform 1 0 3750 0 1 12730
box -6 -8 86 248
use AOI22X1  _11137_
timestamp 0
transform -1 0 4390 0 1 14170
box -6 -8 126 248
use NAND3X1  _11138_
timestamp 0
transform -1 0 2310 0 -1 15610
box -6 -8 106 248
use NAND2X1  _11139_
timestamp 0
transform 1 0 1170 0 -1 17050
box -6 -8 86 248
use OAI21X1  _11140_
timestamp 0
transform 1 0 1010 0 -1 17050
box -6 -8 106 248
use NAND2X1  _11141_
timestamp 0
transform -1 0 4190 0 -1 15610
box -6 -8 86 248
use OAI21X1  _11142_
timestamp 0
transform -1 0 4330 0 -1 15610
box -6 -8 106 248
use MUX2X1  _11143_
timestamp 0
transform 1 0 750 0 1 16570
box -6 -8 126 248
use NAND2X1  _11144_
timestamp 0
transform 1 0 190 0 -1 16570
box -6 -8 86 248
use AND2X2  _11145_
timestamp 0
transform -1 0 1570 0 -1 15610
box -6 -8 106 248
use NOR2X1  _11146_
timestamp 0
transform -1 0 1470 0 -1 13690
box -6 -8 86 248
use NAND2X1  _11147_
timestamp 0
transform 1 0 910 0 1 16570
box -6 -8 86 248
use NAND2X1  _11148_
timestamp 0
transform -1 0 1250 0 1 16570
box -6 -8 86 248
use NAND2X1  _11149_
timestamp 0
transform 1 0 1030 0 1 16570
box -6 -8 86 248
use OAI21X1  _11150_
timestamp 0
transform 1 0 1770 0 -1 15610
box -6 -8 106 248
use OAI21X1  _11151_
timestamp 0
transform -1 0 1770 0 1 13690
box -6 -8 106 248
use OAI21X1  _11152_
timestamp 0
transform 1 0 1630 0 -1 13690
box -6 -8 106 248
use NAND2X1  _11153_
timestamp 0
transform -1 0 2650 0 -1 12250
box -6 -8 86 248
use NOR2X1  _11154_
timestamp 0
transform -1 0 2010 0 -1 14650
box -6 -8 86 248
use NAND2X1  _11155_
timestamp 0
transform 1 0 3410 0 1 15610
box -6 -8 86 248
use OAI21X1  _11156_
timestamp 0
transform 1 0 3250 0 1 15610
box -6 -8 106 248
use NAND2X1  _11157_
timestamp 0
transform 1 0 3550 0 -1 15130
box -6 -8 86 248
use OAI21X1  _11158_
timestamp 0
transform -1 0 3790 0 -1 15130
box -6 -8 106 248
use MUX2X1  _11159_
timestamp 0
transform 1 0 1710 0 1 15610
box -6 -8 126 248
use NAND2X1  _11160_
timestamp 0
transform 1 0 490 0 1 16090
box -6 -8 86 248
use NAND2X1  _11161_
timestamp 0
transform 1 0 890 0 -1 17050
box -6 -8 86 248
use OAI21X1  _11162_
timestamp 0
transform -1 0 850 0 -1 17050
box -6 -8 106 248
use INVX1  _11163_
timestamp 0
transform -1 0 130 0 -1 17050
box -6 -8 66 248
use NAND2X1  _11164_
timestamp 0
transform 1 0 1850 0 1 16570
box -6 -8 86 248
use OAI21X1  _11165_
timestamp 0
transform 1 0 1710 0 1 16570
box -6 -8 106 248
use NAND2X1  _11166_
timestamp 0
transform 1 0 330 0 -1 17050
box -6 -8 86 248
use OAI21X1  _11167_
timestamp 0
transform 1 0 190 0 -1 17050
box -6 -8 106 248
use OAI21X1  _11168_
timestamp 0
transform 1 0 330 0 1 16090
box -6 -8 106 248
use NAND3X1  _11169_
timestamp 0
transform 1 0 1250 0 1 15130
box -6 -8 106 248
use MUX2X1  _11170_
timestamp 0
transform 1 0 590 0 -1 16570
box -6 -8 126 248
use MUX2X1  _11171_
timestamp 0
transform -1 0 870 0 -1 16570
box -6 -8 126 248
use OAI21X1  _11172_
timestamp 0
transform -1 0 1730 0 -1 15610
box -6 -8 106 248
use AOI21X1  _11173_
timestamp 0
transform 1 0 1670 0 1 15130
box -6 -8 106 248
use INVX1  _11174_
timestamp 0
transform 1 0 1870 0 -1 15130
box -6 -8 66 248
use NAND3X1  _11175_
timestamp 0
transform -1 0 1630 0 1 15130
box -6 -8 106 248
use AND2X2  _11176_
timestamp 0
transform 1 0 1970 0 -1 15130
box -6 -8 106 248
use NAND2X1  _11177_
timestamp 0
transform 1 0 1990 0 1 14650
box -6 -8 86 248
use OR2X2  _11178_
timestamp 0
transform -1 0 1930 0 1 14650
box -6 -8 106 248
use AOI21X1  _11179_
timestamp 0
transform 1 0 2130 0 1 14650
box -6 -8 106 248
use OAI21X1  _11180_
timestamp 0
transform 1 0 2410 0 -1 12250
box -6 -8 106 248
use NAND2X1  _11181_
timestamp 0
transform -1 0 2230 0 1 13210
box -6 -8 86 248
use AOI21X1  _11182_
timestamp 0
transform -1 0 1830 0 -1 15130
box -6 -8 106 248
use NAND2X1  _11183_
timestamp 0
transform 1 0 1190 0 -1 15610
box -6 -8 86 248
use NAND2X1  _11184_
timestamp 0
transform 1 0 1570 0 1 16570
box -6 -8 86 248
use OAI21X1  _11185_
timestamp 0
transform 1 0 1410 0 1 16570
box -6 -8 106 248
use NAND2X1  _11186_
timestamp 0
transform 1 0 630 0 1 16570
box -6 -8 86 248
use OAI21X1  _11187_
timestamp 0
transform -1 0 570 0 1 16570
box -6 -8 106 248
use NAND2X1  _11188_
timestamp 0
transform 1 0 1870 0 1 15610
box -6 -8 86 248
use NAND2X1  _11189_
timestamp 0
transform 1 0 1330 0 1 15610
box -6 -8 86 248
use NAND2X1  _11190_
timestamp 0
transform -1 0 1270 0 1 15610
box -6 -8 86 248
use AOI21X1  _11191_
timestamp 0
transform 1 0 930 0 1 15610
box -6 -8 106 248
use INVX1  _11192_
timestamp 0
transform 1 0 810 0 1 15610
box -6 -8 66 248
use NAND3X1  _11193_
timestamp 0
transform 1 0 910 0 -1 15610
box -6 -8 106 248
use AOI21X1  _11194_
timestamp 0
transform -1 0 1430 0 -1 15610
box -6 -8 106 248
use OAI21X1  _11195_
timestamp 0
transform -1 0 1150 0 -1 15610
box -6 -8 106 248
use NAND3X1  _11196_
timestamp 0
transform -1 0 1050 0 1 15130
box -6 -8 106 248
use INVX1  _11197_
timestamp 0
transform 1 0 1070 0 -1 15130
box -6 -8 66 248
use AOI21X1  _11198_
timestamp 0
transform 1 0 1110 0 1 15130
box -6 -8 106 248
use NOR2X1  _11199_
timestamp 0
transform 1 0 1170 0 -1 15130
box -6 -8 86 248
use AND2X2  _11200_
timestamp 0
transform 1 0 1430 0 -1 15130
box -6 -8 106 248
use NOR2X1  _11201_
timestamp 0
transform -1 0 1390 0 -1 15130
box -6 -8 86 248
use OAI21X1  _11202_
timestamp 0
transform 1 0 1570 0 -1 15130
box -6 -8 106 248
use OAI21X1  _11203_
timestamp 0
transform 1 0 2010 0 1 13210
box -6 -8 106 248
use OAI21X1  _11204_
timestamp 0
transform -1 0 1030 0 -1 15130
box -6 -8 106 248
use INVX1  _11205_
timestamp 0
transform -1 0 390 0 -1 15130
box -6 -8 66 248
use NAND2X1  _11206_
timestamp 0
transform 1 0 2030 0 -1 16090
box -6 -8 86 248
use OAI21X1  _11207_
timestamp 0
transform 1 0 1910 0 1 16090
box -6 -8 106 248
use MUX2X1  _11208_
timestamp 0
transform -1 0 750 0 1 16090
box -6 -8 126 248
use NOR2X1  _11209_
timestamp 0
transform 1 0 190 0 -1 16090
box -6 -8 86 248
use NAND2X1  _11210_
timestamp 0
transform -1 0 1670 0 1 15610
box -6 -8 86 248
use NAND2X1  _11211_
timestamp 0
transform -1 0 1410 0 -1 16090
box -6 -8 86 248
use NAND2X1  _11212_
timestamp 0
transform 1 0 1450 0 1 15610
box -6 -8 86 248
use OR2X2  _11213_
timestamp 0
transform -1 0 170 0 1 15610
box -6 -8 106 248
use OAI21X1  _11214_
timestamp 0
transform -1 0 870 0 -1 15610
box -6 -8 106 248
use OR2X2  _11215_
timestamp 0
transform 1 0 350 0 -1 15610
box -6 -8 106 248
use OAI21X1  _11216_
timestamp 0
transform 1 0 350 0 1 15610
box -6 -8 106 248
use AOI21X1  _11217_
timestamp 0
transform 1 0 610 0 1 15130
box -6 -8 106 248
use INVX1  _11218_
timestamp 0
transform -1 0 250 0 1 15130
box -6 -8 66 248
use NAND3X1  _11219_
timestamp 0
transform -1 0 550 0 1 15130
box -6 -8 106 248
use NAND2X1  _11220_
timestamp 0
transform -1 0 150 0 1 15130
box -6 -8 86 248
use OR2X2  _11221_
timestamp 0
transform 1 0 190 0 -1 15130
box -6 -8 106 248
use NAND2X1  _11222_
timestamp 0
transform -1 0 150 0 -1 15130
box -6 -8 86 248
use NAND2X1  _11223_
timestamp 0
transform 1 0 430 0 -1 15130
box -6 -8 86 248
use AOI22X1  _11224_
timestamp 0
transform -1 0 2470 0 -1 12730
box -6 -8 126 248
use AOI21X1  _11225_
timestamp 0
transform -1 0 410 0 1 15130
box -6 -8 106 248
use NAND2X1  _11226_
timestamp 0
transform -1 0 2650 0 1 15610
box -6 -8 86 248
use OAI21X1  _11227_
timestamp 0
transform -1 0 2810 0 1 15610
box -6 -8 106 248
use NAND2X1  _11228_
timestamp 0
transform -1 0 390 0 -1 16570
box -6 -8 86 248
use OAI21X1  _11229_
timestamp 0
transform -1 0 430 0 1 16570
box -6 -8 106 248
use NAND2X1  _11230_
timestamp 0
transform 1 0 50 0 1 16570
box -6 -8 86 248
use OAI21X1  _11231_
timestamp 0
transform -1 0 270 0 1 16570
box -6 -8 106 248
use INVX1  _11232_
timestamp 0
transform 1 0 370 0 1 14650
box -6 -8 66 248
use NAND3X1  _11233_
timestamp 0
transform -1 0 590 0 -1 15610
box -6 -8 106 248
use OAI21X1  _11234_
timestamp 0
transform 1 0 190 0 -1 15610
box -6 -8 106 248
use OR2X2  _11235_
timestamp 0
transform -1 0 290 0 -1 14650
box -6 -8 106 248
use NOR2X1  _11236_
timestamp 0
transform -1 0 130 0 -1 15610
box -6 -8 86 248
use OAI21X1  _11237_
timestamp 0
transform -1 0 170 0 1 14650
box -6 -8 106 248
use NAND3X1  _11238_
timestamp 0
transform -1 0 150 0 -1 14650
box -6 -8 106 248
use OR2X2  _11239_
timestamp 0
transform 1 0 350 0 -1 14650
box -6 -8 106 248
use OAI21X1  _11240_
timestamp 0
transform 1 0 210 0 1 14650
box -6 -8 106 248
use NAND3X1  _11241_
timestamp 0
transform -1 0 170 0 -1 14170
box -6 -8 106 248
use NAND2X1  _11242_
timestamp 0
transform -1 0 130 0 1 13210
box -6 -8 86 248
use OR2X2  _11243_
timestamp 0
transform 1 0 350 0 -1 13210
box -6 -8 106 248
use NAND2X1  _11244_
timestamp 0
transform -1 0 310 0 -1 13210
box -6 -8 86 248
use NAND2X1  _11245_
timestamp 0
transform -1 0 570 0 -1 13210
box -6 -8 86 248
use AOI22X1  _11246_
timestamp 0
transform -1 0 1290 0 1 12730
box -6 -8 126 248
use INVX1  _11247_
timestamp 0
transform -1 0 270 0 1 12250
box -6 -8 66 248
use OAI21X1  _11248_
timestamp 0
transform -1 0 170 0 -1 13210
box -6 -8 106 248
use NAND2X1  _11249_
timestamp 0
transform -1 0 130 0 1 14170
box -6 -8 86 248
use NOR2X1  _11250_
timestamp 0
transform 1 0 1110 0 1 16090
box -6 -8 86 248
use AOI21X1  _11251_
timestamp 0
transform -1 0 910 0 1 16090
box -6 -8 106 248
use NAND2X1  _11252_
timestamp 0
transform -1 0 130 0 1 16090
box -6 -8 86 248
use OAI21X1  _11253_
timestamp 0
transform -1 0 290 0 1 16090
box -6 -8 106 248
use INVX1  _11254_
timestamp 0
transform 1 0 490 0 -1 14650
box -6 -8 66 248
use NAND3X1  _11255_
timestamp 0
transform -1 0 410 0 1 14170
box -6 -8 106 248
use NOR2X1  _11256_
timestamp 0
transform -1 0 310 0 1 15610
box -6 -8 86 248
use NAND3X1  _11257_
timestamp 0
transform 1 0 630 0 -1 15610
box -6 -8 106 248
use OAI21X1  _11258_
timestamp 0
transform -1 0 670 0 -1 15130
box -6 -8 106 248
use NAND2X1  _11259_
timestamp 0
transform 1 0 470 0 1 14650
box -6 -8 86 248
use AOI21X1  _11260_
timestamp 0
transform -1 0 470 0 -1 14170
box -6 -8 106 248
use INVX1  _11261_
timestamp 0
transform -1 0 270 0 -1 13690
box -6 -8 66 248
use NAND3X1  _11262_
timestamp 0
transform 1 0 510 0 -1 14170
box -6 -8 106 248
use NAND2X1  _11263_
timestamp 0
transform -1 0 270 0 1 13210
box -6 -8 86 248
use NOR2X1  _11264_
timestamp 0
transform -1 0 130 0 -1 12730
box -6 -8 86 248
use AND2X2  _11265_
timestamp 0
transform 1 0 190 0 -1 12730
box -6 -8 106 248
use OAI21X1  _11266_
timestamp 0
transform 1 0 330 0 -1 12730
box -6 -8 106 248
use OAI21X1  _11267_
timestamp 0
transform -1 0 170 0 1 12250
box -6 -8 106 248
use INVX1  _11268_
timestamp 0
transform -1 0 1570 0 -1 12250
box -6 -8 66 248
use NAND3X1  _11269_
timestamp 0
transform 1 0 170 0 1 14170
box -6 -8 106 248
use AOI21X1  _11270_
timestamp 0
transform -1 0 1070 0 1 16090
box -6 -8 106 248
use NAND2X1  _11271_
timestamp 0
transform 1 0 570 0 -1 16090
box -6 -8 86 248
use OAI21X1  _11272_
timestamp 0
transform 1 0 510 0 1 15610
box -6 -8 106 248
use NAND3X1  _11273_
timestamp 0
transform 1 0 450 0 1 14170
box -6 -8 106 248
use NOR3X1  _11274_
timestamp 0
transform 1 0 710 0 -1 15130
box -6 -8 186 248
use INVX1  _11275_
timestamp 0
transform -1 0 670 0 1 14650
box -6 -8 66 248
use OAI21X1  _11276_
timestamp 0
transform -1 0 810 0 1 14650
box -6 -8 106 248
use NAND2X1  _11277_
timestamp 0
transform -1 0 550 0 1 13690
box -6 -8 86 248
use NAND2X1  _11278_
timestamp 0
transform -1 0 670 0 -1 13690
box -6 -8 86 248
use NAND3X1  _11279_
timestamp 0
transform 1 0 610 0 1 13690
box -6 -8 106 248
use NAND2X1  _11280_
timestamp 0
transform -1 0 790 0 1 13210
box -6 -8 86 248
use AOI21X1  _11281_
timestamp 0
transform 1 0 210 0 -1 14170
box -6 -8 106 248
use NOR2X1  _11282_
timestamp 0
transform -1 0 250 0 1 13690
box -6 -8 86 248
use OAI21X1  _11283_
timestamp 0
transform -1 0 410 0 1 13210
box -6 -8 106 248
use NAND2X1  _11284_
timestamp 0
transform 1 0 470 0 1 13210
box -6 -8 86 248
use NOR2X1  _11285_
timestamp 0
transform -1 0 670 0 1 13210
box -6 -8 86 248
use AND2X2  _11286_
timestamp 0
transform 1 0 730 0 -1 13210
box -6 -8 106 248
use AND2X2  _11287_
timestamp 0
transform 1 0 70 0 -1 13690
box -6 -8 106 248
use NAND3X1  _11288_
timestamp 0
transform 1 0 310 0 -1 13690
box -6 -8 106 248
use AOI21X1  _11289_
timestamp 0
transform 1 0 310 0 1 13690
box -6 -8 106 248
use OAI21X1  _11290_
timestamp 0
transform 1 0 450 0 -1 13690
box -6 -8 106 248
use NOR2X1  _11291_
timestamp 0
transform 1 0 890 0 -1 13210
box -6 -8 86 248
use OAI21X1  _11292_
timestamp 0
transform 1 0 1010 0 -1 13210
box -6 -8 106 248
use NAND2X1  _11293_
timestamp 0
transform -1 0 1310 0 -1 12250
box -6 -8 86 248
use OAI21X1  _11294_
timestamp 0
transform -1 0 1470 0 -1 12250
box -6 -8 106 248
use INVX1  _11295_
timestamp 0
transform -1 0 1290 0 -1 12730
box -6 -8 66 248
use INVX1  _11296_
timestamp 0
transform -1 0 690 0 -1 13210
box -6 -8 66 248
use NAND2X1  _11297_
timestamp 0
transform 1 0 850 0 1 14650
box -6 -8 86 248
use NOR2X1  _11298_
timestamp 0
transform -1 0 1290 0 -1 16090
box -6 -8 86 248
use INVX1  _11299_
timestamp 0
transform -1 0 1050 0 -1 16090
box -6 -8 66 248
use OAI21X1  _11300_
timestamp 0
transform 1 0 310 0 -1 16090
box -6 -8 106 248
use NAND3X1  _11301_
timestamp 0
transform 1 0 930 0 -1 14170
box -6 -8 106 248
use INVX1  _11302_
timestamp 0
transform 1 0 750 0 -1 14650
box -6 -8 66 248
use OAI21X1  _11303_
timestamp 0
transform 1 0 610 0 -1 14650
box -6 -8 106 248
use NAND2X1  _11304_
timestamp 0
transform -1 0 790 0 1 14170
box -6 -8 86 248
use NAND3X1  _11305_
timestamp 0
transform -1 0 870 0 -1 14170
box -6 -8 106 248
use NAND3X1  _11306_
timestamp 0
transform 1 0 850 0 1 14170
box -6 -8 106 248
use NAND2X1  _11307_
timestamp 0
transform -1 0 670 0 1 14170
box -6 -8 86 248
use NAND3X1  _11308_
timestamp 0
transform -1 0 1110 0 1 14170
box -6 -8 106 248
use NAND2X1  _11309_
timestamp 0
transform 1 0 750 0 1 13690
box -6 -8 86 248
use OAI21X1  _11310_
timestamp 0
transform 1 0 190 0 1 12730
box -6 -8 106 248
use NOR2X1  _11311_
timestamp 0
transform -1 0 130 0 1 12730
box -6 -8 86 248
use INVX1  _11312_
timestamp 0
transform 1 0 470 0 -1 12730
box -6 -8 66 248
use AOI21X1  _11313_
timestamp 0
transform 1 0 590 0 -1 12730
box -6 -8 106 248
use AOI22X1  _11314_
timestamp 0
transform -1 0 950 0 -1 12730
box -6 -8 126 248
use OAI21X1  _11315_
timestamp 0
transform 1 0 730 0 -1 13690
box -6 -8 106 248
use NOR2X1  _11316_
timestamp 0
transform 1 0 830 0 1 13210
box -6 -8 86 248
use AOI21X1  _11317_
timestamp 0
transform 1 0 950 0 1 13210
box -6 -8 106 248
use INVX1  _11318_
timestamp 0
transform -1 0 950 0 1 13690
box -6 -8 66 248
use NAND3X1  _11319_
timestamp 0
transform 1 0 850 0 -1 14650
box -6 -8 106 248
use INVX1  _11320_
timestamp 0
transform -1 0 130 0 -1 16570
box -6 -8 66 248
use OAI21X1  _11321_
timestamp 0
transform -1 0 150 0 -1 16090
box -6 -8 106 248
use INVX1  _11322_
timestamp 0
transform -1 0 1190 0 1 14650
box -6 -8 66 248
use NAND3X1  _11323_
timestamp 0
transform 1 0 1250 0 -1 14650
box -6 -8 106 248
use OAI21X1  _11324_
timestamp 0
transform 1 0 970 0 1 14650
box -6 -8 106 248
use NAND2X1  _11325_
timestamp 0
transform -1 0 1090 0 -1 14650
box -6 -8 86 248
use AOI21X1  _11326_
timestamp 0
transform 1 0 1070 0 -1 14170
box -6 -8 106 248
use NAND3X1  _11327_
timestamp 0
transform -1 0 1430 0 1 14170
box -6 -8 106 248
use NAND2X1  _11328_
timestamp 0
transform -1 0 1210 0 -1 14650
box -6 -8 86 248
use AOI21X1  _11329_
timestamp 0
transform 1 0 1170 0 1 14170
box -6 -8 106 248
use OAI21X1  _11330_
timestamp 0
transform -1 0 830 0 1 12730
box -6 -8 106 248
use INVX1  _11331_
timestamp 0
transform -1 0 790 0 -1 12730
box -6 -8 66 248
use OR2X2  _11332_
timestamp 0
transform 1 0 1310 0 -1 13210
box -6 -8 106 248
use OAI21X1  _11333_
timestamp 0
transform -1 0 430 0 1 12730
box -6 -8 106 248
use OAI22X1  _11334_
timestamp 0
transform -1 0 690 0 1 12250
box -6 -8 126 248
use NAND2X1  _11335_
timestamp 0
transform 1 0 890 0 1 12250
box -6 -8 86 248
use NOR2X1  _11336_
timestamp 0
transform -1 0 550 0 1 12730
box -6 -8 86 248
use NOR2X1  _11337_
timestamp 0
transform -1 0 690 0 1 12730
box -6 -8 86 248
use OAI21X1  _11338_
timestamp 0
transform 1 0 690 0 -1 16090
box -6 -8 106 248
use INVX1  _11339_
timestamp 0
transform 1 0 1410 0 -1 14650
box -6 -8 66 248
use OAI21X1  _11340_
timestamp 0
transform 1 0 1470 0 1 14170
box -6 -8 106 248
use NAND2X1  _11341_
timestamp 0
transform 1 0 1370 0 -1 14170
box -6 -8 86 248
use OR2X2  _11342_
timestamp 0
transform -1 0 1310 0 -1 14170
box -6 -8 106 248
use NAND3X1  _11343_
timestamp 0
transform -1 0 1230 0 1 13690
box -6 -8 106 248
use NAND2X1  _11344_
timestamp 0
transform -1 0 1090 0 1 13690
box -6 -8 86 248
use NAND2X1  _11345_
timestamp 0
transform -1 0 1090 0 -1 13690
box -6 -8 86 248
use NAND2X1  _11346_
timestamp 0
transform 1 0 1170 0 -1 13210
box -6 -8 86 248
use AND2X2  _11347_
timestamp 0
transform -1 0 970 0 1 12730
box -6 -8 106 248
use OAI21X1  _11348_
timestamp 0
transform 1 0 1010 0 1 12730
box -6 -8 106 248
use OAI21X1  _11349_
timestamp 0
transform -1 0 850 0 1 12250
box -6 -8 106 248
use INVX1  _11350_
timestamp 0
transform -1 0 1910 0 -1 12730
box -6 -8 66 248
use INVX1  _11351_
timestamp 0
transform -1 0 1170 0 1 13210
box -6 -8 66 248
use AOI21X1  _11352_
timestamp 0
transform 1 0 1210 0 1 13210
box -6 -8 106 248
use NOR2X1  _11353_
timestamp 0
transform -1 0 970 0 -1 13690
box -6 -8 86 248
use NAND3X1  _11354_
timestamp 0
transform 1 0 1130 0 -1 13690
box -6 -8 106 248
use OAI21X1  _11355_
timestamp 0
transform 1 0 1350 0 1 13210
box -6 -8 106 248
use OAI21X1  _11356_
timestamp 0
transform 1 0 850 0 -1 16090
box -6 -8 106 248
use INVX1  _11357_
timestamp 0
transform 1 0 1090 0 -1 16090
box -6 -8 66 248
use OR2X2  _11358_
timestamp 0
transform 1 0 1250 0 1 14650
box -6 -8 106 248
use OAI21X1  _11359_
timestamp 0
transform 1 0 1390 0 1 14650
box -6 -8 106 248
use NAND2X1  _11360_
timestamp 0
transform -1 0 1630 0 1 14650
box -6 -8 86 248
use OR2X2  _11361_
timestamp 0
transform 1 0 1510 0 -1 14650
box -6 -8 106 248
use NAND3X1  _11362_
timestamp 0
transform -1 0 1710 0 1 14170
box -6 -8 106 248
use AND2X2  _11363_
timestamp 0
transform 1 0 1690 0 1 14650
box -6 -8 106 248
use NOR2X1  _11364_
timestamp 0
transform -1 0 1730 0 -1 14650
box -6 -8 86 248
use OAI21X1  _11365_
timestamp 0
transform 1 0 1790 0 -1 14650
box -6 -8 106 248
use NAND2X1  _11366_
timestamp 0
transform -1 0 1590 0 -1 13690
box -6 -8 86 248
use AND2X2  _11367_
timestamp 0
transform 1 0 1630 0 1 13210
box -6 -8 106 248
use NOR2X1  _11368_
timestamp 0
transform -1 0 1590 0 1 13210
box -6 -8 86 248
use NOR2X1  _11369_
timestamp 0
transform 1 0 1770 0 1 13210
box -6 -8 86 248
use AOI22X1  _11370_
timestamp 0
transform -1 0 1810 0 1 12730
box -6 -8 126 248
use NAND2X1  _11371_
timestamp 0
transform -1 0 1670 0 -1 12730
box -6 -8 86 248
use INVX1  _11372_
timestamp 0
transform -1 0 1530 0 -1 13210
box -6 -8 66 248
use AOI21X1  _11373_
timestamp 0
transform 1 0 1570 0 -1 13210
box -6 -8 106 248
use NAND2X1  _11374_
timestamp 0
transform 1 0 1390 0 1 15130
box -6 -8 86 248
use NOR2X1  _11375_
timestamp 0
transform -1 0 2470 0 1 15130
box -6 -8 86 248
use AOI21X1  _11376_
timestamp 0
transform -1 0 2850 0 1 15130
box -6 -8 106 248
use NOR2X1  _11377_
timestamp 0
transform -1 0 2610 0 1 15130
box -6 -8 86 248
use AND2X2  _11378_
timestamp 0
transform 1 0 1870 0 -1 13210
box -6 -8 106 248
use OAI21X1  _11379_
timestamp 0
transform -1 0 1830 0 -1 13210
box -6 -8 106 248
use OAI21X1  _11380_
timestamp 0
transform -1 0 1810 0 -1 12730
box -6 -8 106 248
use OAI21X1  _11381_
timestamp 0
transform -1 0 2510 0 1 12250
box -6 -8 106 248
use OAI21X1  _11382_
timestamp 0
transform 1 0 4270 0 1 11770
box -6 -8 106 248
use INVX1  _11383_
timestamp 0
transform 1 0 4410 0 1 11770
box -6 -8 66 248
use NOR2X1  _11384_
timestamp 0
transform -1 0 4070 0 -1 11770
box -6 -8 86 248
use NAND2X1  _11385_
timestamp 0
transform 1 0 4510 0 1 11770
box -6 -8 86 248
use NAND2X1  _11386_
timestamp 0
transform 1 0 4770 0 1 11770
box -6 -8 86 248
use NAND2X1  _11387_
timestamp 0
transform 1 0 6010 0 1 11770
box -6 -8 86 248
use OAI21X1  _11388_
timestamp 0
transform 1 0 5430 0 1 11770
box -6 -8 106 248
use NAND2X1  _11389_
timestamp 0
transform -1 0 6210 0 -1 11290
box -6 -8 86 248
use INVX1  _11390_
timestamp 0
transform 1 0 4730 0 1 11290
box -6 -8 66 248
use NOR2X1  _11391_
timestamp 0
transform -1 0 3690 0 1 12730
box -6 -8 86 248
use AOI21X1  _11392_
timestamp 0
transform -1 0 3790 0 1 11290
box -6 -8 106 248
use NOR2X1  _11393_
timestamp 0
transform 1 0 4630 0 -1 11290
box -6 -8 86 248
use OAI21X1  _11394_
timestamp 0
transform 1 0 3830 0 -1 11770
box -6 -8 106 248
use AND2X2  _11395_
timestamp 0
transform 1 0 4750 0 -1 11290
box -6 -8 106 248
use OR2X2  _11396_
timestamp 0
transform -1 0 5010 0 -1 11290
box -6 -8 106 248
use OR2X2  _11397_
timestamp 0
transform 1 0 5190 0 -1 11290
box -6 -8 106 248
use OAI21X1  _11398_
timestamp 0
transform 1 0 5050 0 -1 11290
box -6 -8 106 248
use NAND2X1  _11399_
timestamp 0
transform 1 0 5350 0 -1 11290
box -6 -8 86 248
use NOR2X1  _11400_
timestamp 0
transform 1 0 5470 0 -1 11290
box -6 -8 86 248
use NAND2X1  _11401_
timestamp 0
transform 1 0 4990 0 1 11290
box -6 -8 86 248
use NAND2X1  _11402_
timestamp 0
transform 1 0 5830 0 -1 11290
box -6 -8 86 248
use OAI21X1  _11403_
timestamp 0
transform 1 0 5970 0 -1 11290
box -6 -8 106 248
use INVX1  _11404_
timestamp 0
transform -1 0 4690 0 1 11290
box -6 -8 66 248
use OAI21X1  _11405_
timestamp 0
transform 1 0 4830 0 1 11290
box -6 -8 106 248
use OAI21X1  _11406_
timestamp 0
transform -1 0 2910 0 1 12250
box -6 -8 106 248
use OAI21X1  _11407_
timestamp 0
transform 1 0 3290 0 -1 12250
box -6 -8 106 248
use MUX2X1  _11408_
timestamp 0
transform 1 0 3130 0 -1 12250
box -6 -8 126 248
use NAND2X1  _11409_
timestamp 0
transform -1 0 4190 0 -1 11770
box -6 -8 86 248
use OR2X2  _11410_
timestamp 0
transform 1 0 4250 0 -1 11770
box -6 -8 106 248
use NAND2X1  _11411_
timestamp 0
transform -1 0 4470 0 -1 11770
box -6 -8 86 248
use INVX1  _11412_
timestamp 0
transform 1 0 4410 0 1 11290
box -6 -8 66 248
use NOR2X1  _11413_
timestamp 0
transform 1 0 5250 0 1 11290
box -6 -8 86 248
use NAND2X1  _11414_
timestamp 0
transform -1 0 5190 0 1 11290
box -6 -8 86 248
use NAND2X1  _11415_
timestamp 0
transform -1 0 5470 0 1 11290
box -6 -8 86 248
use OAI22X1  _11416_
timestamp 0
transform -1 0 5630 0 1 11290
box -6 -8 126 248
use NOR2X1  _11417_
timestamp 0
transform -1 0 6770 0 -1 11770
box -6 -8 86 248
use NAND2X1  _11418_
timestamp 0
transform 1 0 5350 0 -1 11770
box -6 -8 86 248
use INVX1  _11419_
timestamp 0
transform -1 0 6350 0 -1 11770
box -6 -8 66 248
use INVX1  _11420_
timestamp 0
transform 1 0 5230 0 -1 12730
box -6 -8 66 248
use NOR2X1  _11421_
timestamp 0
transform -1 0 3690 0 -1 13210
box -6 -8 86 248
use OAI21X1  _11422_
timestamp 0
transform -1 0 3850 0 -1 13210
box -6 -8 106 248
use OAI21X1  _11423_
timestamp 0
transform 1 0 3430 0 -1 12250
box -6 -8 106 248
use OAI21X1  _11424_
timestamp 0
transform 1 0 3630 0 1 12250
box -6 -8 106 248
use NOR2X1  _11425_
timestamp 0
transform 1 0 6690 0 -1 12250
box -6 -8 86 248
use NAND2X1  _11426_
timestamp 0
transform -1 0 6630 0 -1 12250
box -6 -8 86 248
use INVX1  _11427_
timestamp 0
transform 1 0 7210 0 1 11770
box -6 -8 66 248
use NOR2X1  _11428_
timestamp 0
transform 1 0 7070 0 1 11770
box -6 -8 86 248
use OAI21X1  _11429_
timestamp 0
transform -1 0 6490 0 -1 11770
box -6 -8 106 248
use AOI21X1  _11430_
timestamp 0
transform 1 0 6550 0 -1 11770
box -6 -8 106 248
use NOR2X1  _11431_
timestamp 0
transform 1 0 6810 0 -1 11770
box -6 -8 86 248
use NAND2X1  _11432_
timestamp 0
transform 1 0 6150 0 1 11770
box -6 -8 86 248
use INVX1  _11433_
timestamp 0
transform 1 0 6530 0 1 10810
box -6 -8 66 248
use AOI21X1  _11434_
timestamp 0
transform 1 0 3850 0 1 11290
box -6 -8 106 248
use OAI21X1  _11435_
timestamp 0
transform 1 0 3990 0 1 11290
box -6 -8 106 248
use OAI21X1  _11436_
timestamp 0
transform -1 0 4590 0 -1 11290
box -6 -8 106 248
use OR2X2  _11437_
timestamp 0
transform 1 0 6730 0 -1 11290
box -6 -8 106 248
use NAND2X1  _11438_
timestamp 0
transform -1 0 6570 0 -1 11290
box -6 -8 86 248
use NAND2X1  _11439_
timestamp 0
transform 1 0 6890 0 -1 11290
box -6 -8 86 248
use AOI21X1  _11440_
timestamp 0
transform 1 0 6930 0 1 11770
box -6 -8 106 248
use AND2X2  _11441_
timestamp 0
transform -1 0 6250 0 -1 11770
box -6 -8 106 248
use OAI21X1  _11442_
timestamp 0
transform -1 0 6090 0 -1 11770
box -6 -8 106 248
use OAI21X1  _11443_
timestamp 0
transform -1 0 5950 0 -1 11770
box -6 -8 106 248
use OAI21X1  _11444_
timestamp 0
transform 1 0 7030 0 -1 11290
box -6 -8 106 248
use INVX1  _11445_
timestamp 0
transform 1 0 6150 0 1 10810
box -6 -8 66 248
use OAI21X1  _11446_
timestamp 0
transform -1 0 4050 0 -1 14170
box -6 -8 106 248
use OAI21X1  _11447_
timestamp 0
transform -1 0 4030 0 1 13210
box -6 -8 106 248
use OR2X2  _11448_
timestamp 0
transform 1 0 4030 0 -1 13210
box -6 -8 106 248
use NAND2X1  _11449_
timestamp 0
transform 1 0 4190 0 -1 13210
box -6 -8 86 248
use OR2X2  _11450_
timestamp 0
transform 1 0 6390 0 1 10810
box -6 -8 106 248
use NAND2X1  _11451_
timestamp 0
transform -1 0 6350 0 1 10810
box -6 -8 86 248
use NAND2X1  _11452_
timestamp 0
transform 1 0 6630 0 1 10810
box -6 -8 86 248
use INVX1  _11453_
timestamp 0
transform 1 0 6930 0 1 10810
box -6 -8 66 248
use NOR2X1  _11454_
timestamp 0
transform 1 0 7330 0 -1 11290
box -6 -8 86 248
use NAND2X1  _11455_
timestamp 0
transform 1 0 7290 0 1 10810
box -6 -8 86 248
use NAND2X1  _11456_
timestamp 0
transform -1 0 7510 0 1 10810
box -6 -8 86 248
use OAI22X1  _11457_
timestamp 0
transform 1 0 7170 0 -1 11290
box -6 -8 126 248
use NAND2X1  _11458_
timestamp 0
transform -1 0 6510 0 -1 12250
box -6 -8 86 248
use INVX1  _11459_
timestamp 0
transform -1 0 6430 0 1 11290
box -6 -8 66 248
use NAND2X1  _11460_
timestamp 0
transform -1 0 6550 0 1 11290
box -6 -8 86 248
use OAI21X1  _11461_
timestamp 0
transform -1 0 6870 0 1 10810
box -6 -8 106 248
use INVX1  _11462_
timestamp 0
transform -1 0 6670 0 -1 11290
box -6 -8 66 248
use OAI21X1  _11463_
timestamp 0
transform 1 0 6610 0 1 11290
box -6 -8 106 248
use OAI21X1  _11464_
timestamp 0
transform 1 0 3890 0 -1 13210
box -6 -8 106 248
use NOR2X1  _11465_
timestamp 0
transform -1 0 4410 0 -1 13210
box -6 -8 86 248
use NAND2X1  _11466_
timestamp 0
transform -1 0 4670 0 -1 13210
box -6 -8 86 248
use OAI21X1  _11467_
timestamp 0
transform 1 0 4450 0 -1 13210
box -6 -8 106 248
use NAND2X1  _11468_
timestamp 0
transform 1 0 4730 0 -1 13210
box -6 -8 86 248
use NAND2X1  _11469_
timestamp 0
transform -1 0 5290 0 1 12730
box -6 -8 86 248
use OR2X2  _11470_
timestamp 0
transform 1 0 5350 0 1 12730
box -6 -8 106 248
use NAND2X1  _11471_
timestamp 0
transform -1 0 5570 0 1 12730
box -6 -8 86 248
use INVX1  _11472_
timestamp 0
transform 1 0 6110 0 1 12250
box -6 -8 66 248
use NOR2X1  _11473_
timestamp 0
transform 1 0 7070 0 -1 12250
box -6 -8 86 248
use NAND2X1  _11474_
timestamp 0
transform 1 0 6950 0 -1 12250
box -6 -8 86 248
use NAND2X1  _11475_
timestamp 0
transform 1 0 6810 0 1 11770
box -6 -8 86 248
use OAI21X1  _11476_
timestamp 0
transform -1 0 6910 0 -1 12250
box -6 -8 106 248
use INVX1  _11477_
timestamp 0
transform 1 0 5730 0 1 13210
box -6 -8 66 248
use NAND2X1  _11478_
timestamp 0
transform 1 0 6090 0 1 12730
box -6 -8 86 248
use INVX1  _11479_
timestamp 0
transform 1 0 5330 0 -1 12730
box -6 -8 66 248
use NAND2X1  _11480_
timestamp 0
transform -1 0 3510 0 -1 12730
box -6 -8 86 248
use OR2X2  _11481_
timestamp 0
transform 1 0 3550 0 -1 12730
box -6 -8 106 248
use NAND2X1  _11482_
timestamp 0
transform 1 0 3710 0 -1 12730
box -6 -8 86 248
use NOR2X1  _11483_
timestamp 0
transform 1 0 5670 0 -1 12730
box -6 -8 86 248
use INVX1  _11484_
timestamp 0
transform 1 0 5810 0 -1 12730
box -6 -8 66 248
use NAND2X1  _11485_
timestamp 0
transform -1 0 5630 0 -1 12730
box -6 -8 86 248
use NAND2X1  _11486_
timestamp 0
transform 1 0 5910 0 -1 12730
box -6 -8 86 248
use OR2X2  _11487_
timestamp 0
transform 1 0 6170 0 1 13210
box -6 -8 106 248
use AOI21X1  _11488_
timestamp 0
transform -1 0 6110 0 1 13210
box -6 -8 106 248
use AOI22X1  _11489_
timestamp 0
transform 1 0 5850 0 1 13210
box -6 -8 126 248
use NAND2X1  _11490_
timestamp 0
transform -1 0 5550 0 1 12250
box -6 -8 86 248
use NOR2X1  _11491_
timestamp 0
transform -1 0 2630 0 1 12250
box -6 -8 86 248
use INVX1  _11492_
timestamp 0
transform 1 0 2690 0 1 12250
box -6 -8 66 248
use NAND3X1  _11493_
timestamp 0
transform 1 0 3090 0 1 12250
box -6 -8 106 248
use INVX1  _11494_
timestamp 0
transform -1 0 3590 0 1 12250
box -6 -8 66 248
use AOI21X1  _11495_
timestamp 0
transform 1 0 3230 0 1 12250
box -6 -8 106 248
use NOR2X1  _11496_
timestamp 0
transform 1 0 3390 0 1 12250
box -6 -8 86 248
use OAI21X1  _11497_
timestamp 0
transform -1 0 6130 0 -1 12730
box -6 -8 106 248
use NOR2X1  _11498_
timestamp 0
transform -1 0 6050 0 1 12250
box -6 -8 86 248
use AOI21X1  _11499_
timestamp 0
transform -1 0 6190 0 1 11290
box -6 -8 106 248
use NAND3X1  _11500_
timestamp 0
transform -1 0 6330 0 1 11290
box -6 -8 106 248
use OAI21X1  _11501_
timestamp 0
transform -1 0 6030 0 1 11290
box -6 -8 106 248
use NOR2X1  _11502_
timestamp 0
transform 1 0 5090 0 1 12250
box -6 -8 86 248
use NAND2X1  _11503_
timestamp 0
transform -1 0 5050 0 1 12250
box -6 -8 86 248
use NAND2X1  _11504_
timestamp 0
transform -1 0 5290 0 1 12250
box -6 -8 86 248
use OAI21X1  _11505_
timestamp 0
transform 1 0 5330 0 1 12250
box -6 -8 106 248
use AOI21X1  _11506_
timestamp 0
transform -1 0 4450 0 1 12250
box -6 -8 106 248
use OR2X2  _11507_
timestamp 0
transform -1 0 3870 0 1 12250
box -6 -8 106 248
use NAND2X1  _11508_
timestamp 0
transform -1 0 3930 0 -1 12730
box -6 -8 86 248
use NAND2X1  _11509_
timestamp 0
transform -1 0 3990 0 1 12250
box -6 -8 86 248
use AND2X2  _11510_
timestamp 0
transform 1 0 4490 0 1 12250
box -6 -8 106 248
use OAI21X1  _11511_
timestamp 0
transform 1 0 4650 0 1 12250
box -6 -8 106 248
use OAI22X1  _11512_
timestamp 0
transform -1 0 4910 0 1 12250
box -6 -8 126 248
use NAND2X1  _11513_
timestamp 0
transform 1 0 5210 0 -1 11770
box -6 -8 86 248
use OAI21X1  _11514_
timestamp 0
transform 1 0 4030 0 1 12250
box -6 -8 106 248
use NAND3X1  _11515_
timestamp 0
transform 1 0 4190 0 1 12250
box -6 -8 106 248
use INVX1  _11516_
timestamp 0
transform 1 0 4510 0 -1 12250
box -6 -8 66 248
use AOI21X1  _11517_
timestamp 0
transform 1 0 4610 0 -1 12250
box -6 -8 106 248
use INVX1  _11518_
timestamp 0
transform 1 0 3330 0 -1 11770
box -6 -8 66 248
use NAND2X1  _11519_
timestamp 0
transform -1 0 3510 0 -1 11770
box -6 -8 86 248
use NAND2X1  _11520_
timestamp 0
transform -1 0 3650 0 -1 11770
box -6 -8 86 248
use NAND2X1  _11521_
timestamp 0
transform 1 0 3690 0 -1 11770
box -6 -8 86 248
use AND2X2  _11522_
timestamp 0
transform -1 0 4630 0 -1 11770
box -6 -8 106 248
use OAI21X1  _11523_
timestamp 0
transform 1 0 4670 0 -1 11770
box -6 -8 106 248
use OAI21X1  _11524_
timestamp 0
transform 1 0 4810 0 -1 11770
box -6 -8 106 248
use NAND2X1  _11525_
timestamp 0
transform 1 0 5310 0 1 11770
box -6 -8 86 248
use OAI21X1  _11526_
timestamp 0
transform -1 0 4730 0 1 11770
box -6 -8 106 248
use OAI21X1  _11527_
timestamp 0
transform 1 0 5150 0 1 11770
box -6 -8 106 248
use NAND2X1  _11528_
timestamp 0
transform -1 0 4150 0 1 13210
box -6 -8 86 248
use NAND2X1  _11529_
timestamp 0
transform 1 0 2710 0 1 12730
box -6 -8 86 248
use NOR2X1  _11530_
timestamp 0
transform -1 0 3890 0 1 13210
box -6 -8 86 248
use NAND2X1  _11531_
timestamp 0
transform 1 0 2130 0 -1 13690
box -6 -8 86 248
use OAI21X1  _11532_
timestamp 0
transform 1 0 2090 0 -1 14170
box -6 -8 106 248
use NAND2X1  _11533_
timestamp 0
transform 1 0 2830 0 -1 15130
box -6 -8 86 248
use OAI21X1  _11534_
timestamp 0
transform 1 0 2750 0 -1 15610
box -6 -8 106 248
use INVX1  _11535_
timestamp 0
transform -1 0 2150 0 1 12730
box -6 -8 66 248
use OR2X2  _11536_
timestamp 0
transform -1 0 3550 0 1 12730
box -6 -8 106 248
use OAI21X1  _11537_
timestamp 0
transform -1 0 2610 0 -1 13210
box -6 -8 106 248
use OAI21X1  _11538_
timestamp 0
transform -1 0 2750 0 -1 13210
box -6 -8 106 248
use INVX1  _11539_
timestamp 0
transform -1 0 2850 0 -1 13690
box -6 -8 66 248
use OAI21X1  _11540_
timestamp 0
transform -1 0 2590 0 -1 13690
box -6 -8 106 248
use OAI21X1  _11541_
timestamp 0
transform -1 0 2730 0 -1 13690
box -6 -8 106 248
use NAND2X1  _11542_
timestamp 0
transform -1 0 3410 0 1 12730
box -6 -8 86 248
use NAND2X1  _11543_
timestamp 0
transform -1 0 2270 0 1 12730
box -6 -8 86 248
use OAI21X1  _11544_
timestamp 0
transform -1 0 2430 0 1 12730
box -6 -8 106 248
use NAND2X1  _11545_
timestamp 0
transform -1 0 2410 0 1 13690
box -6 -8 86 248
use OAI21X1  _11546_
timestamp 0
transform -1 0 2570 0 1 13690
box -6 -8 106 248
use AND2X2  _11547_
timestamp 0
transform 1 0 2010 0 1 12250
box -6 -8 106 248
use NAND2X1  _11548_
timestamp 0
transform 1 0 2210 0 1 13690
box -6 -8 86 248
use OAI21X1  _11549_
timestamp 0
transform 1 0 2070 0 1 13690
box -6 -8 106 248
use NAND2X1  _11550_
timestamp 0
transform 1 0 2910 0 1 14170
box -6 -8 86 248
use OAI21X1  _11551_
timestamp 0
transform 1 0 2770 0 1 14170
box -6 -8 106 248
use OAI21X1  _11552_
timestamp 0
transform -1 0 3530 0 1 13210
box -6 -8 106 248
use OAI21X1  _11553_
timestamp 0
transform 1 0 3290 0 1 13210
box -6 -8 106 248
use OAI21X1  _11554_
timestamp 0
transform -1 0 3330 0 1 13690
box -6 -8 106 248
use OAI21X1  _11555_
timestamp 0
transform 1 0 3090 0 1 13690
box -6 -8 106 248
use NAND2X1  _11556_
timestamp 0
transform 1 0 2670 0 1 13210
box -6 -8 86 248
use OAI21X1  _11557_
timestamp 0
transform -1 0 2610 0 1 13210
box -6 -8 106 248
use NAND2X1  _11558_
timestamp 0
transform 1 0 2990 0 -1 14650
box -6 -8 86 248
use OAI21X1  _11559_
timestamp 0
transform 1 0 2830 0 -1 14650
box -6 -8 106 248
use NAND2X1  _11560_
timestamp 0
transform -1 0 4210 0 -1 15130
box -6 -8 86 248
use OAI21X1  _11561_
timestamp 0
transform 1 0 3990 0 -1 15130
box -6 -8 106 248
use NAND2X1  _11562_
timestamp 0
transform -1 0 3270 0 -1 15130
box -6 -8 86 248
use OAI21X1  _11563_
timestamp 0
transform 1 0 3150 0 -1 15610
box -6 -8 106 248
use INVX1  _11564_
timestamp 0
transform -1 0 4330 0 -1 13690
box -6 -8 66 248
use OAI21X1  _11565_
timestamp 0
transform 1 0 3750 0 -1 13690
box -6 -8 106 248
use OAI21X1  _11566_
timestamp 0
transform -1 0 4230 0 -1 13690
box -6 -8 106 248
use INVX1  _11567_
timestamp 0
transform 1 0 3570 0 1 13210
box -6 -8 66 248
use OAI21X1  _11568_
timestamp 0
transform -1 0 3410 0 -1 13690
box -6 -8 106 248
use OAI21X1  _11569_
timestamp 0
transform -1 0 3550 0 -1 13690
box -6 -8 106 248
use NAND2X1  _11570_
timestamp 0
transform 1 0 4230 0 -1 14170
box -6 -8 86 248
use OAI21X1  _11571_
timestamp 0
transform 1 0 4350 0 -1 14170
box -6 -8 106 248
use NAND2X1  _11572_
timestamp 0
transform 1 0 3330 0 -1 13210
box -6 -8 86 248
use OAI21X1  _11573_
timestamp 0
transform -1 0 3570 0 -1 13210
box -6 -8 106 248
use NAND2X1  _11574_
timestamp 0
transform 1 0 5030 0 -1 15130
box -6 -8 86 248
use OAI21X1  _11575_
timestamp 0
transform 1 0 4890 0 -1 15130
box -6 -8 106 248
use NAND2X1  _11576_
timestamp 0
transform 1 0 4410 0 -1 15130
box -6 -8 86 248
use OAI21X1  _11577_
timestamp 0
transform 1 0 4270 0 -1 15130
box -6 -8 106 248
use OAI21X1  _11578_
timestamp 0
transform -1 0 4390 0 1 13690
box -6 -8 106 248
use OAI21X1  _11579_
timestamp 0
transform -1 0 4250 0 1 13690
box -6 -8 106 248
use OAI21X1  _11580_
timestamp 0
transform 1 0 3390 0 1 13690
box -6 -8 106 248
use OAI21X1  _11581_
timestamp 0
transform -1 0 3630 0 1 13690
box -6 -8 106 248
use NAND2X1  _11582_
timestamp 0
transform 1 0 5150 0 -1 14170
box -6 -8 86 248
use OAI21X1  _11583_
timestamp 0
transform 1 0 4990 0 -1 14170
box -6 -8 106 248
use NAND2X1  _11584_
timestamp 0
transform -1 0 3750 0 -1 14170
box -6 -8 86 248
use OAI21X1  _11585_
timestamp 0
transform 1 0 3790 0 -1 14170
box -6 -8 106 248
use NAND2X1  _11586_
timestamp 0
transform -1 0 3690 0 1 11770
box -6 -8 86 248
use OAI21X1  _11587_
timestamp 0
transform 1 0 3350 0 1 11770
box -6 -8 106 248
use NAND2X1  _11588_
timestamp 0
transform -1 0 3370 0 -1 12730
box -6 -8 86 248
use OAI21X1  _11589_
timestamp 0
transform -1 0 3250 0 -1 12730
box -6 -8 106 248
use INVX1  _11590_
timestamp 0
transform 1 0 6270 0 1 11770
box -6 -8 66 248
use OAI21X1  _11591_
timestamp 0
transform 1 0 2950 0 1 12250
box -6 -8 106 248
use OAI21X1  _11592_
timestamp 0
transform -1 0 3930 0 -1 12250
box -6 -8 106 248
use INVX1  _11593_
timestamp 0
transform 1 0 4210 0 -1 12730
box -6 -8 66 248
use OAI21X1  _11594_
timestamp 0
transform 1 0 3890 0 1 12730
box -6 -8 106 248
use OAI21X1  _11595_
timestamp 0
transform -1 0 4130 0 1 12730
box -6 -8 106 248
use NAND2X1  _11596_
timestamp 0
transform -1 0 4930 0 1 12730
box -6 -8 86 248
use OAI21X1  _11597_
timestamp 0
transform 1 0 4690 0 1 12730
box -6 -8 106 248
use NAND2X1  _11598_
timestamp 0
transform 1 0 4570 0 1 12730
box -6 -8 86 248
use OAI21X1  _11599_
timestamp 0
transform 1 0 4430 0 1 12730
box -6 -8 106 248
use NAND2X1  _11600_
timestamp 0
transform -1 0 6910 0 -1 10810
box -6 -8 86 248
use OAI21X1  _11601_
timestamp 0
transform 1 0 6690 0 -1 10810
box -6 -8 106 248
use NAND2X1  _11602_
timestamp 0
transform -1 0 5970 0 1 10810
box -6 -8 86 248
use OAI21X1  _11603_
timestamp 0
transform -1 0 6110 0 1 10810
box -6 -8 106 248
use OAI21X1  _11604_
timestamp 0
transform 1 0 3990 0 -1 12250
box -6 -8 106 248
use OAI21X1  _11605_
timestamp 0
transform -1 0 4230 0 -1 12250
box -6 -8 106 248
use OAI21X1  _11606_
timestamp 0
transform 1 0 4830 0 -1 12730
box -6 -8 106 248
use OAI21X1  _11607_
timestamp 0
transform 1 0 4670 0 -1 12730
box -6 -8 106 248
use NAND2X1  _11608_
timestamp 0
transform -1 0 3830 0 1 11770
box -6 -8 86 248
use OAI21X1  _11609_
timestamp 0
transform -1 0 3970 0 1 11770
box -6 -8 106 248
use NAND2X1  _11610_
timestamp 0
transform -1 0 4210 0 1 11290
box -6 -8 86 248
use OAI21X1  _11611_
timestamp 0
transform -1 0 4370 0 1 11290
box -6 -8 106 248
use DFFPOSX1  _11612_
timestamp 0
transform 1 0 4630 0 1 13690
box -6 -8 246 248
use DFFPOSX1  _11613_
timestamp 0
transform 1 0 4830 0 -1 13690
box -6 -8 246 248
use DFFPOSX1  _11614_
timestamp 0
transform 1 0 8070 0 1 11290
box -6 -8 246 248
use DFFPOSX1  _11615_
timestamp 0
transform -1 0 5470 0 -1 14170
box -6 -8 246 248
use DFFPOSX1  _11616_
timestamp 0
transform -1 0 5350 0 -1 15130
box -6 -8 246 248
use DFFPOSX1  _11617_
timestamp 0
transform 1 0 5570 0 -1 14650
box -6 -8 246 248
use DFFPOSX1  _11618_
timestamp 0
transform -1 0 5790 0 -1 16090
box -6 -8 246 248
use DFFPOSX1  _11619_
timestamp 0
transform -1 0 6410 0 1 14650
box -6 -8 246 248
use DFFPOSX1  _11620_
timestamp 0
transform 1 0 5470 0 1 15610
box -6 -8 246 248
use DFFPOSX1  _11621_
timestamp 0
transform 1 0 5510 0 -1 15130
box -6 -8 246 248
use DFFPOSX1  _11622_
timestamp 0
transform -1 0 5930 0 -1 15610
box -6 -8 246 248
use DFFPOSX1  _11623_
timestamp 0
transform -1 0 6210 0 1 14170
box -6 -8 246 248
use DFFPOSX1  _11624_
timestamp 0
transform 1 0 5330 0 -1 14650
box -6 -8 246 248
use DFFPOSX1  _11625_
timestamp 0
transform 1 0 1730 0 -1 13690
box -6 -8 246 248
use DFFPOSX1  _11626_
timestamp 0
transform -1 0 3050 0 1 11770
box -6 -8 246 248
use DFFPOSX1  _11627_
timestamp 0
transform 1 0 1970 0 -1 13210
box -6 -8 246 248
use DFFPOSX1  _11628_
timestamp 0
transform 1 0 2470 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _11629_
timestamp 0
transform 1 0 1290 0 1 12730
box -6 -8 246 248
use DFFPOSX1  _11630_
timestamp 0
transform 1 0 10 0 -1 12250
box -6 -8 246 248
use DFFPOSX1  _11631_
timestamp 0
transform -1 0 1810 0 -1 12250
box -6 -8 246 248
use DFFPOSX1  _11632_
timestamp 0
transform 1 0 950 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _11633_
timestamp 0
transform 1 0 830 0 -1 12250
box -6 -8 246 248
use DFFPOSX1  _11634_
timestamp 0
transform 1 0 270 0 1 12250
box -6 -8 246 248
use DFFPOSX1  _11635_
timestamp 0
transform 1 0 1810 0 1 12730
box -6 -8 246 248
use DFFPOSX1  _11636_
timestamp 0
transform 1 0 970 0 1 12250
box -6 -8 246 248
use DFFPOSX1  _11637_
timestamp 0
transform 1 0 5530 0 1 11770
box -6 -8 246 248
use DFFPOSX1  _11638_
timestamp 0
transform 1 0 6210 0 -1 11290
box -6 -8 246 248
use DFFPOSX1  _11639_
timestamp 0
transform 1 0 5550 0 -1 11290
box -6 -8 246 248
use DFFPOSX1  _11640_
timestamp 0
transform -1 0 7130 0 -1 11770
box -6 -8 246 248
use DFFPOSX1  _11641_
timestamp 0
transform 1 0 5570 0 -1 11770
box -6 -8 246 248
use DFFPOSX1  _11642_
timestamp 0
transform -1 0 7070 0 1 11290
box -6 -8 246 248
use DFFPOSX1  _11643_
timestamp 0
transform -1 0 6670 0 1 12250
box -6 -8 246 248
use DFFPOSX1  _11644_
timestamp 0
transform -1 0 5930 0 -1 13210
box -6 -8 246 248
use DFFPOSX1  _11645_
timestamp 0
transform -1 0 5930 0 1 12250
box -6 -8 246 248
use DFFPOSX1  _11646_
timestamp 0
transform 1 0 4850 0 -1 12250
box -6 -8 246 248
use DFFPOSX1  _11647_
timestamp 0
transform 1 0 4910 0 -1 11770
box -6 -8 246 248
use DFFPOSX1  _11648_
timestamp 0
transform 1 0 4850 0 1 11770
box -6 -8 246 248
use DFFPOSX1  _11649_
timestamp 0
transform -1 0 2430 0 -1 14170
box -6 -8 246 248
use DFFPOSX1  _11650_
timestamp 0
transform -1 0 2410 0 1 15610
box -6 -8 246 248
use DFFPOSX1  _11651_
timestamp 0
transform -1 0 2450 0 -1 13210
box -6 -8 246 248
use DFFPOSX1  _11652_
timestamp 0
transform -1 0 2450 0 -1 13690
box -6 -8 246 248
use DFFPOSX1  _11653_
timestamp 0
transform -1 0 2670 0 1 12730
box -6 -8 246 248
use DFFPOSX1  _11654_
timestamp 0
transform 1 0 2570 0 1 13690
box -6 -8 246 248
use DFFPOSX1  _11655_
timestamp 0
transform -1 0 2010 0 1 13690
box -6 -8 246 248
use DFFPOSX1  _11656_
timestamp 0
transform -1 0 2710 0 1 14170
box -6 -8 246 248
use DFFPOSX1  _11657_
timestamp 0
transform -1 0 3230 0 1 13210
box -6 -8 246 248
use DFFPOSX1  _11658_
timestamp 0
transform -1 0 3050 0 1 13690
box -6 -8 246 248
use DFFPOSX1  _11659_
timestamp 0
transform -1 0 2470 0 1 13210
box -6 -8 246 248
use DFFPOSX1  _11660_
timestamp 0
transform 1 0 2750 0 1 14650
box -6 -8 246 248
use DFFPOSX1  _11661_
timestamp 0
transform -1 0 4090 0 1 15130
box -6 -8 246 248
use DFFPOSX1  _11662_
timestamp 0
transform -1 0 3090 0 -1 15610
box -6 -8 246 248
use DFFPOSX1  _11663_
timestamp 0
transform -1 0 4090 0 -1 13690
box -6 -8 246 248
use DFFPOSX1  _11664_
timestamp 0
transform 1 0 3010 0 -1 13690
box -6 -8 246 248
use DFFPOSX1  _11665_
timestamp 0
transform -1 0 4690 0 -1 14170
box -6 -8 246 248
use DFFPOSX1  _11666_
timestamp 0
transform -1 0 3290 0 -1 13210
box -6 -8 246 248
use DFFPOSX1  _11667_
timestamp 0
transform -1 0 4830 0 -1 15130
box -6 -8 246 248
use DFFPOSX1  _11668_
timestamp 0
transform -1 0 4430 0 1 15130
box -6 -8 246 248
use DFFPOSX1  _11669_
timestamp 0
transform -1 0 4110 0 1 13690
box -6 -8 246 248
use DFFPOSX1  _11670_
timestamp 0
transform -1 0 3870 0 1 13690
box -6 -8 246 248
use DFFPOSX1  _11671_
timestamp 0
transform -1 0 5310 0 1 14170
box -6 -8 246 248
use DFFPOSX1  _11672_
timestamp 0
transform 1 0 3990 0 1 14170
box -6 -8 246 248
use DFFPOSX1  _11673_
timestamp 0
transform 1 0 3030 0 -1 11770
box -6 -8 246 248
use DFFPOSX1  _11674_
timestamp 0
transform -1 0 3270 0 1 12730
box -6 -8 246 248
use DFFPOSX1  _11675_
timestamp 0
transform -1 0 3770 0 -1 12250
box -6 -8 246 248
use DFFPOSX1  _11676_
timestamp 0
transform -1 0 4170 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _11677_
timestamp 0
transform 1 0 4930 0 1 12730
box -6 -8 246 248
use DFFPOSX1  _11678_
timestamp 0
transform 1 0 4130 0 1 12730
box -6 -8 246 248
use DFFPOSX1  _11679_
timestamp 0
transform -1 0 6630 0 -1 10810
box -6 -8 246 248
use DFFPOSX1  _11680_
timestamp 0
transform 1 0 5910 0 -1 10810
box -6 -8 246 248
use DFFPOSX1  _11681_
timestamp 0
transform -1 0 4470 0 -1 12250
box -6 -8 246 248
use DFFPOSX1  _11682_
timestamp 0
transform 1 0 4930 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _11683_
timestamp 0
transform 1 0 3970 0 1 11770
box -6 -8 246 248
use DFFPOSX1  _11684_
timestamp 0
transform -1 0 5610 0 1 10810
box -6 -8 246 248
use DFFPOSX1  _11685_
timestamp 0
transform -1 0 7310 0 1 11290
box -6 -8 246 248
use DFFPOSX1  _11686_
timestamp 0
transform 1 0 4270 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _11687_
timestamp 0
transform 1 0 4930 0 -1 13210
box -6 -8 246 248
use DFFPOSX1  _11688_
timestamp 0
transform 1 0 5050 0 1 13210
box -6 -8 246 248
use DFFPOSX1  _11689_
timestamp 0
transform -1 0 5410 0 -1 13210
box -6 -8 246 248
use DFFPOSX1  _11690_
timestamp 0
transform -1 0 4630 0 1 13210
box -6 -8 246 248
use DFFPOSX1  _11691_
timestamp 0
transform -1 0 4390 0 1 13210
box -6 -8 246 248
use INVX1  _11692_
timestamp 0
transform 1 0 9910 0 -1 8890
box -6 -8 66 248
use INVX2  _11693_
timestamp 0
transform 1 0 11370 0 -1 8410
box -6 -8 66 248
use NOR2X1  _11694_
timestamp 0
transform -1 0 12710 0 1 9850
box -6 -8 86 248
use INVX2  _11695_
timestamp 0
transform 1 0 13310 0 -1 9370
box -6 -8 66 248
use NOR2X1  _11696_
timestamp 0
transform 1 0 11530 0 1 10810
box -6 -8 86 248
use INVX4  _11697_
timestamp 0
transform -1 0 11510 0 -1 7930
box -6 -8 86 248
use NOR2X1  _11698_
timestamp 0
transform -1 0 11870 0 -1 11290
box -6 -8 86 248
use OAI21X1  _11699_
timestamp 0
transform -1 0 11190 0 1 10810
box -6 -8 106 248
use INVX2  _11700_
timestamp 0
transform -1 0 11930 0 -1 8890
box -6 -8 66 248
use AND2X2  _11701_
timestamp 0
transform -1 0 11690 0 1 11290
box -6 -8 106 248
use AOI22X1  _11702_
timestamp 0
transform -1 0 10930 0 1 11290
box -6 -8 126 248
use OAI21X1  _11703_
timestamp 0
transform -1 0 11050 0 1 10810
box -6 -8 106 248
use NOR2X1  _11704_
timestamp 0
transform -1 0 11310 0 -1 8410
box -6 -8 86 248
use AOI22X1  _11705_
timestamp 0
transform -1 0 12030 0 -1 10330
box -6 -8 126 248
use OAI21X1  _11706_
timestamp 0
transform 1 0 12070 0 -1 10330
box -6 -8 106 248
use INVX1  _11707_
timestamp 0
transform 1 0 11530 0 -1 11290
box -6 -8 66 248
use OAI21X1  _11708_
timestamp 0
transform -1 0 12010 0 -1 11290
box -6 -8 106 248
use AOI21X1  _11709_
timestamp 0
transform -1 0 11730 0 -1 11290
box -6 -8 106 248
use INVX1  _11710_
timestamp 0
transform 1 0 9650 0 -1 11290
box -6 -8 66 248
use NAND2X1  _11711_
timestamp 0
transform 1 0 10810 0 -1 11290
box -6 -8 86 248
use OAI21X1  _11712_
timestamp 0
transform -1 0 11050 0 -1 11290
box -6 -8 106 248
use OAI21X1  _11713_
timestamp 0
transform 1 0 11090 0 -1 11290
box -6 -8 106 248
use AOI22X1  _11714_
timestamp 0
transform 1 0 11450 0 -1 10330
box -6 -8 126 248
use NAND2X1  _11715_
timestamp 0
transform 1 0 11230 0 -1 11290
box -6 -8 86 248
use INVX1  _11716_
timestamp 0
transform -1 0 13850 0 1 7450
box -6 -8 66 248
use OAI21X1  _11717_
timestamp 0
transform -1 0 13610 0 1 7450
box -6 -8 106 248
use AOI21X1  _11718_
timestamp 0
transform -1 0 13750 0 1 7450
box -6 -8 106 248
use INVX1  _11719_
timestamp 0
transform -1 0 13630 0 -1 6970
box -6 -8 66 248
use NAND2X1  _11720_
timestamp 0
transform -1 0 13210 0 -1 7450
box -6 -8 86 248
use OAI21X1  _11721_
timestamp 0
transform 1 0 12990 0 -1 7450
box -6 -8 106 248
use OAI21X1  _11722_
timestamp 0
transform -1 0 13050 0 1 7450
box -6 -8 106 248
use AOI22X1  _11723_
timestamp 0
transform -1 0 12550 0 -1 8410
box -6 -8 126 248
use NAND2X1  _11724_
timestamp 0
transform 1 0 12890 0 -1 8410
box -6 -8 86 248
use INVX1  _11725_
timestamp 0
transform -1 0 13430 0 1 6970
box -6 -8 66 248
use OAI21X1  _11726_
timestamp 0
transform 1 0 13210 0 1 7450
box -6 -8 106 248
use AOI21X1  _11727_
timestamp 0
transform 1 0 13350 0 1 7450
box -6 -8 106 248
use INVX1  _11728_
timestamp 0
transform 1 0 12470 0 -1 7450
box -6 -8 66 248
use NAND2X1  _11729_
timestamp 0
transform 1 0 12870 0 -1 7450
box -6 -8 86 248
use OAI21X1  _11730_
timestamp 0
transform 1 0 12710 0 -1 7450
box -6 -8 106 248
use OAI21X1  _11731_
timestamp 0
transform -1 0 12890 0 1 7450
box -6 -8 106 248
use AOI22X1  _11732_
timestamp 0
transform 1 0 12590 0 -1 8410
box -6 -8 126 248
use NAND2X1  _11733_
timestamp 0
transform 1 0 12750 0 -1 8410
box -6 -8 86 248
use INVX1  _11734_
timestamp 0
transform -1 0 13290 0 1 11290
box -6 -8 66 248
use OAI21X1  _11735_
timestamp 0
transform -1 0 13130 0 -1 11290
box -6 -8 106 248
use AOI21X1  _11736_
timestamp 0
transform -1 0 13170 0 1 11290
box -6 -8 106 248
use INVX1  _11737_
timestamp 0
transform -1 0 13470 0 -1 11770
box -6 -8 66 248
use NAND2X1  _11738_
timestamp 0
transform -1 0 12450 0 1 11290
box -6 -8 86 248
use OAI21X1  _11739_
timestamp 0
transform -1 0 12590 0 1 11290
box -6 -8 106 248
use OAI21X1  _11740_
timestamp 0
transform -1 0 12730 0 1 11290
box -6 -8 106 248
use AOI22X1  _11741_
timestamp 0
transform 1 0 13010 0 -1 10810
box -6 -8 126 248
use NAND2X1  _11742_
timestamp 0
transform -1 0 13010 0 1 11290
box -6 -8 86 248
use INVX1  _11743_
timestamp 0
transform -1 0 14650 0 -1 12250
box -6 -8 66 248
use NOR2X1  _11744_
timestamp 0
transform 1 0 12910 0 -1 11290
box -6 -8 86 248
use OAI21X1  _11745_
timestamp 0
transform -1 0 13090 0 1 10810
box -6 -8 106 248
use AOI22X1  _11746_
timestamp 0
transform 1 0 12770 0 1 11290
box -6 -8 126 248
use OAI21X1  _11747_
timestamp 0
transform -1 0 12870 0 -1 11290
box -6 -8 106 248
use AOI22X1  _11748_
timestamp 0
transform -1 0 12730 0 -1 11290
box -6 -8 126 248
use OAI21X1  _11749_
timestamp 0
transform -1 0 14350 0 1 11770
box -6 -8 106 248
use INVX1  _11750_
timestamp 0
transform 1 0 12510 0 1 7930
box -6 -8 66 248
use INVX1  _11751_
timestamp 0
transform 1 0 12770 0 -1 9370
box -6 -8 66 248
use INVX8  _11752_
timestamp 0
transform 1 0 16230 0 1 8890
box -6 -8 126 248
use INVX8  _11753_
timestamp 0
transform -1 0 16290 0 1 9370
box -6 -8 126 248
use INVX1  _11754_
timestamp 0
transform -1 0 14830 0 -1 11290
box -6 -8 66 248
use NAND2X1  _11755_
timestamp 0
transform 1 0 15030 0 -1 11290
box -6 -8 86 248
use OAI21X1  _11756_
timestamp 0
transform 1 0 14870 0 -1 11290
box -6 -8 106 248
use INVX1  _11757_
timestamp 0
transform -1 0 16390 0 -1 12250
box -6 -8 66 248
use NAND2X1  _11758_
timestamp 0
transform -1 0 15790 0 1 10330
box -6 -8 86 248
use OAI21X1  _11759_
timestamp 0
transform 1 0 15830 0 1 10330
box -6 -8 106 248
use MUX2X1  _11760_
timestamp 0
transform 1 0 14870 0 -1 10330
box -6 -8 126 248
use INVX1  _11761_
timestamp 0
transform 1 0 13230 0 1 9850
box -6 -8 66 248
use NAND2X1  _11762_
timestamp 0
transform 1 0 13350 0 1 9850
box -6 -8 86 248
use OAI21X1  _11763_
timestamp 0
transform 1 0 13090 0 1 9850
box -6 -8 106 248
use INVX1  _11764_
timestamp 0
transform 1 0 13150 0 -1 10330
box -6 -8 66 248
use NAND2X1  _11765_
timestamp 0
transform 1 0 13410 0 -1 10330
box -6 -8 86 248
use OAI21X1  _11766_
timestamp 0
transform 1 0 13250 0 -1 10330
box -6 -8 106 248
use MUX2X1  _11767_
timestamp 0
transform -1 0 13050 0 1 9850
box -6 -8 126 248
use MUX2X1  _11768_
timestamp 0
transform 1 0 12750 0 1 9850
box -6 -8 126 248
use NOR2X1  _11769_
timestamp 0
transform 1 0 13170 0 -1 9370
box -6 -8 86 248
use NAND2X1  _11770_
timestamp 0
transform -1 0 12730 0 1 8890
box -6 -8 86 248
use INVX1  _11771_
timestamp 0
transform 1 0 12910 0 1 8890
box -6 -8 66 248
use NAND2X1  _11772_
timestamp 0
transform 1 0 14910 0 -1 9850
box -6 -8 86 248
use OAI21X1  _11773_
timestamp 0
transform -1 0 12550 0 -1 11290
box -6 -8 106 248
use INVX2  _11774_
timestamp 0
transform -1 0 13370 0 -1 11770
box -6 -8 66 248
use OAI21X1  _11775_
timestamp 0
transform -1 0 13110 0 -1 9370
box -6 -8 106 248
use OAI21X1  _11776_
timestamp 0
transform 1 0 12630 0 1 7930
box -6 -8 106 248
use INVX8  _11777_
timestamp 0
transform -1 0 12290 0 1 10810
box -6 -8 126 248
use NAND2X1  _11778_
timestamp 0
transform -1 0 12510 0 1 8410
box -6 -8 86 248
use NOR2X1  _11779_
timestamp 0
transform -1 0 14050 0 1 10330
box -6 -8 86 248
use MUX2X1  _11780_
timestamp 0
transform -1 0 15350 0 1 9370
box -6 -8 126 248
use MUX2X1  _11781_
timestamp 0
transform 1 0 15330 0 -1 9850
box -6 -8 126 248
use MUX2X1  _11782_
timestamp 0
transform -1 0 15190 0 1 9370
box -6 -8 126 248
use INVX2  _11783_
timestamp 0
transform 1 0 12470 0 1 9370
box -6 -8 66 248
use NAND2X1  _11784_
timestamp 0
transform -1 0 13270 0 -1 9850
box -6 -8 86 248
use AOI21X1  _11785_
timestamp 0
transform 1 0 13310 0 -1 9850
box -6 -8 106 248
use NAND3X1  _11786_
timestamp 0
transform -1 0 12990 0 -1 9850
box -6 -8 106 248
use NAND3X1  _11787_
timestamp 0
transform -1 0 13130 0 -1 9850
box -6 -8 106 248
use NAND3X1  _11788_
timestamp 0
transform 1 0 12870 0 1 9370
box -6 -8 106 248
use OAI22X1  _11789_
timestamp 0
transform -1 0 13270 0 1 9370
box -6 -8 126 248
use INVX1  _11790_
timestamp 0
transform -1 0 12370 0 1 8890
box -6 -8 66 248
use INVX8  _11791_
timestamp 0
transform -1 0 12150 0 -1 8410
box -6 -8 126 248
use INVX1  _11792_
timestamp 0
transform 1 0 15630 0 1 10810
box -6 -8 66 248
use NAND2X1  _11793_
timestamp 0
transform -1 0 15530 0 1 10330
box -6 -8 86 248
use OAI21X1  _11794_
timestamp 0
transform -1 0 15670 0 1 10330
box -6 -8 106 248
use INVX1  _11795_
timestamp 0
transform -1 0 15690 0 1 11770
box -6 -8 66 248
use NAND2X1  _11796_
timestamp 0
transform -1 0 15250 0 -1 11290
box -6 -8 86 248
use OAI21X1  _11797_
timestamp 0
transform 1 0 15290 0 -1 11290
box -6 -8 106 248
use MUX2X1  _11798_
timestamp 0
transform 1 0 15670 0 -1 9850
box -6 -8 126 248
use INVX1  _11799_
timestamp 0
transform -1 0 14870 0 1 9850
box -6 -8 66 248
use NAND2X1  _11800_
timestamp 0
transform 1 0 15390 0 1 9850
box -6 -8 86 248
use OAI21X1  _11801_
timestamp 0
transform -1 0 15610 0 1 9850
box -6 -8 106 248
use INVX1  _11802_
timestamp 0
transform 1 0 13470 0 1 9850
box -6 -8 66 248
use NAND2X1  _11803_
timestamp 0
transform -1 0 15010 0 1 9850
box -6 -8 86 248
use OAI21X1  _11804_
timestamp 0
transform 1 0 15050 0 1 9850
box -6 -8 106 248
use MUX2X1  _11805_
timestamp 0
transform -1 0 15330 0 1 9850
box -6 -8 126 248
use MUX2X1  _11806_
timestamp 0
transform -1 0 15270 0 -1 9850
box -6 -8 126 248
use NAND3X1  _11807_
timestamp 0
transform -1 0 13530 0 -1 9370
box -6 -8 106 248
use MUX2X1  _11808_
timestamp 0
transform 1 0 15390 0 1 9370
box -6 -8 126 248
use MUX2X1  _11809_
timestamp 0
transform -1 0 15610 0 -1 9850
box -6 -8 126 248
use MUX2X1  _11810_
timestamp 0
transform -1 0 15690 0 1 9370
box -6 -8 126 248
use MUX2X1  _11811_
timestamp 0
transform 1 0 14650 0 1 9850
box -6 -8 126 248
use MUX2X1  _11812_
timestamp 0
transform 1 0 13470 0 -1 9850
box -6 -8 126 248
use MUX2X1  _11813_
timestamp 0
transform -1 0 14670 0 -1 9850
box -6 -8 126 248
use MUX2X1  _11814_
timestamp 0
transform -1 0 14750 0 1 9370
box -6 -8 126 248
use OAI21X1  _11815_
timestamp 0
transform 1 0 13310 0 1 8890
box -6 -8 106 248
use AOI21X1  _11816_
timestamp 0
transform -1 0 13110 0 1 8890
box -6 -8 106 248
use INVX1  _11817_
timestamp 0
transform -1 0 12450 0 -1 8890
box -6 -8 66 248
use NAND3X1  _11818_
timestamp 0
transform -1 0 13250 0 1 8890
box -6 -8 106 248
use AND2X2  _11819_
timestamp 0
transform 1 0 12510 0 -1 8890
box -6 -8 106 248
use OAI21X1  _11820_
timestamp 0
transform -1 0 12750 0 -1 8890
box -6 -8 106 248
use OR2X2  _11821_
timestamp 0
transform 1 0 12850 0 1 8410
box -6 -8 106 248
use AOI21X1  _11822_
timestamp 0
transform -1 0 12810 0 1 8410
box -6 -8 106 248
use OAI21X1  _11823_
timestamp 0
transform -1 0 12650 0 1 8410
box -6 -8 106 248
use INVX1  _11824_
timestamp 0
transform 1 0 9390 0 1 11290
box -6 -8 66 248
use NAND2X1  _11825_
timestamp 0
transform -1 0 8810 0 1 11290
box -6 -8 86 248
use OAI21X1  _11826_
timestamp 0
transform -1 0 8970 0 1 11290
box -6 -8 106 248
use NAND2X1  _11827_
timestamp 0
transform 1 0 12510 0 -1 7930
box -6 -8 86 248
use AOI21X1  _11828_
timestamp 0
transform 1 0 12770 0 1 8890
box -6 -8 106 248
use MUX2X1  _11829_
timestamp 0
transform 1 0 15350 0 -1 9370
box -6 -8 126 248
use MUX2X1  _11830_
timestamp 0
transform 1 0 15170 0 -1 9370
box -6 -8 126 248
use MUX2X1  _11831_
timestamp 0
transform 1 0 14730 0 -1 9850
box -6 -8 126 248
use NAND2X1  _11832_
timestamp 0
transform 1 0 14950 0 1 9370
box -6 -8 86 248
use OAI22X1  _11833_
timestamp 0
transform -1 0 14910 0 1 9370
box -6 -8 126 248
use AOI21X1  _11834_
timestamp 0
transform -1 0 14930 0 1 8890
box -6 -8 106 248
use AOI21X1  _11835_
timestamp 0
transform -1 0 13870 0 -1 8890
box -6 -8 106 248
use NAND2X1  _11836_
timestamp 0
transform 1 0 13650 0 -1 8890
box -6 -8 86 248
use INVX1  _11837_
timestamp 0
transform 1 0 13570 0 1 8890
box -6 -8 66 248
use OAI21X1  _11838_
timestamp 0
transform 1 0 13590 0 -1 9370
box -6 -8 106 248
use NAND2X1  _11839_
timestamp 0
transform -1 0 13530 0 1 8890
box -6 -8 86 248
use AOI21X1  _11840_
timestamp 0
transform -1 0 13130 0 -1 8890
box -6 -8 106 248
use NAND3X1  _11841_
timestamp 0
transform 1 0 13190 0 -1 8890
box -6 -8 106 248
use INVX1  _11842_
timestamp 0
transform -1 0 13210 0 1 8410
box -6 -8 66 248
use OR2X2  _11843_
timestamp 0
transform 1 0 13270 0 1 8410
box -6 -8 106 248
use NOR2X1  _11844_
timestamp 0
transform 1 0 13250 0 -1 8410
box -6 -8 86 248
use INVX1  _11845_
timestamp 0
transform -1 0 13210 0 -1 8410
box -6 -8 66 248
use OAI21X1  _11846_
timestamp 0
transform -1 0 13110 0 1 8410
box -6 -8 106 248
use AOI21X1  _11847_
timestamp 0
transform -1 0 13110 0 -1 8410
box -6 -8 106 248
use INVX2  _11848_
timestamp 0
transform 1 0 15390 0 1 6970
box -6 -8 66 248
use OAI21X1  _11849_
timestamp 0
transform -1 0 12890 0 -1 7930
box -6 -8 106 248
use OAI21X1  _11850_
timestamp 0
transform -1 0 12750 0 -1 7930
box -6 -8 106 248
use INVX1  _11851_
timestamp 0
transform 1 0 13090 0 1 7450
box -6 -8 66 248
use INVX2  _11852_
timestamp 0
transform 1 0 12930 0 -1 7930
box -6 -8 66 248
use OAI21X1  _11853_
timestamp 0
transform 1 0 13430 0 1 8410
box -6 -8 106 248
use INVX1  _11854_
timestamp 0
transform -1 0 13470 0 -1 7450
box -6 -8 66 248
use INVX1  _11855_
timestamp 0
transform 1 0 16190 0 1 8410
box -6 -8 66 248
use NAND3X1  _11856_
timestamp 0
transform 1 0 13910 0 -1 8890
box -6 -8 106 248
use INVX1  _11857_
timestamp 0
transform -1 0 14810 0 -1 10330
box -6 -8 66 248
use NAND2X1  _11858_
timestamp 0
transform 1 0 14390 0 1 9850
box -6 -8 86 248
use OAI21X1  _11859_
timestamp 0
transform 1 0 14510 0 1 9850
box -6 -8 106 248
use NAND2X1  _11860_
timestamp 0
transform -1 0 15730 0 -1 9370
box -6 -8 86 248
use OAI21X1  _11861_
timestamp 0
transform 1 0 15650 0 1 8890
box -6 -8 106 248
use NOR2X1  _11862_
timestamp 0
transform 1 0 17050 0 1 9370
box -6 -8 86 248
use NOR2X1  _11863_
timestamp 0
transform 1 0 16450 0 1 9370
box -6 -8 86 248
use AOI22X1  _11864_
timestamp 0
transform 1 0 15990 0 1 9370
box -6 -8 126 248
use OAI21X1  _11865_
timestamp 0
transform 1 0 15950 0 1 8890
box -6 -8 106 248
use NAND3X1  _11866_
timestamp 0
transform 1 0 15790 0 -1 7930
box -6 -8 106 248
use INVX1  _11867_
timestamp 0
transform 1 0 17110 0 1 7930
box -6 -8 66 248
use INVX1  _11868_
timestamp 0
transform 1 0 16710 0 -1 8410
box -6 -8 66 248
use OAI21X1  _11869_
timestamp 0
transform 1 0 16810 0 1 7930
box -6 -8 106 248
use NAND3X1  _11870_
timestamp 0
transform -1 0 15910 0 1 7450
box -6 -8 106 248
use AOI21X1  _11871_
timestamp 0
transform -1 0 15770 0 1 7450
box -6 -8 106 248
use INVX1  _11872_
timestamp 0
transform -1 0 14990 0 -1 7450
box -6 -8 66 248
use NAND2X1  _11873_
timestamp 0
transform 1 0 14790 0 -1 7450
box -6 -8 86 248
use AOI21X1  _11874_
timestamp 0
transform -1 0 13770 0 -1 7450
box -6 -8 106 248
use OAI21X1  _11875_
timestamp 0
transform -1 0 13610 0 -1 7450
box -6 -8 106 248
use AOI22X1  _11876_
timestamp 0
transform 1 0 13250 0 -1 7450
box -6 -8 126 248
use AOI21X1  _11877_
timestamp 0
transform 1 0 15190 0 -1 7450
box -6 -8 106 248
use INVX1  _11878_
timestamp 0
transform -1 0 17130 0 -1 8410
box -6 -8 66 248
use INVX1  _11879_
timestamp 0
transform 1 0 14450 0 -1 9850
box -6 -8 66 248
use NAND2X1  _11880_
timestamp 0
transform 1 0 14690 0 -1 9370
box -6 -8 86 248
use OAI21X1  _11881_
timestamp 0
transform 1 0 14490 0 1 9370
box -6 -8 106 248
use NAND2X1  _11882_
timestamp 0
transform -1 0 15590 0 -1 9370
box -6 -8 86 248
use OAI21X1  _11883_
timestamp 0
transform -1 0 15870 0 -1 9370
box -6 -8 106 248
use NAND2X1  _11884_
timestamp 0
transform -1 0 15890 0 1 8890
box -6 -8 86 248
use OAI21X1  _11885_
timestamp 0
transform -1 0 16190 0 1 8890
box -6 -8 106 248
use INVX2  _11886_
timestamp 0
transform -1 0 16890 0 -1 8410
box -6 -8 66 248
use OAI21X1  _11887_
timestamp 0
transform 1 0 16870 0 -1 7930
box -6 -8 106 248
use OR2X2  _11888_
timestamp 0
transform 1 0 16990 0 -1 7450
box -6 -8 106 248
use NOR2X1  _11889_
timestamp 0
transform 1 0 16750 0 -1 7930
box -6 -8 86 248
use OAI21X1  _11890_
timestamp 0
transform 1 0 16750 0 1 7450
box -6 -8 106 248
use NAND3X1  _11891_
timestamp 0
transform 1 0 16830 0 -1 7450
box -6 -8 106 248
use NOR2X1  _11892_
timestamp 0
transform -1 0 16970 0 1 7450
box -6 -8 86 248
use AND2X2  _11893_
timestamp 0
transform -1 0 17130 0 -1 7930
box -6 -8 106 248
use OAI21X1  _11894_
timestamp 0
transform 1 0 17010 0 1 7450
box -6 -8 106 248
use NAND2X1  _11895_
timestamp 0
transform 1 0 17070 0 -1 6970
box -6 -8 86 248
use AOI21X1  _11896_
timestamp 0
transform -1 0 15590 0 -1 6970
box -6 -8 106 248
use OAI21X1  _11897_
timestamp 0
transform -1 0 15430 0 -1 6970
box -6 -8 106 248
use AOI22X1  _11898_
timestamp 0
transform 1 0 14030 0 -1 6970
box -6 -8 126 248
use OAI21X1  _11899_
timestamp 0
transform 1 0 16330 0 -1 6970
box -6 -8 106 248
use INVX1  _11900_
timestamp 0
transform -1 0 17010 0 -1 8890
box -6 -8 66 248
use NAND3X1  _11901_
timestamp 0
transform 1 0 16950 0 1 7930
box -6 -8 106 248
use NAND2X1  _11902_
timestamp 0
transform -1 0 14770 0 1 8890
box -6 -8 86 248
use INVX1  _11903_
timestamp 0
transform 1 0 14990 0 1 8890
box -6 -8 66 248
use AOI21X1  _11904_
timestamp 0
transform 1 0 15370 0 1 8890
box -6 -8 106 248
use NAND2X1  _11905_
timestamp 0
transform 1 0 15530 0 1 8890
box -6 -8 86 248
use OAI21X1  _11906_
timestamp 0
transform 1 0 15590 0 1 8410
box -6 -8 106 248
use NAND3X1  _11907_
timestamp 0
transform 1 0 16610 0 1 7450
box -6 -8 106 248
use NOR3X1  _11908_
timestamp 0
transform -1 0 16750 0 1 7930
box -6 -8 186 248
use INVX1  _11909_
timestamp 0
transform 1 0 16510 0 -1 7930
box -6 -8 66 248
use OAI21X1  _11910_
timestamp 0
transform -1 0 16470 0 -1 7930
box -6 -8 106 248
use NAND3X1  _11911_
timestamp 0
transform -1 0 16450 0 -1 7450
box -6 -8 106 248
use AOI21X1  _11912_
timestamp 0
transform 1 0 16510 0 -1 7450
box -6 -8 106 248
use INVX1  _11913_
timestamp 0
transform 1 0 16810 0 -1 6970
box -6 -8 66 248
use NAND2X1  _11914_
timestamp 0
transform 1 0 16690 0 -1 6970
box -6 -8 86 248
use AND2X2  _11915_
timestamp 0
transform -1 0 15290 0 -1 6970
box -6 -8 106 248
use OAI21X1  _11916_
timestamp 0
transform -1 0 15130 0 -1 6970
box -6 -8 106 248
use OAI21X1  _11917_
timestamp 0
transform -1 0 14830 0 -1 6970
box -6 -8 106 248
use OAI21X1  _11918_
timestamp 0
transform 1 0 12570 0 -1 7450
box -6 -8 106 248
use INVX1  _11919_
timestamp 0
transform 1 0 14450 0 -1 6970
box -6 -8 66 248
use INVX1  _11920_
timestamp 0
transform -1 0 16470 0 1 8410
box -6 -8 66 248
use NAND3X1  _11921_
timestamp 0
transform 1 0 16610 0 -1 7930
box -6 -8 106 248
use AOI21X1  _11922_
timestamp 0
transform -1 0 15330 0 1 8890
box -6 -8 106 248
use NAND2X1  _11923_
timestamp 0
transform -1 0 15290 0 -1 8890
box -6 -8 86 248
use OAI21X1  _11924_
timestamp 0
transform 1 0 15310 0 1 8410
box -6 -8 106 248
use NAND3X1  _11925_
timestamp 0
transform -1 0 16170 0 -1 7930
box -6 -8 106 248
use INVX1  _11926_
timestamp 0
transform 1 0 16090 0 1 7450
box -6 -8 66 248
use OAI21X1  _11927_
timestamp 0
transform 1 0 16470 0 1 7450
box -6 -8 106 248
use NAND2X1  _11928_
timestamp 0
transform 1 0 16190 0 1 7450
box -6 -8 86 248
use NAND3X1  _11929_
timestamp 0
transform -1 0 16310 0 -1 7450
box -6 -8 106 248
use NAND3X1  _11930_
timestamp 0
transform -1 0 16030 0 -1 7930
box -6 -8 106 248
use NAND2X1  _11931_
timestamp 0
transform 1 0 16330 0 1 7450
box -6 -8 86 248
use NAND3X1  _11932_
timestamp 0
transform 1 0 15950 0 1 7450
box -6 -8 106 248
use NAND2X1  _11933_
timestamp 0
transform 1 0 16090 0 -1 6970
box -6 -8 86 248
use AOI21X1  _11934_
timestamp 0
transform -1 0 16770 0 -1 7450
box -6 -8 106 248
use NOR2X1  _11935_
timestamp 0
transform 1 0 16890 0 1 6970
box -6 -8 86 248
use OAI21X1  _11936_
timestamp 0
transform 1 0 16930 0 -1 6970
box -6 -8 106 248
use NAND2X1  _11937_
timestamp 0
transform 1 0 16570 0 -1 6970
box -6 -8 86 248
use AOI21X1  _11938_
timestamp 0
transform -1 0 15890 0 -1 6970
box -6 -8 106 248
use OAI21X1  _11939_
timestamp 0
transform -1 0 15730 0 -1 6970
box -6 -8 106 248
use AOI22X1  _11940_
timestamp 0
transform 1 0 14550 0 -1 6970
box -6 -8 126 248
use INVX1  _11941_
timestamp 0
transform 1 0 12890 0 1 6970
box -6 -8 66 248
use AOI21X1  _11942_
timestamp 0
transform -1 0 16150 0 -1 7450
box -6 -8 106 248
use AND2X2  _11943_
timestamp 0
transform 1 0 17030 0 1 6970
box -6 -8 106 248
use NAND3X1  _11944_
timestamp 0
transform 1 0 16750 0 1 6970
box -6 -8 106 248
use AOI21X1  _11945_
timestamp 0
transform -1 0 16710 0 1 6970
box -6 -8 106 248
use OAI21X1  _11946_
timestamp 0
transform 1 0 16470 0 1 6970
box -6 -8 106 248
use AOI21X1  _11947_
timestamp 0
transform -1 0 16090 0 1 6970
box -6 -8 106 248
use INVX1  _11948_
timestamp 0
transform -1 0 16370 0 1 8410
box -6 -8 66 248
use NAND3X1  _11949_
timestamp 0
transform -1 0 16310 0 -1 7930
box -6 -8 106 248
use INVX1  _11950_
timestamp 0
transform 1 0 14590 0 1 8890
box -6 -8 66 248
use NOR2X1  _11951_
timestamp 0
transform -1 0 15410 0 -1 8890
box -6 -8 86 248
use INVX1  _11952_
timestamp 0
transform 1 0 15450 0 -1 8890
box -6 -8 66 248
use OAI21X1  _11953_
timestamp 0
transform 1 0 15910 0 1 8410
box -6 -8 106 248
use NAND3X1  _11954_
timestamp 0
transform 1 0 15750 0 -1 8410
box -6 -8 106 248
use INVX1  _11955_
timestamp 0
transform 1 0 16610 0 -1 8410
box -6 -8 66 248
use OAI21X1  _11956_
timestamp 0
transform 1 0 16410 0 1 7930
box -6 -8 106 248
use NAND2X1  _11957_
timestamp 0
transform 1 0 16330 0 -1 8410
box -6 -8 86 248
use NAND3X1  _11958_
timestamp 0
transform 1 0 15910 0 -1 8410
box -6 -8 106 248
use NAND3X1  _11959_
timestamp 0
transform -1 0 16290 0 -1 8410
box -6 -8 106 248
use NAND2X1  _11960_
timestamp 0
transform -1 0 16550 0 -1 8410
box -6 -8 86 248
use NAND3X1  _11961_
timestamp 0
transform -1 0 16150 0 -1 8410
box -6 -8 106 248
use NAND2X1  _11962_
timestamp 0
transform 1 0 15870 0 1 6970
box -6 -8 86 248
use INVX1  _11963_
timestamp 0
transform 1 0 15630 0 1 6970
box -6 -8 66 248
use NOR2X1  _11964_
timestamp 0
transform 1 0 15730 0 1 6970
box -6 -8 86 248
use OAI21X1  _11965_
timestamp 0
transform 1 0 15950 0 -1 6970
box -6 -8 106 248
use OAI21X1  _11966_
timestamp 0
transform -1 0 15590 0 1 6970
box -6 -8 106 248
use OAI21X1  _11967_
timestamp 0
transform -1 0 13370 0 1 7930
box -6 -8 106 248
use INVX1  _11968_
timestamp 0
transform 1 0 13810 0 -1 7450
box -6 -8 66 248
use OAI21X1  _11969_
timestamp 0
transform -1 0 14470 0 1 6970
box -6 -8 106 248
use OAI21X1  _11970_
timestamp 0
transform 1 0 12990 0 1 6970
box -6 -8 106 248
use INVX1  _11971_
timestamp 0
transform 1 0 14090 0 1 6970
box -6 -8 66 248
use OAI21X1  _11972_
timestamp 0
transform 1 0 16150 0 1 6970
box -6 -8 106 248
use NOR2X1  _11973_
timestamp 0
transform 1 0 16210 0 -1 6970
box -6 -8 86 248
use AOI21X1  _11974_
timestamp 0
transform 1 0 16310 0 1 6970
box -6 -8 106 248
use INVX1  _11975_
timestamp 0
transform 1 0 15430 0 1 7450
box -6 -8 66 248
use OR2X2  _11976_
timestamp 0
transform -1 0 15810 0 1 7930
box -6 -8 106 248
use OAI21X1  _11977_
timestamp 0
transform -1 0 15850 0 1 8410
box -6 -8 106 248
use NAND3X1  _11978_
timestamp 0
transform -1 0 15670 0 1 7930
box -6 -8 106 248
use NOR2X1  _11979_
timestamp 0
transform 1 0 16030 0 1 7930
box -6 -8 86 248
use INVX1  _11980_
timestamp 0
transform 1 0 15390 0 -1 7930
box -6 -8 66 248
use OAI21X1  _11981_
timestamp 0
transform -1 0 15750 0 -1 7930
box -6 -8 106 248
use NAND3X1  _11982_
timestamp 0
transform -1 0 15350 0 -1 7930
box -6 -8 106 248
use NAND3X1  _11983_
timestamp 0
transform 1 0 15490 0 -1 7930
box -6 -8 106 248
use OAI21X1  _11984_
timestamp 0
transform -1 0 15970 0 1 7930
box -6 -8 106 248
use NAND3X1  _11985_
timestamp 0
transform 1 0 15530 0 1 7450
box -6 -8 106 248
use AND2X2  _11986_
timestamp 0
transform 1 0 15290 0 1 7450
box -6 -8 106 248
use INVX1  _11987_
timestamp 0
transform 1 0 15270 0 1 6970
box -6 -8 66 248
use AOI21X1  _11988_
timestamp 0
transform -1 0 15230 0 1 6970
box -6 -8 106 248
use OAI21X1  _11989_
timestamp 0
transform 1 0 14990 0 1 6970
box -6 -8 106 248
use AOI22X1  _11990_
timestamp 0
transform 1 0 14190 0 1 6970
box -6 -8 126 248
use NAND2X1  _11991_
timestamp 0
transform -1 0 15850 0 -1 7450
box -6 -8 86 248
use AND2X2  _11992_
timestamp 0
transform -1 0 15570 0 -1 7450
box -6 -8 106 248
use AND2X2  _11993_
timestamp 0
transform -1 0 16010 0 -1 7450
box -6 -8 106 248
use NAND3X1  _11994_
timestamp 0
transform -1 0 15710 0 -1 7450
box -6 -8 106 248
use OAI21X1  _11995_
timestamp 0
transform -1 0 15430 0 -1 7450
box -6 -8 106 248
use INVX1  _11996_
timestamp 0
transform -1 0 15230 0 1 7450
box -6 -8 66 248
use AOI21X1  _11997_
timestamp 0
transform -1 0 15130 0 -1 7450
box -6 -8 106 248
use INVX1  _11998_
timestamp 0
transform 1 0 14710 0 -1 7930
box -6 -8 66 248
use NOR3X1  _11999_
timestamp 0
transform -1 0 15710 0 -1 8410
box -6 -8 186 248
use INVX1  _12000_
timestamp 0
transform -1 0 15390 0 1 7930
box -6 -8 66 248
use OAI21X1  _12001_
timestamp 0
transform -1 0 15550 0 1 8410
box -6 -8 106 248
use NAND3X1  _12002_
timestamp 0
transform -1 0 15270 0 1 7930
box -6 -8 106 248
use INVX1  _12003_
timestamp 0
transform -1 0 15210 0 -1 8410
box -6 -8 66 248
use OAI21X1  _12004_
timestamp 0
transform -1 0 15210 0 -1 7930
box -6 -8 106 248
use NAND3X1  _12005_
timestamp 0
transform 1 0 14830 0 -1 7930
box -6 -8 106 248
use NAND3X1  _12006_
timestamp 0
transform 1 0 15030 0 1 7930
box -6 -8 106 248
use OAI21X1  _12007_
timestamp 0
transform -1 0 15530 0 1 7930
box -6 -8 106 248
use NAND3X1  _12008_
timestamp 0
transform 1 0 14730 0 1 7930
box -6 -8 106 248
use AND2X2  _12009_
timestamp 0
transform 1 0 14850 0 1 7450
box -6 -8 106 248
use AND2X2  _12010_
timestamp 0
transform -1 0 14930 0 1 6970
box -6 -8 106 248
use OAI21X1  _12011_
timestamp 0
transform -1 0 14770 0 1 6970
box -6 -8 106 248
use OAI21X1  _12012_
timestamp 0
transform -1 0 14630 0 1 6970
box -6 -8 106 248
use OAI21X1  _12013_
timestamp 0
transform 1 0 13470 0 1 6970
box -6 -8 106 248
use INVX1  _12014_
timestamp 0
transform 1 0 14670 0 -1 8410
box -6 -8 66 248
use OAI21X1  _12015_
timestamp 0
transform 1 0 15150 0 1 8410
box -6 -8 106 248
use INVX1  _12016_
timestamp 0
transform -1 0 14830 0 -1 8410
box -6 -8 66 248
use AOI21X1  _12017_
timestamp 0
transform -1 0 14990 0 1 7930
box -6 -8 106 248
use NAND3X1  _12018_
timestamp 0
transform -1 0 14970 0 -1 8410
box -6 -8 106 248
use NAND2X1  _12019_
timestamp 0
transform 1 0 14590 0 1 7930
box -6 -8 86 248
use NAND2X1  _12020_
timestamp 0
transform 1 0 14550 0 -1 8410
box -6 -8 86 248
use OAI21X1  _12021_
timestamp 0
transform -1 0 14550 0 1 7930
box -6 -8 106 248
use NAND2X1  _12022_
timestamp 0
transform 1 0 14330 0 1 7930
box -6 -8 86 248
use INVX1  _12023_
timestamp 0
transform -1 0 14350 0 -1 7930
box -6 -8 66 248
use AND2X2  _12024_
timestamp 0
transform -1 0 14650 0 -1 7930
box -6 -8 106 248
use NAND2X1  _12025_
timestamp 0
transform -1 0 14250 0 -1 7930
box -6 -8 86 248
use NAND3X1  _12026_
timestamp 0
transform -1 0 14490 0 -1 7930
box -6 -8 106 248
use NAND2X1  _12027_
timestamp 0
transform -1 0 14450 0 -1 7450
box -6 -8 86 248
use AOI21X1  _12028_
timestamp 0
transform 1 0 14970 0 -1 7930
box -6 -8 106 248
use AOI21X1  _12029_
timestamp 0
transform -1 0 15110 0 1 7450
box -6 -8 106 248
use NAND3X1  _12030_
timestamp 0
transform -1 0 14750 0 -1 7450
box -6 -8 106 248
use AOI21X1  _12031_
timestamp 0
transform -1 0 14610 0 -1 7450
box -6 -8 106 248
use AND2X2  _12032_
timestamp 0
transform 1 0 14410 0 1 7450
box -6 -8 106 248
use NAND3X1  _12033_
timestamp 0
transform -1 0 14810 0 1 7450
box -6 -8 106 248
use OAI21X1  _12034_
timestamp 0
transform -1 0 14670 0 1 7450
box -6 -8 106 248
use OAI21X1  _12035_
timestamp 0
transform 1 0 14270 0 1 7450
box -6 -8 106 248
use OR2X2  _12036_
timestamp 0
transform -1 0 14190 0 -1 7450
box -6 -8 106 248
use AOI22X1  _12037_
timestamp 0
transform 1 0 13910 0 -1 7450
box -6 -8 126 248
use NAND2X1  _12038_
timestamp 0
transform -1 0 13110 0 -1 7930
box -6 -8 86 248
use INVX1  _12039_
timestamp 0
transform -1 0 14310 0 -1 7450
box -6 -8 66 248
use NAND2X1  _12040_
timestamp 0
transform 1 0 14690 0 -1 8890
box -6 -8 86 248
use INVX1  _12041_
timestamp 0
transform 1 0 14830 0 -1 8890
box -6 -8 66 248
use NAND2X1  _12042_
timestamp 0
transform -1 0 14510 0 -1 9370
box -6 -8 86 248
use NAND2X1  _12043_
timestamp 0
transform -1 0 14650 0 -1 9370
box -6 -8 86 248
use INVX1  _12044_
timestamp 0
transform 1 0 14230 0 1 8890
box -6 -8 66 248
use NAND2X1  _12045_
timestamp 0
transform -1 0 14270 0 1 7930
box -6 -8 86 248
use NAND2X1  _12046_
timestamp 0
transform -1 0 14150 0 1 7930
box -6 -8 86 248
use NAND2X1  _12047_
timestamp 0
transform -1 0 14010 0 1 7930
box -6 -8 86 248
use INVX1  _12048_
timestamp 0
transform 1 0 13850 0 -1 7930
box -6 -8 66 248
use NOR3X1  _12049_
timestamp 0
transform -1 0 14130 0 -1 7930
box -6 -8 186 248
use AOI21X1  _12050_
timestamp 0
transform -1 0 14230 0 1 7450
box -6 -8 106 248
use OAI21X1  _12051_
timestamp 0
transform -1 0 13790 0 -1 7930
box -6 -8 106 248
use OAI21X1  _12052_
timestamp 0
transform -1 0 13630 0 -1 7930
box -6 -8 106 248
use NAND2X1  _12053_
timestamp 0
transform 1 0 13410 0 -1 7930
box -6 -8 86 248
use NAND2X1  _12054_
timestamp 0
transform 1 0 12870 0 -1 10810
box -6 -8 86 248
use INVX1  _12055_
timestamp 0
transform -1 0 15910 0 -1 8890
box -6 -8 66 248
use NAND2X1  _12056_
timestamp 0
transform 1 0 16050 0 1 8410
box -6 -8 86 248
use OAI21X1  _12057_
timestamp 0
transform 1 0 15950 0 -1 8890
box -6 -8 106 248
use NAND2X1  _12058_
timestamp 0
transform -1 0 16130 0 -1 9370
box -6 -8 86 248
use NOR2X1  _12059_
timestamp 0
transform -1 0 12650 0 1 9370
box -6 -8 86 248
use NOR2X1  _12060_
timestamp 0
transform 1 0 12890 0 -1 9370
box -6 -8 86 248
use AOI22X1  _12061_
timestamp 0
transform -1 0 12730 0 -1 9370
box -6 -8 126 248
use NAND3X1  _12062_
timestamp 0
transform 1 0 16190 0 -1 9370
box -6 -8 106 248
use NAND2X1  _12063_
timestamp 0
transform 1 0 16510 0 1 8410
box -6 -8 86 248
use OAI21X1  _12064_
timestamp 0
transform -1 0 16730 0 1 8410
box -6 -8 106 248
use NAND2X1  _12065_
timestamp 0
transform -1 0 17150 0 1 8890
box -6 -8 86 248
use OAI21X1  _12066_
timestamp 0
transform 1 0 17050 0 -1 8890
box -6 -8 106 248
use MUX2X1  _12067_
timestamp 0
transform 1 0 16750 0 1 9850
box -6 -8 126 248
use NAND2X1  _12068_
timestamp 0
transform 1 0 16690 0 -1 10330
box -6 -8 86 248
use AND2X2  _12069_
timestamp 0
transform -1 0 16350 0 -1 10330
box -6 -8 106 248
use NOR2X1  _12070_
timestamp 0
transform 1 0 12890 0 1 10330
box -6 -8 86 248
use NAND2X1  _12071_
timestamp 0
transform 1 0 17050 0 1 9850
box -6 -8 86 248
use NAND2X1  _12072_
timestamp 0
transform -1 0 17010 0 1 9850
box -6 -8 86 248
use NAND2X1  _12073_
timestamp 0
transform 1 0 17090 0 -1 10330
box -6 -8 86 248
use OAI21X1  _12074_
timestamp 0
transform -1 0 17050 0 -1 10330
box -6 -8 106 248
use OAI21X1  _12075_
timestamp 0
transform -1 0 13110 0 1 10330
box -6 -8 106 248
use OAI21X1  _12076_
timestamp 0
transform -1 0 12830 0 1 10330
box -6 -8 106 248
use NAND2X1  _12077_
timestamp 0
transform -1 0 12670 0 1 10810
box -6 -8 86 248
use NOR2X1  _12078_
timestamp 0
transform -1 0 13230 0 1 10330
box -6 -8 86 248
use NAND2X1  _12079_
timestamp 0
transform 1 0 15610 0 -1 17050
box -6 -8 86 248
use OAI21X1  _12080_
timestamp 0
transform 1 0 17010 0 1 8410
box -6 -8 106 248
use NAND2X1  _12081_
timestamp 0
transform 1 0 13830 0 1 8890
box -6 -8 86 248
use OAI21X1  _12082_
timestamp 0
transform 1 0 13670 0 1 8890
box -6 -8 106 248
use MUX2X1  _12083_
timestamp 0
transform -1 0 16850 0 -1 9370
box -6 -8 126 248
use NAND2X1  _12084_
timestamp 0
transform 1 0 16610 0 -1 9370
box -6 -8 86 248
use NAND2X1  _12085_
timestamp 0
transform -1 0 16170 0 -1 8890
box -6 -8 86 248
use OAI21X1  _12086_
timestamp 0
transform -1 0 16330 0 -1 8890
box -6 -8 106 248
use INVX1  _12087_
timestamp 0
transform -1 0 16770 0 -1 9850
box -6 -8 66 248
use NAND2X1  _12088_
timestamp 0
transform 1 0 16490 0 -1 8890
box -6 -8 86 248
use OAI21X1  _12089_
timestamp 0
transform 1 0 16790 0 -1 8890
box -6 -8 106 248
use NAND2X1  _12090_
timestamp 0
transform 1 0 16990 0 -1 11770
box -6 -8 86 248
use OAI21X1  _12091_
timestamp 0
transform 1 0 16830 0 -1 9850
box -6 -8 106 248
use OAI21X1  _12092_
timestamp 0
transform 1 0 16570 0 -1 9850
box -6 -8 106 248
use NAND3X1  _12093_
timestamp 0
transform -1 0 15550 0 -1 10330
box -6 -8 106 248
use MUX2X1  _12094_
timestamp 0
transform 1 0 16730 0 1 9370
box -6 -8 126 248
use MUX2X1  _12095_
timestamp 0
transform -1 0 16690 0 1 9370
box -6 -8 126 248
use OAI21X1  _12096_
timestamp 0
transform 1 0 16410 0 -1 10330
box -6 -8 106 248
use AOI21X1  _12097_
timestamp 0
transform -1 0 15250 0 -1 10330
box -6 -8 106 248
use INVX1  _12098_
timestamp 0
transform -1 0 15250 0 1 10330
box -6 -8 66 248
use NAND3X1  _12099_
timestamp 0
transform 1 0 15290 0 -1 10330
box -6 -8 106 248
use AND2X2  _12100_
timestamp 0
transform -1 0 15130 0 1 10330
box -6 -8 106 248
use NAND2X1  _12101_
timestamp 0
transform 1 0 13830 0 1 10330
box -6 -8 86 248
use OR2X2  _12102_
timestamp 0
transform -1 0 13770 0 1 10330
box -6 -8 106 248
use AOI21X1  _12103_
timestamp 0
transform -1 0 13630 0 1 10330
box -6 -8 106 248
use OAI21X1  _12104_
timestamp 0
transform -1 0 12810 0 1 10810
box -6 -8 106 248
use NAND2X1  _12105_
timestamp 0
transform -1 0 13270 0 -1 10810
box -6 -8 86 248
use AOI21X1  _12106_
timestamp 0
transform 1 0 15290 0 1 10330
box -6 -8 106 248
use NAND2X1  _12107_
timestamp 0
transform -1 0 16910 0 1 10330
box -6 -8 86 248
use NAND2X1  _12108_
timestamp 0
transform -1 0 15650 0 -1 8890
box -6 -8 86 248
use OAI21X1  _12109_
timestamp 0
transform -1 0 15790 0 -1 8890
box -6 -8 106 248
use NAND2X1  _12110_
timestamp 0
transform 1 0 16610 0 1 9850
box -6 -8 86 248
use OAI21X1  _12111_
timestamp 0
transform 1 0 16170 0 1 9850
box -6 -8 106 248
use NAND2X1  _12112_
timestamp 0
transform -1 0 16430 0 -1 9370
box -6 -8 86 248
use NAND2X1  _12113_
timestamp 0
transform 1 0 16910 0 1 250
box -6 -8 86 248
use NAND2X1  _12114_
timestamp 0
transform -1 0 16550 0 -1 9370
box -6 -8 86 248
use AOI21X1  _12115_
timestamp 0
transform 1 0 16410 0 1 10330
box -6 -8 106 248
use INVX1  _12116_
timestamp 0
transform 1 0 16950 0 -1 10810
box -6 -8 66 248
use NAND3X1  _12117_
timestamp 0
transform -1 0 16910 0 -1 10810
box -6 -8 106 248
use AOI21X1  _12118_
timestamp 0
transform 1 0 16550 0 -1 10330
box -6 -8 106 248
use OAI21X1  _12119_
timestamp 0
transform 1 0 16650 0 -1 10810
box -6 -8 106 248
use NAND3X1  _12120_
timestamp 0
transform 1 0 16510 0 -1 10810
box -6 -8 106 248
use INVX1  _12121_
timestamp 0
transform -1 0 16150 0 -1 10810
box -6 -8 66 248
use AOI21X1  _12122_
timestamp 0
transform 1 0 16350 0 -1 10810
box -6 -8 106 248
use NOR2X1  _12123_
timestamp 0
transform -1 0 16050 0 -1 10810
box -6 -8 86 248
use AND2X2  _12124_
timestamp 0
transform -1 0 15810 0 -1 10810
box -6 -8 106 248
use NOR2X1  _12125_
timestamp 0
transform 1 0 15850 0 -1 10810
box -6 -8 86 248
use OAI21X1  _12126_
timestamp 0
transform -1 0 15650 0 -1 10810
box -6 -8 106 248
use OAI21X1  _12127_
timestamp 0
transform -1 0 13430 0 -1 10810
box -6 -8 106 248
use OAI21X1  _12128_
timestamp 0
transform 1 0 16190 0 -1 10810
box -6 -8 106 248
use INVX1  _12129_
timestamp 0
transform 1 0 17070 0 1 11290
box -6 -8 66 248
use NAND2X1  _12130_
timestamp 0
transform -1 0 15090 0 -1 8410
box -6 -8 86 248
use OAI21X1  _12131_
timestamp 0
transform 1 0 15390 0 -1 8410
box -6 -8 106 248
use MUX2X1  _12132_
timestamp 0
transform -1 0 16390 0 -1 9850
box -6 -8 126 248
use NOR2X1  _12133_
timestamp 0
transform -1 0 16890 0 -1 10330
box -6 -8 86 248
use NAND2X1  _12134_
timestamp 0
transform 1 0 16910 0 -1 9370
box -6 -8 86 248
use NAND2X1  _12135_
timestamp 0
transform 1 0 17030 0 -1 9370
box -6 -8 86 248
use NAND2X1  _12136_
timestamp 0
transform 1 0 16910 0 1 9370
box -6 -8 86 248
use OR2X2  _12137_
timestamp 0
transform 1 0 16930 0 1 10810
box -6 -8 106 248
use OAI21X1  _12138_
timestamp 0
transform 1 0 17050 0 -1 10810
box -6 -8 106 248
use OR2X2  _12139_
timestamp 0
transform 1 0 17090 0 1 10810
box -6 -8 106 248
use OAI21X1  _12140_
timestamp 0
transform 1 0 16790 0 1 10810
box -6 -8 106 248
use AOI21X1  _12141_
timestamp 0
transform -1 0 16670 0 -1 11290
box -6 -8 106 248
use INVX1  _12142_
timestamp 0
transform 1 0 16550 0 1 11290
box -6 -8 66 248
use NAND3X1  _12143_
timestamp 0
transform 1 0 16730 0 -1 11290
box -6 -8 106 248
use NAND2X1  _12144_
timestamp 0
transform 1 0 16650 0 1 11290
box -6 -8 86 248
use OR2X2  _12145_
timestamp 0
transform 1 0 16910 0 1 11290
box -6 -8 106 248
use NAND2X1  _12146_
timestamp 0
transform 1 0 16790 0 1 11290
box -6 -8 86 248
use NAND2X1  _12147_
timestamp 0
transform 1 0 16870 0 -1 11770
box -6 -8 86 248
use AOI22X1  _12148_
timestamp 0
transform 1 0 14410 0 1 11770
box -6 -8 126 248
use AOI21X1  _12149_
timestamp 0
transform 1 0 16410 0 1 11290
box -6 -8 106 248
use NAND2X1  _12150_
timestamp 0
transform -1 0 15010 0 -1 8890
box -6 -8 86 248
use OAI21X1  _12151_
timestamp 0
transform 1 0 15070 0 -1 8890
box -6 -8 106 248
use NAND2X1  _12152_
timestamp 0
transform -1 0 15730 0 1 9850
box -6 -8 86 248
use OAI21X1  _12153_
timestamp 0
transform -1 0 15990 0 1 9850
box -6 -8 106 248
use NAND2X1  _12154_
timestamp 0
transform -1 0 16630 0 1 10330
box -6 -8 86 248
use OAI21X1  _12155_
timestamp 0
transform 1 0 16690 0 1 10330
box -6 -8 106 248
use INVX1  _12156_
timestamp 0
transform 1 0 17110 0 -1 11770
box -6 -8 66 248
use NAND3X1  _12157_
timestamp 0
transform 1 0 16950 0 1 10330
box -6 -8 106 248
use OAI21X1  _12158_
timestamp 0
transform 1 0 17030 0 -1 11290
box -6 -8 106 248
use OR2X2  _12159_
timestamp 0
transform -1 0 16970 0 1 11770
box -6 -8 106 248
use NOR2X1  _12160_
timestamp 0
transform 1 0 16890 0 -1 11290
box -6 -8 86 248
use OAI21X1  _12161_
timestamp 0
transform 1 0 16730 0 -1 11770
box -6 -8 106 248
use NAND3X1  _12162_
timestamp 0
transform 1 0 16730 0 1 11770
box -6 -8 106 248
use OR2X2  _12163_
timestamp 0
transform 1 0 17030 0 1 11770
box -6 -8 106 248
use OAI21X1  _12164_
timestamp 0
transform -1 0 16690 0 -1 11770
box -6 -8 106 248
use NAND3X1  _12165_
timestamp 0
transform -1 0 16690 0 1 11770
box -6 -8 106 248
use NAND2X1  _12166_
timestamp 0
transform -1 0 16230 0 1 11770
box -6 -8 86 248
use OR2X2  _12167_
timestamp 0
transform -1 0 15470 0 1 11770
box -6 -8 106 248
use NAND2X1  _12168_
timestamp 0
transform 1 0 15510 0 1 11770
box -6 -8 86 248
use NAND2X1  _12169_
timestamp 0
transform 1 0 15230 0 1 11770
box -6 -8 86 248
use AOI22X1  _12170_
timestamp 0
transform 1 0 13830 0 1 11770
box -6 -8 126 248
use INVX1  _12171_
timestamp 0
transform 1 0 13990 0 1 11770
box -6 -8 66 248
use OAI21X1  _12172_
timestamp 0
transform 1 0 15890 0 1 11770
box -6 -8 106 248
use NAND2X1  _12173_
timestamp 0
transform -1 0 16210 0 1 11290
box -6 -8 86 248
use NOR2X1  _12174_
timestamp 0
transform -1 0 16070 0 -1 9850
box -6 -8 86 248
use AOI21X1  _12175_
timestamp 0
transform 1 0 16110 0 -1 9850
box -6 -8 106 248
use NAND2X1  _12176_
timestamp 0
transform 1 0 16470 0 1 9850
box -6 -8 86 248
use OAI21X1  _12177_
timestamp 0
transform 1 0 16330 0 1 9850
box -6 -8 106 248
use INVX1  _12178_
timestamp 0
transform 1 0 16170 0 -1 11290
box -6 -8 66 248
use NAND3X1  _12179_
timestamp 0
transform 1 0 16270 0 1 11290
box -6 -8 106 248
use NOR2X1  _12180_
timestamp 0
transform -1 0 16750 0 1 10810
box -6 -8 86 248
use NAND3X1  _12181_
timestamp 0
transform -1 0 16630 0 1 10810
box -6 -8 106 248
use OAI21X1  _12182_
timestamp 0
transform -1 0 16510 0 -1 11290
box -6 -8 106 248
use NAND2X1  _12183_
timestamp 0
transform -1 0 16350 0 -1 11290
box -6 -8 86 248
use AOI21X1  _12184_
timestamp 0
transform -1 0 16390 0 -1 11770
box -6 -8 106 248
use INVX1  _12185_
timestamp 0
transform -1 0 16070 0 -1 11770
box -6 -8 66 248
use NAND3X1  _12186_
timestamp 0
transform -1 0 16550 0 -1 11770
box -6 -8 106 248
use NAND2X1  _12187_
timestamp 0
transform -1 0 15550 0 -1 11770
box -6 -8 86 248
use NOR2X1  _12188_
timestamp 0
transform 1 0 15110 0 1 11770
box -6 -8 86 248
use AND2X2  _12189_
timestamp 0
transform -1 0 15070 0 1 11770
box -6 -8 106 248
use OAI21X1  _12190_
timestamp 0
transform -1 0 14910 0 1 11770
box -6 -8 106 248
use OAI21X1  _12191_
timestamp 0
transform 1 0 14110 0 1 11770
box -6 -8 106 248
use INVX1  _12192_
timestamp 0
transform 1 0 12670 0 -1 11770
box -6 -8 66 248
use NAND3X1  _12193_
timestamp 0
transform -1 0 16090 0 1 11290
box -6 -8 106 248
use AOI21X1  _12194_
timestamp 0
transform 1 0 16030 0 1 9850
box -6 -8 106 248
use NAND2X1  _12195_
timestamp 0
transform -1 0 16210 0 -1 10330
box -6 -8 86 248
use OAI21X1  _12196_
timestamp 0
transform -1 0 16350 0 1 10330
box -6 -8 106 248
use NAND3X1  _12197_
timestamp 0
transform 1 0 15670 0 1 11290
box -6 -8 106 248
use NOR3X1  _12198_
timestamp 0
transform -1 0 16490 0 1 10810
box -6 -8 186 248
use INVX1  _12199_
timestamp 0
transform 1 0 15930 0 -1 11290
box -6 -8 66 248
use OAI21X1  _12200_
timestamp 0
transform -1 0 16130 0 -1 11290
box -6 -8 106 248
use NAND2X1  _12201_
timestamp 0
transform 1 0 15430 0 1 11290
box -6 -8 86 248
use NAND2X1  _12202_
timestamp 0
transform 1 0 15290 0 1 11290
box -6 -8 86 248
use NAND3X1  _12203_
timestamp 0
transform 1 0 15150 0 1 11290
box -6 -8 106 248
use NAND2X1  _12204_
timestamp 0
transform -1 0 15090 0 1 11290
box -6 -8 86 248
use AOI21X1  _12205_
timestamp 0
transform -1 0 16530 0 1 11770
box -6 -8 106 248
use NOR2X1  _12206_
timestamp 0
transform -1 0 16110 0 1 11770
box -6 -8 86 248
use OAI21X1  _12207_
timestamp 0
transform 1 0 15730 0 1 11770
box -6 -8 106 248
use NAND2X1  _12208_
timestamp 0
transform 1 0 15610 0 -1 11770
box -6 -8 86 248
use NOR2X1  _12209_
timestamp 0
transform 1 0 15350 0 -1 11770
box -6 -8 86 248
use AND2X2  _12210_
timestamp 0
transform -1 0 15310 0 -1 11770
box -6 -8 106 248
use AND2X2  _12211_
timestamp 0
transform -1 0 16370 0 1 11770
box -6 -8 106 248
use NAND3X1  _12212_
timestamp 0
transform -1 0 15970 0 -1 11770
box -6 -8 106 248
use AOI21X1  _12213_
timestamp 0
transform -1 0 16230 0 -1 11770
box -6 -8 106 248
use OAI21X1  _12214_
timestamp 0
transform -1 0 15830 0 -1 11770
box -6 -8 106 248
use NOR2X1  _12215_
timestamp 0
transform -1 0 15150 0 -1 11770
box -6 -8 86 248
use OAI21X1  _12216_
timestamp 0
transform -1 0 15010 0 -1 11770
box -6 -8 106 248
use NAND2X1  _12217_
timestamp 0
transform 1 0 13170 0 -1 11770
box -6 -8 86 248
use OAI21X1  _12218_
timestamp 0
transform 1 0 13010 0 -1 11770
box -6 -8 106 248
use INVX1  _12219_
timestamp 0
transform 1 0 13990 0 -1 11770
box -6 -8 66 248
use INVX1  _12220_
timestamp 0
transform -1 0 14870 0 -1 11770
box -6 -8 66 248
use NAND2X1  _12221_
timestamp 0
transform 1 0 16170 0 1 10810
box -6 -8 86 248
use NOR2X1  _12222_
timestamp 0
transform 1 0 15850 0 -1 9850
box -6 -8 86 248
use INVX1  _12223_
timestamp 0
transform -1 0 15830 0 1 9850
box -6 -8 66 248
use OAI21X1  _12224_
timestamp 0
transform -1 0 16090 0 -1 10330
box -6 -8 106 248
use NAND3X1  _12225_
timestamp 0
transform 1 0 15490 0 1 10810
box -6 -8 106 248
use INVX1  _12226_
timestamp 0
transform 1 0 15830 0 -1 11290
box -6 -8 66 248
use OAI21X1  _12227_
timestamp 0
transform -1 0 15930 0 1 11290
box -6 -8 106 248
use NAND2X1  _12228_
timestamp 0
transform -1 0 15670 0 -1 11290
box -6 -8 86 248
use NAND3X1  _12229_
timestamp 0
transform -1 0 15550 0 -1 11290
box -6 -8 106 248
use NAND3X1  _12230_
timestamp 0
transform -1 0 15990 0 1 10810
box -6 -8 106 248
use NAND2X1  _12231_
timestamp 0
transform -1 0 15790 0 -1 11290
box -6 -8 86 248
use NAND3X1  _12232_
timestamp 0
transform -1 0 15850 0 1 10810
box -6 -8 106 248
use NAND2X1  _12233_
timestamp 0
transform 1 0 15550 0 1 11290
box -6 -8 86 248
use OAI21X1  _12234_
timestamp 0
transform -1 0 14630 0 -1 11770
box -6 -8 106 248
use NOR2X1  _12235_
timestamp 0
transform 1 0 14670 0 -1 11770
box -6 -8 86 248
use INVX1  _12236_
timestamp 0
transform -1 0 14470 0 -1 11770
box -6 -8 66 248
use AOI21X1  _12237_
timestamp 0
transform -1 0 14350 0 -1 11770
box -6 -8 106 248
use AOI22X1  _12238_
timestamp 0
transform 1 0 14090 0 -1 11770
box -6 -8 126 248
use OAI21X1  _12239_
timestamp 0
transform 1 0 14870 0 1 11290
box -6 -8 106 248
use NOR2X1  _12240_
timestamp 0
transform -1 0 14810 0 1 11290
box -6 -8 86 248
use AOI21X1  _12241_
timestamp 0
transform -1 0 14690 0 1 11290
box -6 -8 106 248
use INVX1  _12242_
timestamp 0
transform -1 0 14490 0 1 10810
box -6 -8 66 248
use NAND3X1  _12243_
timestamp 0
transform 1 0 16030 0 1 10810
box -6 -8 106 248
use INVX1  _12244_
timestamp 0
transform -1 0 16190 0 1 10330
box -6 -8 66 248
use OAI21X1  _12245_
timestamp 0
transform -1 0 16070 0 1 10330
box -6 -8 106 248
use INVX1  _12246_
timestamp 0
transform -1 0 15290 0 1 10810
box -6 -8 66 248
use NAND3X1  _12247_
timestamp 0
transform -1 0 14930 0 1 10810
box -6 -8 106 248
use OAI21X1  _12248_
timestamp 0
transform -1 0 15450 0 1 10810
box -6 -8 106 248
use NAND2X1  _12249_
timestamp 0
transform -1 0 15170 0 1 10810
box -6 -8 86 248
use AOI21X1  _12250_
timestamp 0
transform -1 0 14630 0 1 10810
box -6 -8 106 248
use NAND3X1  _12251_
timestamp 0
transform -1 0 15350 0 -1 10810
box -6 -8 106 248
use NAND2X1  _12252_
timestamp 0
transform 1 0 14970 0 1 10810
box -6 -8 86 248
use AOI21X1  _12253_
timestamp 0
transform -1 0 14790 0 1 10810
box -6 -8 106 248
use OAI21X1  _12254_
timestamp 0
transform -1 0 14250 0 1 11290
box -6 -8 106 248
use INVX1  _12255_
timestamp 0
transform -1 0 13830 0 1 11290
box -6 -8 66 248
use OR2X2  _12256_
timestamp 0
transform -1 0 14390 0 1 11290
box -6 -8 106 248
use OAI21X1  _12257_
timestamp 0
transform -1 0 13970 0 1 11290
box -6 -8 106 248
use OAI22X1  _12258_
timestamp 0
transform 1 0 13590 0 1 11290
box -6 -8 126 248
use NAND2X1  _12259_
timestamp 0
transform -1 0 13570 0 1 10810
box -6 -8 86 248
use NOR2X1  _12260_
timestamp 0
transform -1 0 14110 0 1 11290
box -6 -8 86 248
use NOR2X1  _12261_
timestamp 0
transform -1 0 14170 0 -1 11290
box -6 -8 86 248
use OAI21X1  _12262_
timestamp 0
transform 1 0 15830 0 -1 10330
box -6 -8 106 248
use INVX1  _12263_
timestamp 0
transform 1 0 14930 0 1 10330
box -6 -8 66 248
use OAI21X1  _12264_
timestamp 0
transform -1 0 15190 0 -1 10810
box -6 -8 106 248
use NAND2X1  _12265_
timestamp 0
transform 1 0 14970 0 -1 10810
box -6 -8 86 248
use OR2X2  _12266_
timestamp 0
transform -1 0 14910 0 -1 10810
box -6 -8 106 248
use NAND3X1  _12267_
timestamp 0
transform -1 0 14650 0 -1 10810
box -6 -8 106 248
use NAND2X1  _12268_
timestamp 0
transform 1 0 14690 0 -1 10810
box -6 -8 86 248
use NAND2X1  _12269_
timestamp 0
transform 1 0 14650 0 1 10330
box -6 -8 86 248
use NAND2X1  _12270_
timestamp 0
transform 1 0 14310 0 1 10810
box -6 -8 86 248
use AND2X2  _12271_
timestamp 0
transform -1 0 14090 0 1 10810
box -6 -8 106 248
use OAI21X1  _12272_
timestamp 0
transform 1 0 14150 0 1 10810
box -6 -8 106 248
use OAI21X1  _12273_
timestamp 0
transform -1 0 13950 0 1 10810
box -6 -8 106 248
use INVX1  _12274_
timestamp 0
transform 1 0 13410 0 -1 11290
box -6 -8 66 248
use INVX1  _12275_
timestamp 0
transform -1 0 14290 0 -1 11290
box -6 -8 66 248
use AOI21X1  _12276_
timestamp 0
transform 1 0 14330 0 -1 11290
box -6 -8 106 248
use NOR2X1  _12277_
timestamp 0
transform -1 0 14530 0 1 11290
box -6 -8 86 248
use NAND3X1  _12278_
timestamp 0
transform 1 0 14630 0 -1 11290
box -6 -8 106 248
use OAI21X1  _12279_
timestamp 0
transform -1 0 14590 0 -1 11290
box -6 -8 106 248
use OAI21X1  _12280_
timestamp 0
transform 1 0 15690 0 -1 10330
box -6 -8 106 248
use INVX1  _12281_
timestamp 0
transform -1 0 15650 0 -1 10330
box -6 -8 66 248
use OR2X2  _12282_
timestamp 0
transform 1 0 15410 0 -1 10810
box -6 -8 106 248
use OAI21X1  _12283_
timestamp 0
transform -1 0 14870 0 1 10330
box -6 -8 106 248
use NAND2X1  _12284_
timestamp 0
transform 1 0 14530 0 1 10330
box -6 -8 86 248
use OR2X2  _12285_
timestamp 0
transform -1 0 14690 0 -1 10330
box -6 -8 106 248
use NAND3X1  _12286_
timestamp 0
transform 1 0 14450 0 -1 10330
box -6 -8 106 248
use AND2X2  _12287_
timestamp 0
transform -1 0 14350 0 1 10330
box -6 -8 106 248
use NOR2X1  _12288_
timestamp 0
transform 1 0 14390 0 1 10330
box -6 -8 86 248
use OAI21X1  _12289_
timestamp 0
transform -1 0 14210 0 1 10330
box -6 -8 106 248
use NAND2X1  _12290_
timestamp 0
transform 1 0 14290 0 -1 10810
box -6 -8 86 248
use AND2X2  _12291_
timestamp 0
transform -1 0 13930 0 -1 11290
box -6 -8 106 248
use NOR2X1  _12292_
timestamp 0
transform 1 0 13970 0 -1 11290
box -6 -8 86 248
use NOR2X1  _12293_
timestamp 0
transform -1 0 13770 0 -1 11290
box -6 -8 86 248
use AOI22X1  _12294_
timestamp 0
transform 1 0 13530 0 -1 11290
box -6 -8 126 248
use NAND2X1  _12295_
timestamp 0
transform -1 0 13210 0 1 10810
box -6 -8 86 248
use INVX1  _12296_
timestamp 0
transform -1 0 14490 0 -1 10810
box -6 -8 66 248
use AOI21X1  _12297_
timestamp 0
transform -1 0 14250 0 -1 10810
box -6 -8 106 248
use NAND2X1  _12298_
timestamp 0
transform 1 0 14310 0 -1 9850
box -6 -8 86 248
use NOR2X1  _12299_
timestamp 0
transform 1 0 14170 0 -1 9850
box -6 -8 86 248
use AOI21X1  _12300_
timestamp 0
transform 1 0 14290 0 -1 10330
box -6 -8 106 248
use NOR2X1  _12301_
timestamp 0
transform -1 0 14250 0 -1 10330
box -6 -8 86 248
use AND2X2  _12302_
timestamp 0
transform -1 0 14110 0 -1 10810
box -6 -8 106 248
use OAI21X1  _12303_
timestamp 0
transform -1 0 13970 0 -1 10810
box -6 -8 106 248
use OAI21X1  _12304_
timestamp 0
transform -1 0 13810 0 -1 10810
box -6 -8 106 248
use OAI21X1  _12305_
timestamp 0
transform -1 0 12010 0 1 9370
box -6 -8 106 248
use OAI21X1  _12306_
timestamp 0
transform 1 0 10710 0 1 9370
box -6 -8 106 248
use INVX1  _12307_
timestamp 0
transform 1 0 10850 0 1 9370
box -6 -8 66 248
use NOR2X1  _12308_
timestamp 0
transform -1 0 11050 0 1 9370
box -6 -8 86 248
use NAND2X1  _12309_
timestamp 0
transform 1 0 11090 0 1 9370
box -6 -8 86 248
use NAND2X1  _12310_
timestamp 0
transform 1 0 11230 0 1 9370
box -6 -8 86 248
use NAND2X1  _12311_
timestamp 0
transform 1 0 11530 0 1 9850
box -6 -8 86 248
use OAI21X1  _12312_
timestamp 0
transform 1 0 11290 0 -1 9850
box -6 -8 106 248
use NAND2X1  _12313_
timestamp 0
transform -1 0 11370 0 1 8890
box -6 -8 86 248
use INVX1  _12314_
timestamp 0
transform -1 0 11010 0 -1 9370
box -6 -8 66 248
use NOR2X1  _12315_
timestamp 0
transform 1 0 10770 0 -1 9850
box -6 -8 86 248
use AOI21X1  _12316_
timestamp 0
transform -1 0 10710 0 -1 9850
box -6 -8 106 248
use NOR2X1  _12317_
timestamp 0
transform -1 0 10150 0 1 9370
box -6 -8 86 248
use OAI21X1  _12318_
timestamp 0
transform -1 0 10430 0 1 9370
box -6 -8 106 248
use AND2X2  _12319_
timestamp 0
transform -1 0 10290 0 1 9370
box -6 -8 106 248
use OR2X2  _12320_
timestamp 0
transform 1 0 10290 0 -1 9370
box -6 -8 106 248
use OR2X2  _12321_
timestamp 0
transform -1 0 10310 0 1 8890
box -6 -8 106 248
use OAI21X1  _12322_
timestamp 0
transform -1 0 10230 0 -1 9370
box -6 -8 106 248
use NAND2X1  _12323_
timestamp 0
transform -1 0 10170 0 1 8890
box -6 -8 86 248
use NOR2X1  _12324_
timestamp 0
transform -1 0 10950 0 1 8890
box -6 -8 86 248
use NAND2X1  _12325_
timestamp 0
transform -1 0 10830 0 1 8890
box -6 -8 86 248
use NAND2X1  _12326_
timestamp 0
transform -1 0 11070 0 1 8890
box -6 -8 86 248
use OAI21X1  _12327_
timestamp 0
transform 1 0 11130 0 1 8890
box -6 -8 106 248
use INVX1  _12328_
timestamp 0
transform 1 0 10470 0 1 8890
box -6 -8 66 248
use OAI21X1  _12329_
timestamp 0
transform 1 0 10590 0 1 8890
box -6 -8 106 248
use OAI21X1  _12330_
timestamp 0
transform -1 0 12570 0 -1 9370
box -6 -8 106 248
use OAI21X1  _12331_
timestamp 0
transform -1 0 11630 0 -1 8890
box -6 -8 106 248
use MUX2X1  _12332_
timestamp 0
transform -1 0 11810 0 -1 8890
box -6 -8 126 248
use NAND2X1  _12333_
timestamp 0
transform 1 0 11250 0 1 8410
box -6 -8 86 248
use OR2X2  _12334_
timestamp 0
transform -1 0 11210 0 1 8410
box -6 -8 106 248
use NAND2X1  _12335_
timestamp 0
transform 1 0 10970 0 1 8410
box -6 -8 86 248
use INVX1  _12336_
timestamp 0
transform -1 0 10930 0 1 8410
box -6 -8 66 248
use NOR2X1  _12337_
timestamp 0
transform -1 0 10430 0 1 8890
box -6 -8 86 248
use NAND2X1  _12338_
timestamp 0
transform -1 0 10490 0 -1 8890
box -6 -8 86 248
use NAND2X1  _12339_
timestamp 0
transform 1 0 10290 0 -1 8890
box -6 -8 86 248
use OAI22X1  _12340_
timestamp 0
transform 1 0 10110 0 -1 8890
box -6 -8 126 248
use NOR2X1  _12341_
timestamp 0
transform 1 0 11190 0 -1 10330
box -6 -8 86 248
use NAND2X1  _12342_
timestamp 0
transform -1 0 10730 0 -1 8890
box -6 -8 86 248
use INVX1  _12343_
timestamp 0
transform 1 0 11030 0 -1 9850
box -6 -8 66 248
use INVX1  _12344_
timestamp 0
transform 1 0 11690 0 -1 9850
box -6 -8 66 248
use NOR2X1  _12345_
timestamp 0
transform 1 0 12630 0 -1 9850
box -6 -8 86 248
use OAI21X1  _12346_
timestamp 0
transform -1 0 12450 0 -1 9850
box -6 -8 106 248
use OAI21X1  _12347_
timestamp 0
transform 1 0 11950 0 1 9850
box -6 -8 106 248
use OAI21X1  _12348_
timestamp 0
transform -1 0 12150 0 -1 9850
box -6 -8 106 248
use NOR2X1  _12349_
timestamp 0
transform 1 0 11550 0 -1 9850
box -6 -8 86 248
use NAND2X1  _12350_
timestamp 0
transform -1 0 11510 0 -1 9850
box -6 -8 86 248
use INVX1  _12351_
timestamp 0
transform -1 0 10710 0 1 9850
box -6 -8 66 248
use NOR2X1  _12352_
timestamp 0
transform -1 0 10830 0 1 9850
box -6 -8 86 248
use OAI21X1  _12353_
timestamp 0
transform 1 0 11150 0 -1 9850
box -6 -8 106 248
use AOI21X1  _12354_
timestamp 0
transform 1 0 11150 0 1 9850
box -6 -8 106 248
use NOR2X1  _12355_
timestamp 0
transform -1 0 11130 0 -1 10330
box -6 -8 86 248
use NAND2X1  _12356_
timestamp 0
transform 1 0 10690 0 1 11290
box -6 -8 86 248
use INVX1  _12357_
timestamp 0
transform -1 0 10010 0 1 10330
box -6 -8 66 248
use AOI21X1  _12358_
timestamp 0
transform -1 0 10590 0 1 9850
box -6 -8 106 248
use OAI21X1  _12359_
timestamp 0
transform -1 0 10430 0 1 9850
box -6 -8 106 248
use OAI21X1  _12360_
timestamp 0
transform -1 0 10150 0 1 9850
box -6 -8 106 248
use OR2X2  _12361_
timestamp 0
transform -1 0 9790 0 1 10330
box -6 -8 106 248
use NAND2X1  _12362_
timestamp 0
transform -1 0 9910 0 1 10330
box -6 -8 86 248
use NAND2X1  _12363_
timestamp 0
transform -1 0 9870 0 -1 10810
box -6 -8 86 248
use AOI21X1  _12364_
timestamp 0
transform -1 0 10990 0 -1 9850
box -6 -8 106 248
use AND2X2  _12365_
timestamp 0
transform 1 0 9990 0 1 11290
box -6 -8 106 248
use OAI21X1  _12366_
timestamp 0
transform 1 0 10130 0 1 11290
box -6 -8 106 248
use OAI21X1  _12367_
timestamp 0
transform 1 0 10290 0 1 11290
box -6 -8 106 248
use OAI21X1  _12368_
timestamp 0
transform -1 0 9650 0 1 10810
box -6 -8 106 248
use INVX1  _12369_
timestamp 0
transform -1 0 9990 0 1 9850
box -6 -8 66 248
use OAI21X1  _12370_
timestamp 0
transform 1 0 12710 0 1 9370
box -6 -8 106 248
use OAI21X1  _12371_
timestamp 0
transform 1 0 12050 0 1 9370
box -6 -8 106 248
use OR2X2  _12372_
timestamp 0
transform 1 0 12210 0 1 9370
box -6 -8 106 248
use NAND2X1  _12373_
timestamp 0
transform -1 0 12430 0 1 9370
box -6 -8 86 248
use OR2X2  _12374_
timestamp 0
transform -1 0 10290 0 1 9850
box -6 -8 106 248
use NAND2X1  _12375_
timestamp 0
transform -1 0 10330 0 -1 9850
box -6 -8 86 248
use NAND2X1  _12376_
timestamp 0
transform 1 0 10290 0 -1 10330
box -6 -8 86 248
use INVX1  _12377_
timestamp 0
transform 1 0 9930 0 -1 10810
box -6 -8 66 248
use NOR2X1  _12378_
timestamp 0
transform -1 0 9370 0 1 10810
box -6 -8 86 248
use NAND2X1  _12379_
timestamp 0
transform -1 0 9510 0 1 10810
box -6 -8 86 248
use NAND2X1  _12380_
timestamp 0
transform -1 0 9590 0 -1 11290
box -6 -8 86 248
use OAI22X1  _12381_
timestamp 0
transform -1 0 9470 0 -1 11290
box -6 -8 126 248
use NAND2X1  _12382_
timestamp 0
transform 1 0 10690 0 -1 11290
box -6 -8 86 248
use INVX1  _12383_
timestamp 0
transform 1 0 9690 0 1 10810
box -6 -8 66 248
use NAND2X1  _12384_
timestamp 0
transform 1 0 9810 0 1 10810
box -6 -8 86 248
use OAI21X1  _12385_
timestamp 0
transform 1 0 10050 0 1 10330
box -6 -8 106 248
use INVX1  _12386_
timestamp 0
transform -1 0 9990 0 1 10810
box -6 -8 66 248
use OAI21X1  _12387_
timestamp 0
transform -1 0 9870 0 -1 11290
box -6 -8 106 248
use OAI21X1  _12388_
timestamp 0
transform -1 0 12590 0 -1 9850
box -6 -8 106 248
use NOR2X1  _12389_
timestamp 0
transform 1 0 12510 0 1 9850
box -6 -8 86 248
use NAND2X1  _12390_
timestamp 0
transform 1 0 12210 0 1 9850
box -6 -8 86 248
use OAI21X1  _12391_
timestamp 0
transform -1 0 12450 0 1 9850
box -6 -8 106 248
use NAND2X1  _12392_
timestamp 0
transform -1 0 12170 0 1 9850
box -6 -8 86 248
use NAND2X1  _12393_
timestamp 0
transform 1 0 11030 0 1 9850
box -6 -8 86 248
use OR2X2  _12394_
timestamp 0
transform -1 0 10990 0 1 9850
box -6 -8 106 248
use NAND2X1  _12395_
timestamp 0
transform 1 0 10870 0 -1 10810
box -6 -8 86 248
use INVX1  _12396_
timestamp 0
transform -1 0 10110 0 1 10810
box -6 -8 66 248
use NOR2X1  _12397_
timestamp 0
transform -1 0 10130 0 -1 11290
box -6 -8 86 248
use NAND2X1  _12398_
timestamp 0
transform -1 0 10010 0 -1 11290
box -6 -8 86 248
use NAND2X1  _12399_
timestamp 0
transform -1 0 10250 0 -1 11290
box -6 -8 86 248
use OAI21X1  _12400_
timestamp 0
transform 1 0 10290 0 -1 11290
box -6 -8 106 248
use INVX1  _12401_
timestamp 0
transform 1 0 10410 0 1 10810
box -6 -8 66 248
use NAND2X1  _12402_
timestamp 0
transform 1 0 10750 0 -1 10810
box -6 -8 86 248
use INVX1  _12403_
timestamp 0
transform 1 0 11350 0 -1 9370
box -6 -8 66 248
use NAND2X1  _12404_
timestamp 0
transform -1 0 10630 0 -1 10330
box -6 -8 86 248
use OR2X2  _12405_
timestamp 0
transform -1 0 10510 0 -1 10330
box -6 -8 106 248
use NAND2X1  _12406_
timestamp 0
transform 1 0 10690 0 -1 10330
box -6 -8 86 248
use NOR2X1  _12407_
timestamp 0
transform -1 0 10890 0 -1 10330
box -6 -8 86 248
use INVX1  _12408_
timestamp 0
transform -1 0 10690 0 1 10330
box -6 -8 66 248
use NAND2X1  _12409_
timestamp 0
transform -1 0 11010 0 -1 10330
box -6 -8 86 248
use NAND2X1  _12410_
timestamp 0
transform -1 0 10570 0 1 10330
box -6 -8 86 248
use OR2X2  _12411_
timestamp 0
transform 1 0 10610 0 -1 10810
box -6 -8 106 248
use AOI21X1  _12412_
timestamp 0
transform -1 0 10570 0 -1 10810
box -6 -8 106 248
use AOI22X1  _12413_
timestamp 0
transform 1 0 10530 0 1 10810
box -6 -8 126 248
use NAND2X1  _12414_
timestamp 0
transform 1 0 11150 0 -1 10810
box -6 -8 86 248
use NOR2X1  _12415_
timestamp 0
transform 1 0 11910 0 -1 9850
box -6 -8 86 248
use INVX1  _12416_
timestamp 0
transform -1 0 11850 0 -1 9850
box -6 -8 66 248
use NAND3X1  _12417_
timestamp 0
transform -1 0 11770 0 1 9850
box -6 -8 106 248
use INVX1  _12418_
timestamp 0
transform 1 0 11650 0 1 10330
box -6 -8 66 248
use AOI21X1  _12419_
timestamp 0
transform 1 0 11810 0 1 9850
box -6 -8 106 248
use NOR2X1  _12420_
timestamp 0
transform -1 0 11850 0 -1 10330
box -6 -8 86 248
use OAI21X1  _12421_
timestamp 0
transform -1 0 10430 0 1 10330
box -6 -8 106 248
use NOR2X1  _12422_
timestamp 0
transform -1 0 10430 0 -1 10810
box -6 -8 86 248
use AOI21X1  _12423_
timestamp 0
transform 1 0 10190 0 1 10330
box -6 -8 106 248
use NAND3X1  _12424_
timestamp 0
transform 1 0 10030 0 -1 10810
box -6 -8 106 248
use OAI21X1  _12425_
timestamp 0
transform 1 0 10190 0 -1 10810
box -6 -8 106 248
use NOR2X1  _12426_
timestamp 0
transform 1 0 11270 0 -1 10810
box -6 -8 86 248
use NAND2X1  _12427_
timestamp 0
transform -1 0 11190 0 1 10330
box -6 -8 86 248
use NAND2X1  _12428_
timestamp 0
transform -1 0 11050 0 1 10330
box -6 -8 86 248
use OAI21X1  _12429_
timestamp 0
transform 1 0 11010 0 -1 10810
box -6 -8 106 248
use AOI21X1  _12430_
timestamp 0
transform -1 0 11750 0 -1 10810
box -6 -8 106 248
use OR2X2  _12431_
timestamp 0
transform -1 0 11850 0 1 10330
box -6 -8 106 248
use NAND2X1  _12432_
timestamp 0
transform -1 0 11710 0 -1 10330
box -6 -8 86 248
use NAND2X1  _12433_
timestamp 0
transform -1 0 11310 0 1 10330
box -6 -8 86 248
use AND2X2  _12434_
timestamp 0
transform -1 0 11350 0 1 10810
box -6 -8 106 248
use OAI21X1  _12435_
timestamp 0
transform 1 0 11390 0 1 10810
box -6 -8 106 248
use OAI22X1  _12436_
timestamp 0
transform -1 0 11470 0 -1 11290
box -6 -8 126 248
use NAND2X1  _12437_
timestamp 0
transform -1 0 11890 0 -1 10810
box -6 -8 86 248
use OAI21X1  _12438_
timestamp 0
transform 1 0 11510 0 1 10330
box -6 -8 106 248
use NAND3X1  _12439_
timestamp 0
transform -1 0 11470 0 1 10330
box -6 -8 106 248
use INVX1  _12440_
timestamp 0
transform -1 0 11450 0 -1 10810
box -6 -8 66 248
use AOI21X1  _12441_
timestamp 0
transform 1 0 11510 0 -1 10810
box -6 -8 106 248
use INVX1  _12442_
timestamp 0
transform -1 0 12210 0 1 10330
box -6 -8 66 248
use NAND2X1  _12443_
timestamp 0
transform 1 0 12210 0 -1 10330
box -6 -8 86 248
use NAND2X1  _12444_
timestamp 0
transform -1 0 12110 0 1 10330
box -6 -8 86 248
use NAND2X1  _12445_
timestamp 0
transform 1 0 12390 0 -1 10810
box -6 -8 86 248
use AND2X2  _12446_
timestamp 0
transform -1 0 12210 0 -1 10810
box -6 -8 106 248
use OAI21X1  _12447_
timestamp 0
transform -1 0 12130 0 1 10810
box -6 -8 106 248
use OAI21X1  _12448_
timestamp 0
transform -1 0 12050 0 -1 10810
box -6 -8 106 248
use NAND2X1  _12449_
timestamp 0
transform 1 0 12210 0 -1 11290
box -6 -8 86 248
use OAI21X1  _12450_
timestamp 0
transform 1 0 12250 0 -1 10810
box -6 -8 106 248
use OAI21X1  _12451_
timestamp 0
transform 1 0 12070 0 -1 11290
box -6 -8 106 248
use NAND2X1  _12452_
timestamp 0
transform 1 0 11790 0 -1 7930
box -6 -8 86 248
use NAND2X1  _12453_
timestamp 0
transform -1 0 11790 0 1 7930
box -6 -8 86 248
use NOR2X1  _12454_
timestamp 0
transform 1 0 11830 0 1 7930
box -6 -8 86 248
use NAND2X1  _12455_
timestamp 0
transform -1 0 13950 0 1 9850
box -6 -8 86 248
use OAI21X1  _12456_
timestamp 0
transform -1 0 14110 0 1 9850
box -6 -8 106 248
use NAND2X1  _12457_
timestamp 0
transform -1 0 14030 0 1 8890
box -6 -8 86 248
use OAI21X1  _12458_
timestamp 0
transform -1 0 14190 0 1 8890
box -6 -8 106 248
use INVX1  _12459_
timestamp 0
transform 1 0 14050 0 -1 10330
box -6 -8 66 248
use OR2X2  _12460_
timestamp 0
transform -1 0 11830 0 -1 8410
box -6 -8 106 248
use OAI21X1  _12461_
timestamp 0
transform 1 0 14010 0 -1 9370
box -6 -8 106 248
use OAI21X1  _12462_
timestamp 0
transform 1 0 13870 0 -1 9370
box -6 -8 106 248
use INVX1  _12463_
timestamp 0
transform 1 0 14170 0 -1 9370
box -6 -8 66 248
use OAI21X1  _12464_
timestamp 0
transform 1 0 13730 0 -1 9370
box -6 -8 106 248
use OAI21X1  _12465_
timestamp 0
transform -1 0 13670 0 1 9370
box -6 -8 106 248
use NAND2X1  _12466_
timestamp 0
transform 1 0 12310 0 1 8410
box -6 -8 86 248
use NAND2X1  _12467_
timestamp 0
transform -1 0 14890 0 -1 9370
box -6 -8 86 248
use OAI21X1  _12468_
timestamp 0
transform 1 0 14290 0 -1 9370
box -6 -8 106 248
use NAND2X1  _12469_
timestamp 0
transform 1 0 14350 0 1 9370
box -6 -8 86 248
use OAI21X1  _12470_
timestamp 0
transform 1 0 13970 0 1 9370
box -6 -8 106 248
use AND2X2  _12471_
timestamp 0
transform 1 0 12190 0 -1 9850
box -6 -8 106 248
use NAND2X1  _12472_
timestamp 0
transform 1 0 16450 0 -1 12250
box -6 -8 86 248
use OAI21X1  _12473_
timestamp 0
transform -1 0 16670 0 -1 12250
box -6 -8 106 248
use NAND2X1  _12474_
timestamp 0
transform 1 0 15190 0 -1 12250
box -6 -8 86 248
use OAI21X1  _12475_
timestamp 0
transform -1 0 15670 0 -1 12250
box -6 -8 106 248
use OAI21X1  _12476_
timestamp 0
transform 1 0 13570 0 1 9850
box -6 -8 106 248
use OAI21X1  _12477_
timestamp 0
transform -1 0 13830 0 1 9850
box -6 -8 106 248
use OAI21X1  _12478_
timestamp 0
transform 1 0 13630 0 -1 9850
box -6 -8 106 248
use OAI21X1  _12479_
timestamp 0
transform -1 0 13890 0 -1 9850
box -6 -8 106 248
use NAND2X1  _12480_
timestamp 0
transform -1 0 12970 0 -1 10330
box -6 -8 86 248
use OAI21X1  _12481_
timestamp 0
transform 1 0 13010 0 -1 10330
box -6 -8 106 248
use NAND2X1  _12482_
timestamp 0
transform 1 0 13690 0 -1 10330
box -6 -8 86 248
use OAI21X1  _12483_
timestamp 0
transform 1 0 13530 0 -1 10330
box -6 -8 106 248
use NAND2X1  _12484_
timestamp 0
transform -1 0 14110 0 -1 8410
box -6 -8 86 248
use OAI21X1  _12485_
timestamp 0
transform -1 0 14250 0 -1 8410
box -6 -8 106 248
use NAND2X1  _12486_
timestamp 0
transform 1 0 14170 0 -1 8890
box -6 -8 86 248
use OAI21X1  _12487_
timestamp 0
transform -1 0 14410 0 -1 8890
box -6 -8 106 248
use INVX1  _12488_
timestamp 0
transform -1 0 13970 0 -1 8410
box -6 -8 66 248
use OAI21X1  _12489_
timestamp 0
transform -1 0 13870 0 -1 8410
box -6 -8 106 248
use OAI21X1  _12490_
timestamp 0
transform 1 0 13610 0 -1 8410
box -6 -8 106 248
use INVX1  _12491_
timestamp 0
transform -1 0 14130 0 -1 8890
box -6 -8 66 248
use OAI21X1  _12492_
timestamp 0
transform 1 0 13410 0 1 7930
box -6 -8 106 248
use OAI21X1  _12493_
timestamp 0
transform -1 0 13650 0 1 7930
box -6 -8 106 248
use NAND2X1  _12494_
timestamp 0
transform -1 0 14570 0 1 8410
box -6 -8 86 248
use OAI21X1  _12495_
timestamp 0
transform 1 0 14090 0 1 8410
box -6 -8 106 248
use NAND2X1  _12496_
timestamp 0
transform -1 0 14850 0 1 8410
box -6 -8 86 248
use OAI21X1  _12497_
timestamp 0
transform 1 0 14610 0 1 8410
box -6 -8 106 248
use NAND2X1  _12498_
timestamp 0
transform 1 0 16370 0 -1 8890
box -6 -8 86 248
use OAI21X1  _12499_
timestamp 0
transform -1 0 16730 0 -1 8890
box -6 -8 106 248
use NAND2X1  _12500_
timestamp 0
transform 1 0 16530 0 1 8890
box -6 -8 86 248
use OAI21X1  _12501_
timestamp 0
transform -1 0 16770 0 1 8890
box -6 -8 106 248
use OAI21X1  _12502_
timestamp 0
transform -1 0 13430 0 -1 8890
box -6 -8 106 248
use OAI21X1  _12503_
timestamp 0
transform -1 0 13590 0 -1 8890
box -6 -8 106 248
use OAI21X1  _12504_
timestamp 0
transform 1 0 13570 0 1 8410
box -6 -8 106 248
use OAI21X1  _12505_
timestamp 0
transform -1 0 13810 0 1 8410
box -6 -8 106 248
use NAND2X1  _12506_
timestamp 0
transform -1 0 12190 0 -1 8890
box -6 -8 86 248
use OAI21X1  _12507_
timestamp 0
transform -1 0 12330 0 -1 8890
box -6 -8 106 248
use NAND2X1  _12508_
timestamp 0
transform -1 0 11890 0 1 8890
box -6 -8 86 248
use OAI21X1  _12509_
timestamp 0
transform -1 0 12030 0 1 8890
box -6 -8 106 248
use NAND2X1  _12510_
timestamp 0
transform 1 0 12490 0 -1 10330
box -6 -8 86 248
use OAI21X1  _12511_
timestamp 0
transform 1 0 12330 0 -1 10330
box -6 -8 106 248
use NAND2X1  _12512_
timestamp 0
transform 1 0 11890 0 1 8410
box -6 -8 86 248
use OAI21X1  _12513_
timestamp 0
transform -1 0 12070 0 1 7930
box -6 -8 106 248
use INVX1  _12514_
timestamp 0
transform 1 0 12070 0 -1 9370
box -6 -8 66 248
use OAI21X1  _12515_
timestamp 0
transform -1 0 12430 0 -1 9370
box -6 -8 106 248
use OAI21X1  _12516_
timestamp 0
transform 1 0 12170 0 -1 9370
box -6 -8 106 248
use INVX1  _12517_
timestamp 0
transform 1 0 11690 0 1 8890
box -6 -8 66 248
use OAI21X1  _12518_
timestamp 0
transform -1 0 12270 0 1 8410
box -6 -8 106 248
use OAI21X1  _12519_
timestamp 0
transform 1 0 12010 0 1 8410
box -6 -8 106 248
use NAND2X1  _12520_
timestamp 0
transform 1 0 11030 0 -1 8890
box -6 -8 86 248
use OAI21X1  _12521_
timestamp 0
transform -1 0 11250 0 -1 8890
box -6 -8 106 248
use NAND2X1  _12522_
timestamp 0
transform 1 0 11430 0 1 8890
box -6 -8 86 248
use OAI21X1  _12523_
timestamp 0
transform -1 0 11650 0 1 8890
box -6 -8 106 248
use NAND2X1  _12524_
timestamp 0
transform -1 0 9490 0 1 10330
box -6 -8 86 248
use OAI21X1  _12525_
timestamp 0
transform -1 0 9650 0 1 10330
box -6 -8 106 248
use NAND2X1  _12526_
timestamp 0
transform -1 0 9730 0 1 9850
box -6 -8 86 248
use OAI21X1  _12527_
timestamp 0
transform -1 0 9890 0 1 9850
box -6 -8 106 248
use OAI21X1  _12528_
timestamp 0
transform 1 0 11370 0 1 8410
box -6 -8 106 248
use OAI21X1  _12529_
timestamp 0
transform -1 0 11850 0 1 8410
box -6 -8 106 248
use OAI21X1  _12530_
timestamp 0
transform -1 0 11710 0 1 9370
box -6 -8 106 248
use OAI21X1  _12531_
timestamp 0
transform -1 0 11850 0 1 9370
box -6 -8 106 248
use NAND2X1  _12532_
timestamp 0
transform 1 0 11210 0 -1 9370
box -6 -8 86 248
use OAI21X1  _12533_
timestamp 0
transform 1 0 11050 0 -1 9370
box -6 -8 106 248
use NAND2X1  _12534_
timestamp 0
transform 1 0 10830 0 -1 9370
box -6 -8 86 248
use OAI21X1  _12535_
timestamp 0
transform -1 0 10770 0 -1 9370
box -6 -8 106 248
use DFFPOSX1  _12536_
timestamp 0
transform 1 0 12210 0 1 7930
box -6 -8 246 248
use DFFPOSX1  _12537_
timestamp 0
transform 1 0 12150 0 -1 8410
box -6 -8 246 248
use DFFPOSX1  _12538_
timestamp 0
transform 1 0 8970 0 1 11290
box -6 -8 246 248
use DFFPOSX1  _12539_
timestamp 0
transform 1 0 12230 0 -1 7930
box -6 -8 246 248
use DFFPOSX1  _12540_
timestamp 0
transform 1 0 12490 0 1 7450
box -6 -8 246 248
use DFFPOSX1  _12541_
timestamp 0
transform -1 0 13870 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _12542_
timestamp 0
transform 1 0 12190 0 -1 7450
box -6 -8 246 248
use DFFPOSX1  _12543_
timestamp 0
transform -1 0 14390 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _12544_
timestamp 0
transform 1 0 12590 0 1 6970
box -6 -8 246 248
use DFFPOSX1  _12545_
timestamp 0
transform -1 0 14050 0 1 6970
box -6 -8 246 248
use DFFPOSX1  _12546_
timestamp 0
transform -1 0 13810 0 1 6970
box -6 -8 246 248
use DFFPOSX1  _12547_
timestamp 0
transform -1 0 14090 0 1 7450
box -6 -8 246 248
use DFFPOSX1  _12548_
timestamp 0
transform -1 0 13350 0 -1 7930
box -6 -8 246 248
use DFFPOSX1  _12549_
timestamp 0
transform 1 0 12590 0 -1 10810
box -6 -8 246 248
use DFFPOSX1  _12550_
timestamp 0
transform 1 0 12290 0 1 10810
box -6 -8 246 248
use DFFPOSX1  _12551_
timestamp 0
transform -1 0 13670 0 -1 10810
box -6 -8 246 248
use DFFPOSX1  _12552_
timestamp 0
transform -1 0 14770 0 1 11770
box -6 -8 246 248
use DFFPOSX1  _12553_
timestamp 0
transform -1 0 13770 0 1 11770
box -6 -8 246 248
use DFFPOSX1  _12554_
timestamp 0
transform -1 0 13710 0 -1 11770
box -6 -8 246 248
use DFFPOSX1  _12555_
timestamp 0
transform -1 0 12970 0 -1 11770
box -6 -8 246 248
use DFFPOSX1  _12556_
timestamp 0
transform -1 0 13950 0 -1 11770
box -6 -8 246 248
use DFFPOSX1  _12557_
timestamp 0
transform -1 0 13530 0 1 11290
box -6 -8 246 248
use DFFPOSX1  _12558_
timestamp 0
transform -1 0 13810 0 1 10810
box -6 -8 246 248
use DFFPOSX1  _12559_
timestamp 0
transform -1 0 13370 0 -1 11290
box -6 -8 246 248
use DFFPOSX1  _12560_
timestamp 0
transform -1 0 13450 0 1 10810
box -6 -8 246 248
use DFFPOSX1  _12561_
timestamp 0
transform 1 0 11250 0 1 9850
box -6 -8 246 248
use DFFPOSX1  _12562_
timestamp 0
transform -1 0 11650 0 -1 9370
box -6 -8 246 248
use DFFPOSX1  _12563_
timestamp 0
transform 1 0 9630 0 -1 8890
box -6 -8 246 248
use DFFPOSX1  _12564_
timestamp 0
transform 1 0 10690 0 1 10330
box -6 -8 246 248
use DFFPOSX1  _12565_
timestamp 0
transform 1 0 10390 0 1 11290
box -6 -8 246 248
use DFFPOSX1  _12566_
timestamp 0
transform 1 0 9070 0 -1 11290
box -6 -8 246 248
use DFFPOSX1  _12567_
timestamp 0
transform 1 0 10390 0 -1 11290
box -6 -8 246 248
use DFFPOSX1  _12568_
timestamp 0
transform 1 0 10110 0 1 10810
box -6 -8 246 248
use DFFPOSX1  _12569_
timestamp 0
transform 1 0 10650 0 1 10810
box -6 -8 246 248
use DFFPOSX1  _12570_
timestamp 0
transform 1 0 11310 0 1 11290
box -6 -8 246 248
use DFFPOSX1  _12571_
timestamp 0
transform -1 0 11850 0 1 10810
box -6 -8 246 248
use DFFPOSX1  _12572_
timestamp 0
transform -1 0 12170 0 1 11290
box -6 -8 246 248
use DFFPOSX1  _12573_
timestamp 0
transform 1 0 14110 0 1 9850
box -6 -8 246 248
use DFFPOSX1  _12574_
timestamp 0
transform 1 0 14290 0 1 8890
box -6 -8 246 248
use DFFPOSX1  _12575_
timestamp 0
transform 1 0 13670 0 1 9370
box -6 -8 246 248
use DFFPOSX1  _12576_
timestamp 0
transform 1 0 13270 0 1 9370
box -6 -8 246 248
use DFFPOSX1  _12577_
timestamp 0
transform 1 0 14890 0 -1 9370
box -6 -8 246 248
use DFFPOSX1  _12578_
timestamp 0
transform 1 0 14070 0 1 9370
box -6 -8 246 248
use DFFPOSX1  _12579_
timestamp 0
transform -1 0 16910 0 -1 12250
box -6 -8 246 248
use DFFPOSX1  _12580_
timestamp 0
transform -1 0 15910 0 -1 12250
box -6 -8 246 248
use DFFPOSX1  _12581_
timestamp 0
transform 1 0 13770 0 -1 10330
box -6 -8 246 248
use DFFPOSX1  _12582_
timestamp 0
transform 1 0 13890 0 -1 9850
box -6 -8 246 248
use DFFPOSX1  _12583_
timestamp 0
transform 1 0 12450 0 1 10330
box -6 -8 246 248
use DFFPOSX1  _12584_
timestamp 0
transform -1 0 13470 0 1 10330
box -6 -8 246 248
use DFFPOSX1  _12585_
timestamp 0
transform 1 0 14250 0 -1 8410
box -6 -8 246 248
use DFFPOSX1  _12586_
timestamp 0
transform 1 0 14410 0 -1 8890
box -6 -8 246 248
use DFFPOSX1  _12587_
timestamp 0
transform 1 0 13330 0 -1 8410
box -6 -8 246 248
use DFFPOSX1  _12588_
timestamp 0
transform 1 0 13650 0 1 7930
box -6 -8 246 248
use DFFPOSX1  _12589_
timestamp 0
transform 1 0 14190 0 1 8410
box -6 -8 246 248
use DFFPOSX1  _12590_
timestamp 0
transform 1 0 14850 0 1 8410
box -6 -8 246 248
use DFFPOSX1  _12591_
timestamp 0
transform 1 0 16730 0 1 8410
box -6 -8 246 248
use DFFPOSX1  _12592_
timestamp 0
transform 1 0 16770 0 1 8890
box -6 -8 246 248
use DFFPOSX1  _12593_
timestamp 0
transform 1 0 12750 0 -1 8890
box -6 -8 246 248
use DFFPOSX1  _12594_
timestamp 0
transform 1 0 13810 0 1 8410
box -6 -8 246 248
use DFFPOSX1  _12595_
timestamp 0
transform 1 0 12370 0 1 8890
box -6 -8 246 248
use DFFPOSX1  _12596_
timestamp 0
transform 1 0 12030 0 1 8890
box -6 -8 246 248
use DFFPOSX1  _12597_
timestamp 0
transform -1 0 12450 0 1 10330
box -6 -8 246 248
use DFFPOSX1  _12598_
timestamp 0
transform 1 0 11870 0 -1 7930
box -6 -8 246 248
use DFFPOSX1  _12599_
timestamp 0
transform -1 0 12030 0 -1 9370
box -6 -8 246 248
use DFFPOSX1  _12600_
timestamp 0
transform 1 0 11430 0 -1 8410
box -6 -8 246 248
use DFFPOSX1  _12601_
timestamp 0
transform 1 0 10730 0 -1 8890
box -6 -8 246 248
use DFFPOSX1  _12602_
timestamp 0
transform -1 0 11490 0 -1 8890
box -6 -8 246 248
use DFFPOSX1  _12603_
timestamp 0
transform -1 0 10250 0 -1 10330
box -6 -8 246 248
use DFFPOSX1  _12604_
timestamp 0
transform -1 0 10190 0 -1 9850
box -6 -8 246 248
use DFFPOSX1  _12605_
timestamp 0
transform -1 0 11710 0 1 8410
box -6 -8 246 248
use DFFPOSX1  _12606_
timestamp 0
transform 1 0 11310 0 1 9370
box -6 -8 246 248
use DFFPOSX1  _12607_
timestamp 0
transform 1 0 10430 0 1 9370
box -6 -8 246 248
use DFFPOSX1  _12608_
timestamp 0
transform -1 0 10630 0 -1 9370
box -6 -8 246 248
use DFFPOSX1  _12609_
timestamp 0
transform 1 0 9250 0 -1 10330
box -6 -8 246 248
use DFFPOSX1  _12610_
timestamp 0
transform 1 0 10710 0 -1 8410
box -6 -8 246 248
use DFFPOSX1  _12611_
timestamp 0
transform 1 0 10950 0 -1 8410
box -6 -8 246 248
use DFFPOSX1  _12612_
timestamp 0
transform 1 0 11070 0 1 11290
box -6 -8 246 248
use DFFPOSX1  _12613_
timestamp 0
transform 1 0 11690 0 1 11290
box -6 -8 246 248
use DFFPOSX1  _12614_
timestamp 0
transform -1 0 12010 0 1 7450
box -6 -8 246 248
use DFFPOSX1  _12615_
timestamp 0
transform -1 0 11750 0 -1 7930
box -6 -8 246 248
use INVX2  _12616_
timestamp 0
transform 1 0 11290 0 1 13690
box -6 -8 66 248
use NOR2X1  _12617_
timestamp 0
transform -1 0 11490 0 1 13690
box -6 -8 86 248
use INVX2  _12618_
timestamp 0
transform 1 0 12370 0 -1 14170
box -6 -8 66 248
use INVX4  _12619_
timestamp 0
transform 1 0 11530 0 1 16090
box -6 -8 86 248
use NOR2X1  _12620_
timestamp 0
transform -1 0 11170 0 1 16090
box -6 -8 86 248
use INVX2  _12621_
timestamp 0
transform -1 0 10910 0 1 16090
box -6 -8 66 248
use AND2X2  _12622_
timestamp 0
transform 1 0 10950 0 1 16090
box -6 -8 106 248
use NOR2X1  _12623_
timestamp 0
transform -1 0 11130 0 1 13690
box -6 -8 86 248
use INVX1  _12624_
timestamp 0
transform -1 0 11610 0 1 13690
box -6 -8 66 248
use OAI21X1  _12625_
timestamp 0
transform -1 0 11810 0 1 14170
box -6 -8 106 248
use AOI21X1  _12626_
timestamp 0
transform -1 0 11670 0 1 14170
box -6 -8 106 248
use INVX1  _12627_
timestamp 0
transform -1 0 10670 0 1 11770
box -6 -8 66 248
use NAND2X1  _12628_
timestamp 0
transform -1 0 11590 0 -1 14170
box -6 -8 86 248
use OAI21X1  _12629_
timestamp 0
transform 1 0 11370 0 -1 14170
box -6 -8 106 248
use OAI21X1  _12630_
timestamp 0
transform -1 0 11310 0 -1 14170
box -6 -8 106 248
use AOI22X1  _12631_
timestamp 0
transform 1 0 11230 0 -1 13690
box -6 -8 126 248
use NAND2X1  _12632_
timestamp 0
transform 1 0 11170 0 1 13690
box -6 -8 86 248
use INVX1  _12633_
timestamp 0
transform 1 0 11670 0 1 16090
box -6 -8 66 248
use OAI21X1  _12634_
timestamp 0
transform -1 0 11250 0 -1 16090
box -6 -8 106 248
use AOI21X1  _12635_
timestamp 0
transform -1 0 11390 0 -1 16090
box -6 -8 106 248
use INVX1  _12636_
timestamp 0
transform -1 0 11710 0 1 15130
box -6 -8 66 248
use NAND2X1  _12637_
timestamp 0
transform -1 0 11890 0 -1 15610
box -6 -8 86 248
use OAI21X1  _12638_
timestamp 0
transform 1 0 11670 0 -1 15610
box -6 -8 106 248
use OAI21X1  _12639_
timestamp 0
transform -1 0 11350 0 1 15610
box -6 -8 106 248
use AOI22X1  _12640_
timestamp 0
transform -1 0 11790 0 -1 14650
box -6 -8 126 248
use NAND2X1  _12641_
timestamp 0
transform -1 0 11390 0 -1 15130
box -6 -8 86 248
use INVX1  _12642_
timestamp 0
transform 1 0 10970 0 1 16570
box -6 -8 66 248
use OAI21X1  _12643_
timestamp 0
transform -1 0 11430 0 -1 16570
box -6 -8 106 248
use AOI21X1  _12644_
timestamp 0
transform -1 0 11110 0 -1 16570
box -6 -8 106 248
use INVX1  _12645_
timestamp 0
transform -1 0 11230 0 -1 15610
box -6 -8 66 248
use NAND2X1  _12646_
timestamp 0
transform -1 0 11610 0 1 15610
box -6 -8 86 248
use OAI21X1  _12647_
timestamp 0
transform 1 0 11390 0 1 15610
box -6 -8 106 248
use OAI21X1  _12648_
timestamp 0
transform 1 0 11110 0 1 15610
box -6 -8 106 248
use AOI22X1  _12649_
timestamp 0
transform 1 0 11430 0 1 14650
box -6 -8 126 248
use NAND2X1  _12650_
timestamp 0
transform -1 0 11030 0 -1 15130
box -6 -8 86 248
use INVX1  _12651_
timestamp 0
transform -1 0 10510 0 -1 17050
box -6 -8 66 248
use OAI21X1  _12652_
timestamp 0
transform 1 0 11170 0 -1 16570
box -6 -8 106 248
use AOI21X1  _12653_
timestamp 0
transform 1 0 11210 0 1 16090
box -6 -8 106 248
use INVX1  _12654_
timestamp 0
transform -1 0 11550 0 1 16570
box -6 -8 66 248
use NAND2X1  _12655_
timestamp 0
transform 1 0 11230 0 1 16570
box -6 -8 86 248
use OAI21X1  _12656_
timestamp 0
transform -1 0 11450 0 1 16570
box -6 -8 106 248
use OAI21X1  _12657_
timestamp 0
transform 1 0 11370 0 1 16090
box -6 -8 106 248
use AOI22X1  _12658_
timestamp 0
transform 1 0 12110 0 1 14650
box -6 -8 126 248
use NAND2X1  _12659_
timestamp 0
transform -1 0 11470 0 1 15130
box -6 -8 86 248
use INVX1  _12660_
timestamp 0
transform -1 0 12590 0 1 14170
box -6 -8 66 248
use NOR2X1  _12661_
timestamp 0
transform 1 0 12150 0 1 16570
box -6 -8 86 248
use OAI21X1  _12662_
timestamp 0
transform -1 0 12490 0 -1 16570
box -6 -8 106 248
use AOI22X1  _12663_
timestamp 0
transform -1 0 12110 0 1 16570
box -6 -8 126 248
use OAI21X1  _12664_
timestamp 0
transform -1 0 12210 0 -1 16570
box -6 -8 106 248
use AOI22X1  _12665_
timestamp 0
transform 1 0 11970 0 -1 14650
box -6 -8 126 248
use OAI21X1  _12666_
timestamp 0
transform -1 0 11930 0 -1 14650
box -6 -8 106 248
use INVX1  _12667_
timestamp 0
transform -1 0 12090 0 -1 14170
box -6 -8 66 248
use INVX1  _12668_
timestamp 0
transform -1 0 13390 0 -1 13210
box -6 -8 66 248
use INVX8  _12669_
timestamp 0
transform -1 0 17150 0 1 14170
box -6 -8 126 248
use INVX8  _12670_
timestamp 0
transform 1 0 16050 0 1 12730
box -6 -8 126 248
use INVX1  _12671_
timestamp 0
transform 1 0 16730 0 -1 13690
box -6 -8 66 248
use NAND2X1  _12672_
timestamp 0
transform -1 0 16630 0 1 13210
box -6 -8 86 248
use OAI21X1  _12673_
timestamp 0
transform -1 0 16770 0 1 13210
box -6 -8 106 248
use INVX1  _12674_
timestamp 0
transform 1 0 16910 0 1 14170
box -6 -8 66 248
use NAND2X1  _12675_
timestamp 0
transform 1 0 17090 0 -1 13210
box -6 -8 86 248
use OAI21X1  _12676_
timestamp 0
transform 1 0 16950 0 -1 13210
box -6 -8 106 248
use MUX2X1  _12677_
timestamp 0
transform -1 0 16710 0 -1 13210
box -6 -8 126 248
use INVX1  _12678_
timestamp 0
transform 1 0 16450 0 -1 12730
box -6 -8 66 248
use NAND2X1  _12679_
timestamp 0
transform -1 0 16270 0 -1 12730
box -6 -8 86 248
use OAI21X1  _12680_
timestamp 0
transform -1 0 16410 0 -1 12730
box -6 -8 106 248
use INVX1  _12681_
timestamp 0
transform 1 0 15970 0 1 12250
box -6 -8 66 248
use NAND2X1  _12682_
timestamp 0
transform 1 0 16710 0 -1 12730
box -6 -8 86 248
use OAI21X1  _12683_
timestamp 0
transform 1 0 16570 0 -1 12730
box -6 -8 106 248
use MUX2X1  _12684_
timestamp 0
transform 1 0 16370 0 1 12730
box -6 -8 126 248
use MUX2X1  _12685_
timestamp 0
transform -1 0 16370 0 -1 13210
box -6 -8 126 248
use NOR2X1  _12686_
timestamp 0
transform -1 0 13210 0 1 13210
box -6 -8 86 248
use NAND2X1  _12687_
timestamp 0
transform -1 0 13330 0 1 13210
box -6 -8 86 248
use INVX1  _12688_
timestamp 0
transform -1 0 12730 0 1 13690
box -6 -8 66 248
use NAND2X1  _12689_
timestamp 0
transform -1 0 14990 0 1 12250
box -6 -8 86 248
use OAI21X1  _12690_
timestamp 0
transform -1 0 12870 0 1 16570
box -6 -8 106 248
use INVX2  _12691_
timestamp 0
transform 1 0 12930 0 1 16570
box -6 -8 66 248
use OAI21X1  _12692_
timestamp 0
transform -1 0 12610 0 1 13690
box -6 -8 106 248
use OAI21X1  _12693_
timestamp 0
transform 1 0 12090 0 1 13690
box -6 -8 106 248
use INVX8  _12694_
timestamp 0
transform -1 0 11690 0 -1 15130
box -6 -8 126 248
use NAND2X1  _12695_
timestamp 0
transform 1 0 11390 0 -1 14650
box -6 -8 86 248
use NOR2X1  _12696_
timestamp 0
transform -1 0 12950 0 1 14170
box -6 -8 86 248
use MUX2X1  _12697_
timestamp 0
transform -1 0 16170 0 1 13210
box -6 -8 126 248
use MUX2X1  _12698_
timestamp 0
transform -1 0 16550 0 -1 13210
box -6 -8 126 248
use MUX2X1  _12699_
timestamp 0
transform -1 0 16010 0 1 13210
box -6 -8 126 248
use INVX2  _12700_
timestamp 0
transform 1 0 16210 0 -1 12250
box -6 -8 66 248
use NAND2X1  _12701_
timestamp 0
transform 1 0 16050 0 -1 12730
box -6 -8 86 248
use AOI21X1  _12702_
timestamp 0
transform -1 0 16010 0 -1 12730
box -6 -8 106 248
use NAND3X1  _12703_
timestamp 0
transform -1 0 15890 0 1 12730
box -6 -8 106 248
use NAND3X1  _12704_
timestamp 0
transform -1 0 16630 0 1 12730
box -6 -8 106 248
use NAND3X1  _12705_
timestamp 0
transform -1 0 16330 0 1 12730
box -6 -8 106 248
use OAI22X1  _12706_
timestamp 0
transform -1 0 15750 0 1 12730
box -6 -8 126 248
use INVX1  _12707_
timestamp 0
transform 1 0 14510 0 -1 12730
box -6 -8 66 248
use INVX8  _12708_
timestamp 0
transform 1 0 14470 0 1 14650
box -6 -8 126 248
use INVX1  _12709_
timestamp 0
transform 1 0 16390 0 1 15610
box -6 -8 66 248
use NAND2X1  _12710_
timestamp 0
transform 1 0 15790 0 1 15130
box -6 -8 86 248
use OAI21X1  _12711_
timestamp 0
transform 1 0 15910 0 1 15130
box -6 -8 106 248
use INVX1  _12712_
timestamp 0
transform -1 0 16750 0 1 12730
box -6 -8 66 248
use NAND2X1  _12713_
timestamp 0
transform 1 0 16830 0 1 13690
box -6 -8 86 248
use OAI21X1  _12714_
timestamp 0
transform 1 0 16690 0 1 13690
box -6 -8 106 248
use MUX2X1  _12715_
timestamp 0
transform 1 0 16330 0 1 13690
box -6 -8 126 248
use INVX1  _12716_
timestamp 0
transform 1 0 17050 0 -1 250
box -6 -8 66 248
use NAND2X1  _12717_
timestamp 0
transform 1 0 17110 0 1 13690
box -6 -8 86 248
use OAI21X1  _12718_
timestamp 0
transform 1 0 16950 0 1 13690
box -6 -8 106 248
use INVX1  _12719_
timestamp 0
transform 1 0 16730 0 1 12250
box -6 -8 66 248
use NAND2X1  _12720_
timestamp 0
transform 1 0 16810 0 -1 250
box -6 -8 86 248
use OAI21X1  _12721_
timestamp 0
transform 1 0 17010 0 1 16570
box -6 -8 106 248
use MUX2X1  _12722_
timestamp 0
transform 1 0 16970 0 -1 13690
box -6 -8 126 248
use MUX2X1  _12723_
timestamp 0
transform 1 0 16550 0 -1 13690
box -6 -8 126 248
use NAND3X1  _12724_
timestamp 0
transform -1 0 14550 0 1 13210
box -6 -8 106 248
use MUX2X1  _12725_
timestamp 0
transform -1 0 15890 0 1 13690
box -6 -8 126 248
use MUX2X1  _12726_
timestamp 0
transform -1 0 17110 0 1 13210
box -6 -8 126 248
use MUX2X1  _12727_
timestamp 0
transform 1 0 16390 0 1 13210
box -6 -8 126 248
use MUX2X1  _12728_
timestamp 0
transform -1 0 16610 0 -1 250
box -6 -8 126 248
use MUX2X1  _12729_
timestamp 0
transform 1 0 16770 0 -1 13210
box -6 -8 126 248
use MUX2X1  _12730_
timestamp 0
transform -1 0 16930 0 1 13210
box -6 -8 126 248
use MUX2X1  _12731_
timestamp 0
transform -1 0 16350 0 1 13210
box -6 -8 126 248
use OAI21X1  _12732_
timestamp 0
transform 1 0 14130 0 -1 13210
box -6 -8 106 248
use AOI21X1  _12733_
timestamp 0
transform -1 0 14030 0 1 13210
box -6 -8 106 248
use INVX1  _12734_
timestamp 0
transform -1 0 13870 0 1 13210
box -6 -8 66 248
use NAND3X1  _12735_
timestamp 0
transform -1 0 14170 0 1 13210
box -6 -8 106 248
use AND2X2  _12736_
timestamp 0
transform -1 0 13770 0 1 13210
box -6 -8 106 248
use OAI21X1  _12737_
timestamp 0
transform -1 0 13670 0 -1 13210
box -6 -8 106 248
use OR2X2  _12738_
timestamp 0
transform -1 0 13150 0 1 13690
box -6 -8 106 248
use AOI21X1  _12739_
timestamp 0
transform -1 0 12870 0 1 13690
box -6 -8 106 248
use OAI21X1  _12740_
timestamp 0
transform -1 0 11610 0 -1 14650
box -6 -8 106 248
use INVX1  _12741_
timestamp 0
transform -1 0 9090 0 1 10810
box -6 -8 66 248
use NAND2X1  _12742_
timestamp 0
transform 1 0 9250 0 1 11290
box -6 -8 86 248
use OAI21X1  _12743_
timestamp 0
transform 1 0 9150 0 1 10810
box -6 -8 106 248
use NAND2X1  _12744_
timestamp 0
transform -1 0 11810 0 -1 15130
box -6 -8 86 248
use AOI21X1  _12745_
timestamp 0
transform -1 0 13490 0 1 13210
box -6 -8 106 248
use MUX2X1  _12746_
timestamp 0
transform 1 0 15570 0 1 13210
box -6 -8 126 248
use MUX2X1  _12747_
timestamp 0
transform -1 0 15850 0 1 13210
box -6 -8 126 248
use MUX2X1  _12748_
timestamp 0
transform -1 0 15830 0 -1 13210
box -6 -8 126 248
use NAND2X1  _12749_
timestamp 0
transform -1 0 15470 0 -1 13210
box -6 -8 86 248
use OAI22X1  _12750_
timestamp 0
transform 1 0 15530 0 -1 13210
box -6 -8 126 248
use AOI21X1  _12751_
timestamp 0
transform 1 0 15250 0 -1 13210
box -6 -8 106 248
use AOI21X1  _12752_
timestamp 0
transform -1 0 13950 0 -1 13210
box -6 -8 106 248
use NAND2X1  _12753_
timestamp 0
transform 1 0 13710 0 -1 13210
box -6 -8 86 248
use INVX1  _12754_
timestamp 0
transform 1 0 14210 0 1 13210
box -6 -8 66 248
use OAI21X1  _12755_
timestamp 0
transform -1 0 14710 0 1 13210
box -6 -8 106 248
use NAND2X1  _12756_
timestamp 0
transform 1 0 14310 0 1 13210
box -6 -8 86 248
use AOI21X1  _12757_
timestamp 0
transform -1 0 13570 0 -1 13690
box -6 -8 106 248
use NAND3X1  _12758_
timestamp 0
transform -1 0 13710 0 -1 13690
box -6 -8 106 248
use INVX1  _12759_
timestamp 0
transform -1 0 13270 0 -1 13690
box -6 -8 66 248
use OR2X2  _12760_
timestamp 0
transform -1 0 13030 0 -1 13690
box -6 -8 106 248
use NOR2X1  _12761_
timestamp 0
transform -1 0 12990 0 1 13690
box -6 -8 86 248
use INVX1  _12762_
timestamp 0
transform -1 0 12470 0 1 13690
box -6 -8 66 248
use OAI21X1  _12763_
timestamp 0
transform 1 0 13070 0 -1 13690
box -6 -8 106 248
use AOI21X1  _12764_
timestamp 0
transform -1 0 12350 0 1 13690
box -6 -8 106 248
use INVX2  _12765_
timestamp 0
transform 1 0 12510 0 -1 15130
box -6 -8 66 248
use OAI21X1  _12766_
timestamp 0
transform -1 0 12350 0 -1 15130
box -6 -8 106 248
use OAI21X1  _12767_
timestamp 0
transform -1 0 12210 0 -1 15130
box -6 -8 106 248
use INVX1  _12768_
timestamp 0
transform 1 0 11830 0 1 14650
box -6 -8 66 248
use INVX2  _12769_
timestamp 0
transform 1 0 12410 0 -1 15130
box -6 -8 66 248
use OAI21X1  _12770_
timestamp 0
transform 1 0 13310 0 -1 13690
box -6 -8 106 248
use INVX1  _12771_
timestamp 0
transform -1 0 12830 0 -1 14170
box -6 -8 66 248
use INVX1  _12772_
timestamp 0
transform 1 0 15010 0 1 13690
box -6 -8 66 248
use NAND3X1  _12773_
timestamp 0
transform -1 0 14090 0 -1 13210
box -6 -8 106 248
use INVX1  _12774_
timestamp 0
transform 1 0 15190 0 -1 15610
box -6 -8 66 248
use NAND2X1  _12775_
timestamp 0
transform -1 0 15430 0 1 14650
box -6 -8 86 248
use OAI21X1  _12776_
timestamp 0
transform 1 0 15490 0 1 14650
box -6 -8 106 248
use NAND2X1  _12777_
timestamp 0
transform 1 0 15650 0 1 13690
box -6 -8 86 248
use OAI21X1  _12778_
timestamp 0
transform 1 0 15510 0 1 13690
box -6 -8 106 248
use NOR2X1  _12779_
timestamp 0
transform 1 0 17050 0 -1 14170
box -6 -8 86 248
use NOR2X1  _12780_
timestamp 0
transform 1 0 16830 0 -1 13690
box -6 -8 86 248
use AOI22X1  _12781_
timestamp 0
transform 1 0 16510 0 1 13690
box -6 -8 126 248
use OAI21X1  _12782_
timestamp 0
transform 1 0 15250 0 1 13690
box -6 -8 106 248
use NAND3X1  _12783_
timestamp 0
transform -1 0 13310 0 1 13690
box -6 -8 106 248
use INVX1  _12784_
timestamp 0
transform -1 0 13050 0 1 14170
box -6 -8 66 248
use INVX1  _12785_
timestamp 0
transform -1 0 13310 0 1 14170
box -6 -8 66 248
use OAI21X1  _12786_
timestamp 0
transform 1 0 13110 0 1 14170
box -6 -8 106 248
use NAND3X1  _12787_
timestamp 0
transform -1 0 13330 0 -1 14170
box -6 -8 106 248
use AOI21X1  _12788_
timestamp 0
transform 1 0 13390 0 -1 14170
box -6 -8 106 248
use INVX1  _12789_
timestamp 0
transform -1 0 13050 0 -1 14170
box -6 -8 66 248
use NAND2X1  _12790_
timestamp 0
transform -1 0 12950 0 -1 14170
box -6 -8 86 248
use AOI21X1  _12791_
timestamp 0
transform -1 0 12730 0 -1 14170
box -6 -8 106 248
use OAI21X1  _12792_
timestamp 0
transform -1 0 12570 0 -1 14170
box -6 -8 106 248
use AOI22X1  _12793_
timestamp 0
transform 1 0 11950 0 1 14650
box -6 -8 126 248
use AOI21X1  _12794_
timestamp 0
transform -1 0 13190 0 -1 14170
box -6 -8 106 248
use INVX1  _12795_
timestamp 0
transform -1 0 14150 0 -1 14170
box -6 -8 66 248
use INVX1  _12796_
timestamp 0
transform 1 0 14990 0 -1 15130
box -6 -8 66 248
use NAND2X1  _12797_
timestamp 0
transform 1 0 15410 0 1 14170
box -6 -8 86 248
use OAI21X1  _12798_
timestamp 0
transform 1 0 15270 0 1 14170
box -6 -8 106 248
use NAND2X1  _12799_
timestamp 0
transform -1 0 15470 0 1 13690
box -6 -8 86 248
use OAI21X1  _12800_
timestamp 0
transform -1 0 15510 0 -1 14170
box -6 -8 106 248
use NAND2X1  _12801_
timestamp 0
transform 1 0 15610 0 -1 13690
box -6 -8 86 248
use OAI21X1  _12802_
timestamp 0
transform -1 0 15210 0 1 13690
box -6 -8 106 248
use INVX2  _12803_
timestamp 0
transform -1 0 13570 0 1 13690
box -6 -8 66 248
use OAI21X1  _12804_
timestamp 0
transform -1 0 13750 0 1 14170
box -6 -8 106 248
use OR2X2  _12805_
timestamp 0
transform -1 0 13610 0 1 14170
box -6 -8 106 248
use NOR2X1  _12806_
timestamp 0
transform 1 0 13950 0 -1 14170
box -6 -8 86 248
use OAI21X1  _12807_
timestamp 0
transform 1 0 12830 0 -1 14650
box -6 -8 106 248
use NAND3X1  _12808_
timestamp 0
transform 1 0 13410 0 1 14650
box -6 -8 106 248
use NOR2X1  _12809_
timestamp 0
transform 1 0 13530 0 -1 14170
box -6 -8 86 248
use AND2X2  _12810_
timestamp 0
transform 1 0 13670 0 -1 14170
box -6 -8 106 248
use OAI21X1  _12811_
timestamp 0
transform 1 0 13810 0 -1 14170
box -6 -8 106 248
use NAND2X1  _12812_
timestamp 0
transform 1 0 12770 0 -1 15130
box -6 -8 86 248
use AOI21X1  _12813_
timestamp 0
transform -1 0 12970 0 1 15130
box -6 -8 106 248
use OAI21X1  _12814_
timestamp 0
transform 1 0 12730 0 1 15130
box -6 -8 106 248
use AOI22X1  _12815_
timestamp 0
transform 1 0 11990 0 1 15130
box -6 -8 126 248
use OAI21X1  _12816_
timestamp 0
transform -1 0 12710 0 -1 15130
box -6 -8 106 248
use INVX1  _12817_
timestamp 0
transform -1 0 14630 0 -1 14650
box -6 -8 66 248
use NAND3X1  _12818_
timestamp 0
transform 1 0 13350 0 1 14170
box -6 -8 106 248
use NAND2X1  _12819_
timestamp 0
transform 1 0 15690 0 1 14170
box -6 -8 86 248
use INVX1  _12820_
timestamp 0
transform 1 0 15830 0 -1 14170
box -6 -8 66 248
use AOI21X1  _12821_
timestamp 0
transform 1 0 15690 0 -1 14170
box -6 -8 106 248
use NAND2X1  _12822_
timestamp 0
transform 1 0 16430 0 -1 13690
box -6 -8 86 248
use OAI21X1  _12823_
timestamp 0
transform -1 0 15630 0 1 14170
box -6 -8 106 248
use NAND3X1  _12824_
timestamp 0
transform -1 0 13910 0 1 14170
box -6 -8 106 248
use NOR3X1  _12825_
timestamp 0
transform 1 0 13610 0 1 13690
box -6 -8 186 248
use INVX1  _12826_
timestamp 0
transform -1 0 14170 0 1 14170
box -6 -8 66 248
use OAI21X1  _12827_
timestamp 0
transform -1 0 13670 0 -1 14650
box -6 -8 106 248
use NAND3X1  _12828_
timestamp 0
transform -1 0 13370 0 -1 14650
box -6 -8 106 248
use AOI21X1  _12829_
timestamp 0
transform -1 0 13230 0 -1 14650
box -6 -8 106 248
use INVX1  _12830_
timestamp 0
transform -1 0 13370 0 1 14650
box -6 -8 66 248
use NAND2X1  _12831_
timestamp 0
transform 1 0 13150 0 1 15130
box -6 -8 86 248
use AND2X2  _12832_
timestamp 0
transform -1 0 12670 0 1 15130
box -6 -8 106 248
use OAI21X1  _12833_
timestamp 0
transform -1 0 12530 0 1 15130
box -6 -8 106 248
use OAI21X1  _12834_
timestamp 0
transform -1 0 12390 0 1 15130
box -6 -8 106 248
use OAI21X1  _12835_
timestamp 0
transform 1 0 11510 0 -1 15610
box -6 -8 106 248
use INVX1  _12836_
timestamp 0
transform 1 0 12190 0 -1 15610
box -6 -8 66 248
use INVX1  _12837_
timestamp 0
transform -1 0 13610 0 1 15130
box -6 -8 66 248
use NAND3X1  _12838_
timestamp 0
transform 1 0 13430 0 -1 14650
box -6 -8 106 248
use AOI21X1  _12839_
timestamp 0
transform -1 0 15650 0 -1 14170
box -6 -8 106 248
use NAND2X1  _12840_
timestamp 0
transform 1 0 15350 0 -1 13690
box -6 -8 86 248
use OAI21X1  _12841_
timestamp 0
transform -1 0 15450 0 -1 14650
box -6 -8 106 248
use NAND3X1  _12842_
timestamp 0
transform -1 0 13590 0 -1 15130
box -6 -8 106 248
use INVX1  _12843_
timestamp 0
transform -1 0 14190 0 1 14650
box -6 -8 66 248
use OAI21X1  _12844_
timestamp 0
transform 1 0 13950 0 1 14170
box -6 -8 106 248
use NAND2X1  _12845_
timestamp 0
transform 1 0 13850 0 1 14650
box -6 -8 86 248
use NAND3X1  _12846_
timestamp 0
transform -1 0 13370 0 1 15130
box -6 -8 106 248
use NAND3X1  _12847_
timestamp 0
transform -1 0 13790 0 1 14650
box -6 -8 106 248
use NAND2X1  _12848_
timestamp 0
transform 1 0 13990 0 1 14650
box -6 -8 86 248
use NAND3X1  _12849_
timestamp 0
transform -1 0 13650 0 1 14650
box -6 -8 106 248
use NAND2X1  _12850_
timestamp 0
transform -1 0 12850 0 -1 15610
box -6 -8 86 248
use AOI21X1  _12851_
timestamp 0
transform -1 0 13070 0 -1 14650
box -6 -8 106 248
use NOR2X1  _12852_
timestamp 0
transform 1 0 13030 0 1 14650
box -6 -8 86 248
use OAI21X1  _12853_
timestamp 0
transform 1 0 12910 0 -1 15130
box -6 -8 106 248
use NAND2X1  _12854_
timestamp 0
transform -1 0 13090 0 1 15130
box -6 -8 86 248
use AOI21X1  _12855_
timestamp 0
transform -1 0 12550 0 1 15610
box -6 -8 106 248
use OAI21X1  _12856_
timestamp 0
transform -1 0 12570 0 -1 15610
box -6 -8 106 248
use AOI22X1  _12857_
timestamp 0
transform 1 0 12310 0 -1 15610
box -6 -8 126 248
use INVX1  _12858_
timestamp 0
transform 1 0 11890 0 1 15610
box -6 -8 66 248
use AOI21X1  _12859_
timestamp 0
transform 1 0 13410 0 1 15130
box -6 -8 106 248
use AND2X2  _12860_
timestamp 0
transform -1 0 13450 0 -1 15130
box -6 -8 106 248
use NAND3X1  _12861_
timestamp 0
transform -1 0 13290 0 -1 15130
box -6 -8 106 248
use AOI21X1  _12862_
timestamp 0
transform 1 0 13170 0 1 14650
box -6 -8 106 248
use OAI21X1  _12863_
timestamp 0
transform 1 0 13050 0 -1 15130
box -6 -8 106 248
use AOI21X1  _12864_
timestamp 0
transform -1 0 13250 0 -1 15610
box -6 -8 106 248
use INVX1  _12865_
timestamp 0
transform -1 0 13990 0 1 15130
box -6 -8 66 248
use NAND3X1  _12866_
timestamp 0
transform 1 0 13710 0 -1 14650
box -6 -8 106 248
use INVX1  _12867_
timestamp 0
transform 1 0 15250 0 1 14650
box -6 -8 66 248
use NOR2X1  _12868_
timestamp 0
transform -1 0 15430 0 -1 15130
box -6 -8 86 248
use INVX1  _12869_
timestamp 0
transform -1 0 15330 0 1 15130
box -6 -8 66 248
use OAI21X1  _12870_
timestamp 0
transform 1 0 14730 0 -1 15130
box -6 -8 106 248
use NAND3X1  _12871_
timestamp 0
transform -1 0 13890 0 1 15130
box -6 -8 106 248
use INVX1  _12872_
timestamp 0
transform -1 0 14410 0 -1 15130
box -6 -8 66 248
use OAI21X1  _12873_
timestamp 0
transform 1 0 13630 0 -1 15130
box -6 -8 106 248
use NAND2X1  _12874_
timestamp 0
transform 1 0 13790 0 -1 15130
box -6 -8 86 248
use NAND3X1  _12875_
timestamp 0
transform -1 0 13750 0 1 15130
box -6 -8 106 248
use NAND3X1  _12876_
timestamp 0
transform 1 0 14070 0 -1 15130
box -6 -8 106 248
use NAND2X1  _12877_
timestamp 0
transform 1 0 14210 0 -1 15130
box -6 -8 86 248
use NAND3X1  _12878_
timestamp 0
transform -1 0 14010 0 -1 15130
box -6 -8 106 248
use NAND2X1  _12879_
timestamp 0
transform -1 0 13110 0 1 15610
box -6 -8 86 248
use INVX1  _12880_
timestamp 0
transform -1 0 12950 0 -1 15610
box -6 -8 66 248
use NOR2X1  _12881_
timestamp 0
transform 1 0 13010 0 -1 15610
box -6 -8 86 248
use OAI21X1  _12882_
timestamp 0
transform 1 0 12610 0 -1 15610
box -6 -8 106 248
use OAI21X1  _12883_
timestamp 0
transform -1 0 12390 0 1 15610
box -6 -8 106 248
use OAI21X1  _12884_
timestamp 0
transform -1 0 12190 0 -1 16090
box -6 -8 106 248
use INVX1  _12885_
timestamp 0
transform -1 0 12030 0 -1 16090
box -6 -8 66 248
use OAI21X1  _12886_
timestamp 0
transform -1 0 12250 0 1 15610
box -6 -8 106 248
use OAI21X1  _12887_
timestamp 0
transform 1 0 11990 0 1 15610
box -6 -8 106 248
use INVX1  _12888_
timestamp 0
transform -1 0 11510 0 -1 16090
box -6 -8 66 248
use OAI21X1  _12889_
timestamp 0
transform 1 0 12870 0 1 15610
box -6 -8 106 248
use NOR2X1  _12890_
timestamp 0
transform -1 0 12670 0 1 15610
box -6 -8 86 248
use AOI21X1  _12891_
timestamp 0
transform -1 0 12830 0 1 15610
box -6 -8 106 248
use INVX1  _12892_
timestamp 0
transform 1 0 13590 0 1 15610
box -6 -8 66 248
use OR2X2  _12893_
timestamp 0
transform -1 0 13970 0 -1 15610
box -6 -8 106 248
use OAI21X1  _12894_
timestamp 0
transform 1 0 14690 0 1 15130
box -6 -8 106 248
use NAND3X1  _12895_
timestamp 0
transform -1 0 13810 0 1 15610
box -6 -8 106 248
use NOR2X1  _12896_
timestamp 0
transform 1 0 14010 0 -1 15610
box -6 -8 86 248
use INVX1  _12897_
timestamp 0
transform 1 0 14170 0 1 15610
box -6 -8 66 248
use OAI21X1  _12898_
timestamp 0
transform 1 0 14030 0 1 15610
box -6 -8 106 248
use NAND3X1  _12899_
timestamp 0
transform -1 0 13550 0 1 15610
box -6 -8 106 248
use NAND3X1  _12900_
timestamp 0
transform -1 0 13970 0 1 15610
box -6 -8 106 248
use OAI21X1  _12901_
timestamp 0
transform -1 0 13810 0 -1 15610
box -6 -8 106 248
use NAND3X1  _12902_
timestamp 0
transform -1 0 13670 0 -1 16090
box -6 -8 106 248
use AND2X2  _12903_
timestamp 0
transform -1 0 13490 0 1 16090
box -6 -8 106 248
use INVX1  _12904_
timestamp 0
transform -1 0 12590 0 -1 16090
box -6 -8 66 248
use AOI21X1  _12905_
timestamp 0
transform -1 0 12490 0 -1 16090
box -6 -8 106 248
use OAI21X1  _12906_
timestamp 0
transform -1 0 12330 0 -1 16090
box -6 -8 106 248
use AOI22X1  _12907_
timestamp 0
transform 1 0 11810 0 -1 16090
box -6 -8 126 248
use NAND2X1  _12908_
timestamp 0
transform 1 0 13590 0 -1 15610
box -6 -8 86 248
use AND2X2  _12909_
timestamp 0
transform -1 0 13550 0 -1 15610
box -6 -8 106 248
use AND2X2  _12910_
timestamp 0
transform 1 0 13310 0 -1 15610
box -6 -8 106 248
use NAND3X1  _12911_
timestamp 0
transform -1 0 13410 0 1 15610
box -6 -8 106 248
use OAI21X1  _12912_
timestamp 0
transform 1 0 13170 0 1 15610
box -6 -8 106 248
use INVX1  _12913_
timestamp 0
transform -1 0 13410 0 -1 16090
box -6 -8 66 248
use AOI21X1  _12914_
timestamp 0
transform 1 0 13230 0 1 16090
box -6 -8 106 248
use INVX1  _12915_
timestamp 0
transform 1 0 14290 0 -1 15610
box -6 -8 66 248
use NOR3X1  _12916_
timestamp 0
transform 1 0 14030 0 1 15130
box -6 -8 186 248
use INVX1  _12917_
timestamp 0
transform 1 0 14710 0 -1 15610
box -6 -8 66 248
use OAI21X1  _12918_
timestamp 0
transform 1 0 14970 0 1 15130
box -6 -8 106 248
use NAND3X1  _12919_
timestamp 0
transform -1 0 14650 0 -1 15610
box -6 -8 106 248
use INVX1  _12920_
timestamp 0
transform 1 0 14810 0 -1 15610
box -6 -8 66 248
use OAI21X1  _12921_
timestamp 0
transform 1 0 14570 0 1 15610
box -6 -8 106 248
use NAND3X1  _12922_
timestamp 0
transform 1 0 14430 0 1 15610
box -6 -8 106 248
use NAND3X1  _12923_
timestamp 0
transform 1 0 14390 0 -1 15610
box -6 -8 106 248
use OAI21X1  _12924_
timestamp 0
transform 1 0 14550 0 1 15130
box -6 -8 106 248
use NAND3X1  _12925_
timestamp 0
transform -1 0 14230 0 -1 15610
box -6 -8 106 248
use AND2X2  _12926_
timestamp 0
transform -1 0 13650 0 1 16090
box -6 -8 106 248
use AND2X2  _12927_
timestamp 0
transform -1 0 12190 0 1 16090
box -6 -8 106 248
use OAI21X1  _12928_
timestamp 0
transform -1 0 12330 0 1 16090
box -6 -8 106 248
use OAI21X1  _12929_
timestamp 0
transform -1 0 12050 0 1 16090
box -6 -8 106 248
use OAI21X1  _12930_
timestamp 0
transform 1 0 11070 0 1 16570
box -6 -8 106 248
use INVX1  _12931_
timestamp 0
transform 1 0 15110 0 -1 15130
box -6 -8 66 248
use OAI21X1  _12932_
timestamp 0
transform -1 0 15310 0 -1 15130
box -6 -8 106 248
use INVX1  _12933_
timestamp 0
transform -1 0 15170 0 1 15610
box -6 -8 66 248
use AOI21X1  _12934_
timestamp 0
transform 1 0 14970 0 1 15610
box -6 -8 106 248
use NAND3X1  _12935_
timestamp 0
transform 1 0 14810 0 1 15610
box -6 -8 106 248
use NAND2X1  _12936_
timestamp 0
transform -1 0 14090 0 -1 16090
box -6 -8 86 248
use NAND2X1  _12937_
timestamp 0
transform 1 0 15210 0 1 15610
box -6 -8 86 248
use OAI21X1  _12938_
timestamp 0
transform -1 0 14650 0 -1 16090
box -6 -8 106 248
use NAND2X1  _12939_
timestamp 0
transform 1 0 14410 0 -1 16090
box -6 -8 86 248
use INVX1  _12940_
timestamp 0
transform 1 0 14710 0 1 15610
box -6 -8 66 248
use AND2X2  _12941_
timestamp 0
transform -1 0 13950 0 -1 16090
box -6 -8 106 248
use NAND2X1  _12942_
timestamp 0
transform -1 0 14210 0 -1 16090
box -6 -8 86 248
use NAND3X1  _12943_
timestamp 0
transform -1 0 14370 0 -1 16090
box -6 -8 106 248
use NAND2X1  _12944_
timestamp 0
transform -1 0 12990 0 -1 16090
box -6 -8 86 248
use AOI21X1  _12945_
timestamp 0
transform -1 0 14370 0 1 15610
box -6 -8 106 248
use AOI21X1  _12946_
timestamp 0
transform -1 0 13310 0 -1 16090
box -6 -8 106 248
use NAND3X1  _12947_
timestamp 0
transform -1 0 13190 0 1 16090
box -6 -8 106 248
use AOI21X1  _12948_
timestamp 0
transform -1 0 13050 0 1 16090
box -6 -8 106 248
use AND2X2  _12949_
timestamp 0
transform -1 0 12870 0 -1 16090
box -6 -8 106 248
use NAND3X1  _12950_
timestamp 0
transform -1 0 13150 0 -1 16090
box -6 -8 106 248
use OAI21X1  _12951_
timestamp 0
transform -1 0 12730 0 -1 16090
box -6 -8 106 248
use OAI21X1  _12952_
timestamp 0
transform -1 0 12630 0 1 16090
box -6 -8 106 248
use OR2X2  _12953_
timestamp 0
transform -1 0 12490 0 1 16090
box -6 -8 106 248
use AOI22X1  _12954_
timestamp 0
transform 1 0 11770 0 1 16090
box -6 -8 126 248
use NAND2X1  _12955_
timestamp 0
transform 1 0 11970 0 -1 16570
box -6 -8 86 248
use INVX1  _12956_
timestamp 0
transform -1 0 12890 0 1 16090
box -6 -8 66 248
use NAND2X1  _12957_
timestamp 0
transform 1 0 15130 0 1 15130
box -6 -8 86 248
use INVX1  _12958_
timestamp 0
transform 1 0 15470 0 -1 15130
box -6 -8 66 248
use NAND2X1  _12959_
timestamp 0
transform -1 0 14950 0 -1 15130
box -6 -8 86 248
use NAND2X1  _12960_
timestamp 0
transform -1 0 14930 0 1 15130
box -6 -8 86 248
use INVX1  _12961_
timestamp 0
transform 1 0 13810 0 1 16090
box -6 -8 66 248
use NAND2X1  _12962_
timestamp 0
transform 1 0 13930 0 1 16090
box -6 -8 86 248
use NAND2X1  _12963_
timestamp 0
transform -1 0 13790 0 -1 16090
box -6 -8 86 248
use NAND2X1  _12964_
timestamp 0
transform -1 0 13770 0 1 16090
box -6 -8 86 248
use INVX1  _12965_
timestamp 0
transform 1 0 13210 0 -1 16570
box -6 -8 66 248
use NOR3X1  _12966_
timestamp 0
transform -1 0 13010 0 -1 16570
box -6 -8 186 248
use AOI21X1  _12967_
timestamp 0
transform 1 0 12690 0 1 16090
box -6 -8 106 248
use OAI21X1  _12968_
timestamp 0
transform -1 0 13150 0 -1 16570
box -6 -8 106 248
use OAI21X1  _12969_
timestamp 0
transform -1 0 12790 0 -1 16570
box -6 -8 106 248
use NAND2X1  _12970_
timestamp 0
transform 1 0 12250 0 -1 16570
box -6 -8 86 248
use NAND2X1  _12971_
timestamp 0
transform -1 0 12990 0 1 14650
box -6 -8 86 248
use INVX1  _12972_
timestamp 0
transform 1 0 15750 0 -1 13690
box -6 -8 66 248
use NAND2X1  _12973_
timestamp 0
transform -1 0 15930 0 -1 13690
box -6 -8 86 248
use OAI21X1  _12974_
timestamp 0
transform -1 0 16090 0 -1 13690
box -6 -8 106 248
use NAND2X1  _12975_
timestamp 0
transform 1 0 16290 0 -1 13690
box -6 -8 86 248
use NOR2X1  _12976_
timestamp 0
transform 1 0 14070 0 -1 12730
box -6 -8 86 248
use NOR2X1  _12977_
timestamp 0
transform -1 0 14170 0 1 12250
box -6 -8 86 248
use AOI22X1  _12978_
timestamp 0
transform 1 0 14190 0 -1 12730
box -6 -8 126 248
use NAND3X1  _12979_
timestamp 0
transform -1 0 16250 0 -1 13690
box -6 -8 106 248
use NAND2X1  _12980_
timestamp 0
transform -1 0 14530 0 -1 15130
box -6 -8 86 248
use OAI21X1  _12981_
timestamp 0
transform 1 0 14590 0 -1 15130
box -6 -8 106 248
use NAND2X1  _12982_
timestamp 0
transform -1 0 14830 0 1 14170
box -6 -8 86 248
use OAI21X1  _12983_
timestamp 0
transform -1 0 14970 0 1 14170
box -6 -8 106 248
use MUX2X1  _12984_
timestamp 0
transform 1 0 16250 0 -1 15130
box -6 -8 126 248
use NAND2X1  _12985_
timestamp 0
transform -1 0 16490 0 -1 15130
box -6 -8 86 248
use AND2X2  _12986_
timestamp 0
transform 1 0 16670 0 -1 250
box -6 -8 106 248
use NOR2X1  _12987_
timestamp 0
transform -1 0 15890 0 1 14170
box -6 -8 86 248
use NAND2X1  _12988_
timestamp 0
transform -1 0 15950 0 -1 15130
box -6 -8 86 248
use NAND2X1  _12989_
timestamp 0
transform 1 0 16110 0 -1 15130
box -6 -8 86 248
use NAND2X1  _12990_
timestamp 0
transform 1 0 15990 0 -1 15130
box -6 -8 86 248
use OAI21X1  _12991_
timestamp 0
transform 1 0 16070 0 1 14650
box -6 -8 106 248
use OAI21X1  _12992_
timestamp 0
transform -1 0 15890 0 1 14650
box -6 -8 106 248
use OAI21X1  _12993_
timestamp 0
transform -1 0 15750 0 1 14650
box -6 -8 106 248
use NAND2X1  _12994_
timestamp 0
transform 1 0 12370 0 -1 14650
box -6 -8 86 248
use NOR2X1  _12995_
timestamp 0
transform -1 0 16010 0 1 14650
box -6 -8 86 248
use NAND2X1  _12996_
timestamp 0
transform -1 0 15210 0 -1 14170
box -6 -8 86 248
use OAI21X1  _12997_
timestamp 0
transform -1 0 15350 0 -1 14170
box -6 -8 106 248
use NAND2X1  _12998_
timestamp 0
transform -1 0 15570 0 -1 13690
box -6 -8 86 248
use OAI21X1  _12999_
timestamp 0
transform 1 0 15210 0 -1 13690
box -6 -8 106 248
use MUX2X1  _13000_
timestamp 0
transform -1 0 16610 0 -1 14170
box -6 -8 126 248
use NAND2X1  _13001_
timestamp 0
transform 1 0 16610 0 -1 14650
box -6 -8 86 248
use NAND2X1  _13002_
timestamp 0
transform 1 0 14410 0 1 15130
box -6 -8 86 248
use OAI21X1  _13003_
timestamp 0
transform 1 0 14270 0 1 15130
box -6 -8 106 248
use INVX1  _13004_
timestamp 0
transform 1 0 16050 0 1 14170
box -6 -8 66 248
use NAND2X1  _13005_
timestamp 0
transform -1 0 14310 0 1 14170
box -6 -8 86 248
use OAI21X1  _13006_
timestamp 0
transform -1 0 14450 0 1 14170
box -6 -8 106 248
use NAND2X1  _13007_
timestamp 0
transform 1 0 16470 0 1 14170
box -6 -8 86 248
use OAI21X1  _13008_
timestamp 0
transform 1 0 16310 0 1 14170
box -6 -8 106 248
use OAI21X1  _13009_
timestamp 0
transform 1 0 16470 0 -1 14650
box -6 -8 106 248
use NAND3X1  _13010_
timestamp 0
transform -1 0 17110 0 1 12250
box -6 -8 106 248
use MUX2X1  _13011_
timestamp 0
transform 1 0 16150 0 1 14170
box -6 -8 126 248
use MUX2X1  _13012_
timestamp 0
transform -1 0 16850 0 1 14170
box -6 -8 126 248
use OAI21X1  _13013_
timestamp 0
transform 1 0 16530 0 1 14650
box -6 -8 106 248
use AOI21X1  _13014_
timestamp 0
transform -1 0 16290 0 -1 14650
box -6 -8 106 248
use INVX1  _13015_
timestamp 0
transform 1 0 15950 0 -1 14650
box -6 -8 66 248
use NAND3X1  _13016_
timestamp 0
transform -1 0 16430 0 -1 14650
box -6 -8 106 248
use AND2X2  _13017_
timestamp 0
transform -1 0 15890 0 -1 14650
box -6 -8 106 248
use NAND2X1  _13018_
timestamp 0
transform 1 0 15650 0 -1 14650
box -6 -8 86 248
use OR2X2  _13019_
timestamp 0
transform -1 0 15610 0 -1 14650
box -6 -8 106 248
use AOI21X1  _13020_
timestamp 0
transform 1 0 14410 0 -1 14650
box -6 -8 106 248
use OAI21X1  _13021_
timestamp 0
transform -1 0 12590 0 -1 14650
box -6 -8 106 248
use NAND2X1  _13022_
timestamp 0
transform -1 0 12370 0 1 14650
box -6 -8 86 248
use AOI21X1  _13023_
timestamp 0
transform 1 0 16050 0 -1 14650
box -6 -8 106 248
use NAND2X1  _13024_
timestamp 0
transform 1 0 16670 0 -1 17050
box -6 -8 86 248
use NAND2X1  _13025_
timestamp 0
transform 1 0 15050 0 -1 15610
box -6 -8 86 248
use OAI21X1  _13026_
timestamp 0
transform 1 0 14910 0 -1 15610
box -6 -8 106 248
use NAND2X1  _13027_
timestamp 0
transform 1 0 16150 0 -1 15610
box -6 -8 86 248
use OAI21X1  _13028_
timestamp 0
transform 1 0 15990 0 -1 15610
box -6 -8 106 248
use NAND2X1  _13029_
timestamp 0
transform -1 0 16290 0 1 13690
box -6 -8 86 248
use NAND2X1  _13030_
timestamp 0
transform 1 0 16350 0 -1 14170
box -6 -8 86 248
use NAND2X1  _13031_
timestamp 0
transform -1 0 16310 0 -1 14170
box -6 -8 86 248
use AOI21X1  _13032_
timestamp 0
transform -1 0 16290 0 1 15130
box -6 -8 106 248
use INVX1  _13033_
timestamp 0
transform 1 0 17090 0 -1 12250
box -6 -8 66 248
use NAND3X1  _13034_
timestamp 0
transform -1 0 16910 0 -1 17050
box -6 -8 106 248
use AOI21X1  _13035_
timestamp 0
transform 1 0 16810 0 1 14650
box -6 -8 106 248
use OAI21X1  _13036_
timestamp 0
transform 1 0 16970 0 1 14650
box -6 -8 106 248
use NAND3X1  _13037_
timestamp 0
transform 1 0 16770 0 1 250
box -6 -8 106 248
use INVX1  _13038_
timestamp 0
transform 1 0 16870 0 -1 14650
box -6 -8 66 248
use AOI21X1  _13039_
timestamp 0
transform 1 0 16970 0 -1 14650
box -6 -8 106 248
use NOR2X1  _13040_
timestamp 0
transform -1 0 16810 0 -1 14650
box -6 -8 86 248
use AND2X2  _13041_
timestamp 0
transform -1 0 16490 0 1 14650
box -6 -8 106 248
use NOR2X1  _13042_
timestamp 0
transform 1 0 15050 0 -1 17050
box -6 -8 86 248
use OAI21X1  _13043_
timestamp 0
transform -1 0 16330 0 1 14650
box -6 -8 106 248
use OAI21X1  _13044_
timestamp 0
transform -1 0 12870 0 1 14650
box -6 -8 106 248
use OAI21X1  _13045_
timestamp 0
transform 1 0 16670 0 1 14650
box -6 -8 106 248
use INVX1  _13046_
timestamp 0
transform -1 0 16770 0 -1 15610
box -6 -8 66 248
use NAND2X1  _13047_
timestamp 0
transform -1 0 15410 0 1 15610
box -6 -8 86 248
use OAI21X1  _13048_
timestamp 0
transform -1 0 15570 0 1 15610
box -6 -8 106 248
use MUX2X1  _13049_
timestamp 0
transform -1 0 15630 0 1 15130
box -6 -8 126 248
use NOR2X1  _13050_
timestamp 0
transform 1 0 16070 0 1 15130
box -6 -8 86 248
use NAND2X1  _13051_
timestamp 0
transform 1 0 16650 0 -1 14170
box -6 -8 86 248
use NAND2X1  _13052_
timestamp 0
transform -1 0 16850 0 -1 14170
box -6 -8 86 248
use NAND2X1  _13053_
timestamp 0
transform -1 0 16990 0 -1 14170
box -6 -8 86 248
use OR2X2  _13054_
timestamp 0
transform 1 0 16970 0 -1 15130
box -6 -8 106 248
use OAI21X1  _13055_
timestamp 0
transform 1 0 16970 0 -1 17050
box -6 -8 106 248
use OR2X2  _13056_
timestamp 0
transform -1 0 16610 0 -1 17050
box -6 -8 106 248
use OAI21X1  _13057_
timestamp 0
transform 1 0 17030 0 1 3130
box -6 -8 106 248
use AOI21X1  _13058_
timestamp 0
transform 1 0 17050 0 1 15130
box -6 -8 106 248
use INVX1  _13059_
timestamp 0
transform 1 0 16950 0 -1 15610
box -6 -8 66 248
use NAND3X1  _13060_
timestamp 0
transform -1 0 16990 0 1 15130
box -6 -8 106 248
use NAND2X1  _13061_
timestamp 0
transform 1 0 17050 0 -1 15610
box -6 -8 86 248
use OR2X2  _13062_
timestamp 0
transform -1 0 16710 0 1 15130
box -6 -8 106 248
use NAND2X1  _13063_
timestamp 0
transform 1 0 16750 0 1 15130
box -6 -8 86 248
use NAND2X1  _13064_
timestamp 0
transform 1 0 16470 0 1 15130
box -6 -8 86 248
use AOI22X1  _13065_
timestamp 0
transform 1 0 12650 0 -1 14650
box -6 -8 126 248
use AOI21X1  _13066_
timestamp 0
transform 1 0 16810 0 -1 15610
box -6 -8 106 248
use NAND2X1  _13067_
timestamp 0
transform -1 0 15470 0 1 15130
box -6 -8 86 248
use OAI21X1  _13068_
timestamp 0
transform 1 0 15290 0 -1 15610
box -6 -8 106 248
use NAND2X1  _13069_
timestamp 0
transform -1 0 15810 0 -1 15610
box -6 -8 86 248
use OAI21X1  _13070_
timestamp 0
transform -1 0 15950 0 -1 15610
box -6 -8 106 248
use NAND2X1  _13071_
timestamp 0
transform 1 0 16410 0 -1 15610
box -6 -8 86 248
use OAI21X1  _13072_
timestamp 0
transform 1 0 16550 0 -1 15610
box -6 -8 106 248
use INVX1  _13073_
timestamp 0
transform 1 0 17070 0 -1 16090
box -6 -8 66 248
use NAND3X1  _13074_
timestamp 0
transform 1 0 16550 0 -1 15130
box -6 -8 106 248
use OAI21X1  _13075_
timestamp 0
transform -1 0 17010 0 1 15610
box -6 -8 106 248
use OR2X2  _13076_
timestamp 0
transform -1 0 17030 0 -1 16090
box -6 -8 106 248
use NOR2X1  _13077_
timestamp 0
transform -1 0 17150 0 1 15610
box -6 -8 86 248
use OAI21X1  _13078_
timestamp 0
transform -1 0 16890 0 -1 16090
box -6 -8 106 248
use NAND3X1  _13079_
timestamp 0
transform -1 0 16750 0 -1 16090
box -6 -8 106 248
use OR2X2  _13080_
timestamp 0
transform -1 0 17010 0 1 16090
box -6 -8 106 248
use OAI21X1  _13081_
timestamp 0
transform -1 0 16870 0 1 16090
box -6 -8 106 248
use NAND3X1  _13082_
timestamp 0
transform -1 0 16810 0 -1 16570
box -6 -8 106 248
use NAND2X1  _13083_
timestamp 0
transform -1 0 16670 0 -1 16570
box -6 -8 86 248
use OR2X2  _13084_
timestamp 0
transform 1 0 14490 0 -1 17050
box -6 -8 106 248
use NAND2X1  _13085_
timestamp 0
transform -1 0 16390 0 1 16570
box -6 -8 86 248
use NAND2X1  _13086_
timestamp 0
transform -1 0 16270 0 1 16570
box -6 -8 86 248
use AOI22X1  _13087_
timestamp 0
transform 1 0 11830 0 1 16570
box -6 -8 126 248
use INVX1  _13088_
timestamp 0
transform -1 0 12330 0 1 16570
box -6 -8 66 248
use OAI21X1  _13089_
timestamp 0
transform 1 0 16450 0 1 16570
box -6 -8 106 248
use NAND2X1  _13090_
timestamp 0
transform 1 0 17050 0 1 16090
box -6 -8 86 248
use NOR2X1  _13091_
timestamp 0
transform -1 0 15670 0 -1 15130
box -6 -8 86 248
use AOI21X1  _13092_
timestamp 0
transform -1 0 15530 0 -1 15610
box -6 -8 106 248
use NAND2X1  _13093_
timestamp 0
transform 1 0 16350 0 1 15130
box -6 -8 86 248
use OAI21X1  _13094_
timestamp 0
transform 1 0 16270 0 -1 15610
box -6 -8 106 248
use INVX1  _13095_
timestamp 0
transform -1 0 16550 0 1 16090
box -6 -8 66 248
use NAND3X1  _13096_
timestamp 0
transform 1 0 17030 0 -1 16570
box -6 -8 106 248
use NOR2X1  _13097_
timestamp 0
transform -1 0 16930 0 -1 15130
box -6 -8 86 248
use NAND3X1  _13098_
timestamp 0
transform 1 0 16710 0 -1 15130
box -6 -8 106 248
use OAI21X1  _13099_
timestamp 0
transform 1 0 16770 0 1 15610
box -6 -8 106 248
use NAND2X1  _13100_
timestamp 0
transform 1 0 16650 0 1 15610
box -6 -8 86 248
use AOI21X1  _13101_
timestamp 0
transform -1 0 16690 0 1 16570
box -6 -8 106 248
use INVX1  _13102_
timestamp 0
transform -1 0 16130 0 1 16570
box -6 -8 66 248
use NAND3X1  _13103_
timestamp 0
transform 1 0 16750 0 1 16570
box -6 -8 106 248
use NAND2X1  _13104_
timestamp 0
transform 1 0 15950 0 1 16570
box -6 -8 86 248
use NOR2X1  _13105_
timestamp 0
transform 1 0 15830 0 1 16570
box -6 -8 86 248
use AND2X2  _13106_
timestamp 0
transform -1 0 15770 0 1 16570
box -6 -8 106 248
use OAI21X1  _13107_
timestamp 0
transform -1 0 15630 0 1 16570
box -6 -8 106 248
use OAI21X1  _13108_
timestamp 0
transform 1 0 12630 0 1 16570
box -6 -8 106 248
use INVX1  _13109_
timestamp 0
transform 1 0 9550 0 -1 17050
box -6 -8 66 248
use NAND3X1  _13110_
timestamp 0
transform 1 0 16610 0 1 16090
box -6 -8 106 248
use AOI21X1  _13111_
timestamp 0
transform 1 0 15570 0 -1 15610
box -6 -8 106 248
use NAND2X1  _13112_
timestamp 0
transform -1 0 16210 0 1 15610
box -6 -8 86 248
use OAI21X1  _13113_
timestamp 0
transform 1 0 16250 0 1 15610
box -6 -8 106 248
use NAND3X1  _13114_
timestamp 0
transform -1 0 16350 0 -1 16090
box -6 -8 106 248
use NOR3X1  _13115_
timestamp 0
transform -1 0 16590 0 -1 16090
box -6 -8 186 248
use INVX1  _13116_
timestamp 0
transform 1 0 16390 0 1 16090
box -6 -8 66 248
use OAI21X1  _13117_
timestamp 0
transform 1 0 16250 0 1 16090
box -6 -8 106 248
use NAND2X1  _13118_
timestamp 0
transform -1 0 16070 0 -1 16090
box -6 -8 86 248
use NAND2X1  _13119_
timestamp 0
transform 1 0 15990 0 1 15610
box -6 -8 86 248
use NAND3X1  _13120_
timestamp 0
transform -1 0 16210 0 -1 16090
box -6 -8 106 248
use NAND2X1  _13121_
timestamp 0
transform 1 0 13650 0 -1 17050
box -6 -8 86 248
use AOI21X1  _13122_
timestamp 0
transform 1 0 16870 0 -1 16570
box -6 -8 106 248
use NOR2X1  _13123_
timestamp 0
transform 1 0 14930 0 -1 17050
box -6 -8 86 248
use OAI21X1  _13124_
timestamp 0
transform -1 0 14430 0 -1 17050
box -6 -8 106 248
use NAND2X1  _13125_
timestamp 0
transform -1 0 14110 0 -1 17050
box -6 -8 86 248
use NOR2X1  _13126_
timestamp 0
transform 1 0 13770 0 -1 17050
box -6 -8 86 248
use AND2X2  _13127_
timestamp 0
transform -1 0 13190 0 -1 17050
box -6 -8 106 248
use AND2X2  _13128_
timestamp 0
transform -1 0 16550 0 -1 16570
box -6 -8 106 248
use NAND3X1  _13129_
timestamp 0
transform -1 0 14750 0 -1 17050
box -6 -8 106 248
use AOI21X1  _13130_
timestamp 0
transform -1 0 14890 0 -1 17050
box -6 -8 106 248
use OAI21X1  _13131_
timestamp 0
transform -1 0 14270 0 -1 17050
box -6 -8 106 248
use NOR2X1  _13132_
timestamp 0
transform -1 0 13030 0 -1 17050
box -6 -8 86 248
use OAI21X1  _13133_
timestamp 0
transform -1 0 12230 0 -1 17050
box -6 -8 106 248
use NAND2X1  _13134_
timestamp 0
transform 1 0 9810 0 -1 17050
box -6 -8 86 248
use OAI21X1  _13135_
timestamp 0
transform 1 0 9650 0 -1 17050
box -6 -8 106 248
use INVX1  _13136_
timestamp 0
transform 1 0 11330 0 -1 17050
box -6 -8 66 248
use INVX1  _13137_
timestamp 0
transform -1 0 12490 0 -1 17050
box -6 -8 66 248
use NAND2X1  _13138_
timestamp 0
transform 1 0 15990 0 1 16090
box -6 -8 86 248
use NOR2X1  _13139_
timestamp 0
transform -1 0 15810 0 -1 15130
box -6 -8 86 248
use INVX1  _13140_
timestamp 0
transform 1 0 15670 0 1 15130
box -6 -8 66 248
use OAI21X1  _13141_
timestamp 0
transform 1 0 15570 0 -1 16090
box -6 -8 106 248
use NAND3X1  _13142_
timestamp 0
transform -1 0 15730 0 -1 16570
box -6 -8 106 248
use INVX1  _13143_
timestamp 0
transform 1 0 16130 0 1 16090
box -6 -8 66 248
use OAI21X1  _13144_
timestamp 0
transform -1 0 16410 0 -1 16570
box -6 -8 106 248
use NAND2X1  _13145_
timestamp 0
transform 1 0 16190 0 -1 16570
box -6 -8 86 248
use NAND3X1  _13146_
timestamp 0
transform -1 0 15490 0 1 16570
box -6 -8 106 248
use NAND3X1  _13147_
timestamp 0
transform -1 0 15870 0 -1 16570
box -6 -8 106 248
use NAND2X1  _13148_
timestamp 0
transform -1 0 16150 0 -1 16570
box -6 -8 86 248
use NAND3X1  _13149_
timestamp 0
transform 1 0 15910 0 -1 16570
box -6 -8 106 248
use NAND2X1  _13150_
timestamp 0
transform 1 0 13910 0 -1 17050
box -6 -8 86 248
use OAI21X1  _13151_
timestamp 0
transform -1 0 11970 0 -1 17050
box -6 -8 106 248
use NOR2X1  _13152_
timestamp 0
transform 1 0 12010 0 -1 17050
box -6 -8 86 248
use INVX1  _13153_
timestamp 0
transform -1 0 11830 0 -1 17050
box -6 -8 66 248
use AOI21X1  _13154_
timestamp 0
transform -1 0 11710 0 -1 17050
box -6 -8 106 248
use AOI22X1  _13155_
timestamp 0
transform 1 0 11450 0 -1 17050
box -6 -8 126 248
use OAI21X1  _13156_
timestamp 0
transform 1 0 13390 0 -1 17050
box -6 -8 106 248
use NOR2X1  _13157_
timestamp 0
transform -1 0 13610 0 -1 17050
box -6 -8 86 248
use AOI21X1  _13158_
timestamp 0
transform -1 0 13350 0 -1 17050
box -6 -8 106 248
use INVX1  _13159_
timestamp 0
transform -1 0 15170 0 1 16570
box -6 -8 66 248
use NAND3X1  _13160_
timestamp 0
transform -1 0 15950 0 1 16090
box -6 -8 106 248
use INVX1  _13161_
timestamp 0
transform -1 0 15930 0 1 15610
box -6 -8 66 248
use OAI21X1  _13162_
timestamp 0
transform -1 0 15830 0 -1 16090
box -6 -8 106 248
use INVX1  _13163_
timestamp 0
transform -1 0 15170 0 -1 16570
box -6 -8 66 248
use NAND3X1  _13164_
timestamp 0
transform 1 0 15210 0 -1 16570
box -6 -8 106 248
use OAI21X1  _13165_
timestamp 0
transform -1 0 15590 0 -1 16570
box -6 -8 106 248
use NAND2X1  _13166_
timestamp 0
transform 1 0 15350 0 -1 16570
box -6 -8 86 248
use AOI21X1  _13167_
timestamp 0
transform -1 0 15330 0 1 16570
box -6 -8 106 248
use NAND3X1  _13168_
timestamp 0
transform -1 0 15070 0 -1 16570
box -6 -8 106 248
use NAND2X1  _13169_
timestamp 0
transform -1 0 15070 0 1 16570
box -6 -8 86 248
use AOI21X1  _13170_
timestamp 0
transform -1 0 14950 0 1 16570
box -6 -8 106 248
use OAI21X1  _13171_
timestamp 0
transform -1 0 12630 0 -1 17050
box -6 -8 106 248
use INVX1  _13172_
timestamp 0
transform -1 0 11030 0 -1 17050
box -6 -8 66 248
use OR2X2  _13173_
timestamp 0
transform 1 0 12670 0 -1 17050
box -6 -8 106 248
use OAI21X1  _13174_
timestamp 0
transform -1 0 12390 0 -1 17050
box -6 -8 106 248
use OAI22X1  _13175_
timestamp 0
transform 1 0 10790 0 -1 17050
box -6 -8 126 248
use NAND2X1  _13176_
timestamp 0
transform -1 0 13390 0 -1 16570
box -6 -8 86 248
use NOR2X1  _13177_
timestamp 0
transform 1 0 12830 0 -1 17050
box -6 -8 86 248
use NOR2X1  _13178_
timestamp 0
transform -1 0 13930 0 1 16570
box -6 -8 86 248
use OAI21X1  _13179_
timestamp 0
transform -1 0 15370 0 -1 16090
box -6 -8 106 248
use INVX1  _13180_
timestamp 0
transform 1 0 15450 0 1 16090
box -6 -8 66 248
use OAI21X1  _13181_
timestamp 0
transform 1 0 15690 0 1 16090
box -6 -8 106 248
use NAND2X1  _13182_
timestamp 0
transform 1 0 15550 0 1 16090
box -6 -8 86 248
use OR2X2  _13183_
timestamp 0
transform -1 0 15410 0 1 16090
box -6 -8 106 248
use NAND3X1  _13184_
timestamp 0
transform -1 0 15150 0 1 16090
box -6 -8 106 248
use NAND2X1  _13185_
timestamp 0
transform 1 0 15190 0 1 16090
box -6 -8 86 248
use NAND2X1  _13186_
timestamp 0
transform 1 0 14850 0 -1 16570
box -6 -8 86 248
use NAND2X1  _13187_
timestamp 0
transform -1 0 14550 0 -1 16570
box -6 -8 86 248
use AND2X2  _13188_
timestamp 0
transform -1 0 13910 0 -1 16570
box -6 -8 106 248
use OAI21X1  _13189_
timestamp 0
transform 1 0 13970 0 -1 16570
box -6 -8 106 248
use OAI21X1  _13190_
timestamp 0
transform -1 0 13770 0 -1 16570
box -6 -8 106 248
use INVX1  _13191_
timestamp 0
transform -1 0 10250 0 -1 17050
box -6 -8 66 248
use INVX1  _13192_
timestamp 0
transform -1 0 14650 0 -1 16570
box -6 -8 66 248
use AOI21X1  _13193_
timestamp 0
transform -1 0 14670 0 1 16570
box -6 -8 106 248
use NOR2X1  _13194_
timestamp 0
transform 1 0 14710 0 1 16570
box -6 -8 86 248
use NAND3X1  _13195_
timestamp 0
transform -1 0 14790 0 -1 16570
box -6 -8 106 248
use OAI21X1  _13196_
timestamp 0
transform 1 0 14410 0 1 16570
box -6 -8 106 248
use OAI21X1  _13197_
timestamp 0
transform -1 0 15830 0 1 15610
box -6 -8 106 248
use INVX1  _13198_
timestamp 0
transform -1 0 15690 0 1 15610
box -6 -8 66 248
use OR2X2  _13199_
timestamp 0
transform -1 0 15510 0 -1 16090
box -6 -8 106 248
use OAI21X1  _13200_
timestamp 0
transform -1 0 15210 0 -1 16090
box -6 -8 106 248
use NAND2X1  _13201_
timestamp 0
transform 1 0 14910 0 1 16090
box -6 -8 86 248
use OR2X2  _13202_
timestamp 0
transform -1 0 14850 0 1 16090
box -6 -8 106 248
use NAND3X1  _13203_
timestamp 0
transform -1 0 14710 0 1 16090
box -6 -8 106 248
use AND2X2  _13204_
timestamp 0
transform -1 0 14930 0 -1 16090
box -6 -8 106 248
use NOR2X1  _13205_
timestamp 0
transform 1 0 14990 0 -1 16090
box -6 -8 86 248
use OAI21X1  _13206_
timestamp 0
transform -1 0 14790 0 -1 16090
box -6 -8 106 248
use NAND2X1  _13207_
timestamp 0
transform 1 0 14350 0 -1 16570
box -6 -8 86 248
use AND2X2  _13208_
timestamp 0
transform -1 0 14230 0 1 16570
box -6 -8 106 248
use NOR2X1  _13209_
timestamp 0
transform 1 0 14270 0 1 16570
box -6 -8 86 248
use NOR2X1  _13210_
timestamp 0
transform -1 0 14070 0 1 16570
box -6 -8 86 248
use AOI22X1  _13211_
timestamp 0
transform 1 0 10290 0 -1 17050
box -6 -8 126 248
use NAND2X1  _13212_
timestamp 0
transform -1 0 13130 0 1 16570
box -6 -8 86 248
use INVX1  _13213_
timestamp 0
transform -1 0 14310 0 -1 16570
box -6 -8 66 248
use AOI21X1  _13214_
timestamp 0
transform -1 0 14210 0 -1 16570
box -6 -8 106 248
use NAND2X1  _13215_
timestamp 0
transform -1 0 14550 0 1 16090
box -6 -8 86 248
use NOR2X1  _13216_
timestamp 0
transform 1 0 14330 0 1 16090
box -6 -8 86 248
use AOI21X1  _13217_
timestamp 0
transform -1 0 14290 0 1 16090
box -6 -8 106 248
use NOR2X1  _13218_
timestamp 0
transform -1 0 14130 0 1 16090
box -6 -8 86 248
use AND2X2  _13219_
timestamp 0
transform -1 0 13810 0 1 16570
box -6 -8 106 248
use OAI21X1  _13220_
timestamp 0
transform -1 0 13670 0 1 16570
box -6 -8 106 248
use OAI21X1  _13221_
timestamp 0
transform -1 0 13510 0 1 16570
box -6 -8 106 248
use OAI21X1  _13222_
timestamp 0
transform -1 0 13470 0 1 12250
box -6 -8 106 248
use OAI21X1  _13223_
timestamp 0
transform -1 0 13370 0 -1 12730
box -6 -8 106 248
use INVX1  _13224_
timestamp 0
transform -1 0 12830 0 1 12730
box -6 -8 66 248
use NAND2X1  _13225_
timestamp 0
transform 1 0 11610 0 1 13210
box -6 -8 86 248
use INVX1  _13226_
timestamp 0
transform -1 0 13290 0 -1 13210
box -6 -8 66 248
use NOR2X1  _13227_
timestamp 0
transform -1 0 13170 0 1 12250
box -6 -8 86 248
use AOI21X1  _13228_
timestamp 0
transform 1 0 13350 0 -1 12250
box -6 -8 106 248
use NOR2X1  _13229_
timestamp 0
transform -1 0 13750 0 -1 12730
box -6 -8 86 248
use OAI21X1  _13230_
timestamp 0
transform -1 0 13310 0 1 12250
box -6 -8 106 248
use AND2X2  _13231_
timestamp 0
transform -1 0 13030 0 1 12250
box -6 -8 106 248
use OR2X2  _13232_
timestamp 0
transform -1 0 11730 0 -1 12730
box -6 -8 106 248
use OR2X2  _13233_
timestamp 0
transform 1 0 11210 0 -1 12730
box -6 -8 106 248
use OAI21X1  _13234_
timestamp 0
transform -1 0 11590 0 -1 12730
box -6 -8 106 248
use NAND2X1  _13235_
timestamp 0
transform -1 0 11430 0 -1 12730
box -6 -8 86 248
use NOR2X1  _13236_
timestamp 0
transform -1 0 11510 0 -1 13210
box -6 -8 86 248
use NAND2X1  _13237_
timestamp 0
transform -1 0 11370 0 -1 13210
box -6 -8 86 248
use NAND2X1  _13238_
timestamp 0
transform -1 0 11250 0 -1 13210
box -6 -8 86 248
use OAI21X1  _13239_
timestamp 0
transform 1 0 11570 0 -1 13210
box -6 -8 106 248
use INVX1  _13240_
timestamp 0
transform -1 0 11050 0 -1 12730
box -6 -8 66 248
use OAI21X1  _13241_
timestamp 0
transform 1 0 10990 0 1 12730
box -6 -8 106 248
use OAI21X1  _13242_
timestamp 0
transform -1 0 13890 0 -1 12730
box -6 -8 106 248
use OAI21X1  _13243_
timestamp 0
transform 1 0 11790 0 -1 12730
box -6 -8 106 248
use MUX2X1  _13244_
timestamp 0
transform -1 0 12050 0 -1 12730
box -6 -8 126 248
use NAND2X1  _13245_
timestamp 0
transform -1 0 11370 0 1 12730
box -6 -8 86 248
use OR2X2  _13246_
timestamp 0
transform -1 0 11250 0 1 12730
box -6 -8 106 248
use NAND2X1  _13247_
timestamp 0
transform 1 0 10550 0 1 12730
box -6 -8 86 248
use INVX1  _13248_
timestamp 0
transform -1 0 10510 0 1 12730
box -6 -8 66 248
use NAND2X1  _13249_
timestamp 0
transform -1 0 10390 0 1 12730
box -6 -8 86 248
use NOR2X1  _13250_
timestamp 0
transform 1 0 11250 0 1 13210
box -6 -8 86 248
use NAND2X1  _13251_
timestamp 0
transform -1 0 10270 0 1 12730
box -6 -8 86 248
use INVX1  _13252_
timestamp 0
transform -1 0 10130 0 1 12730
box -6 -8 66 248
use INVX1  _13253_
timestamp 0
transform -1 0 12170 0 -1 12730
box -6 -8 66 248
use NOR2X1  _13254_
timestamp 0
transform 1 0 14510 0 1 12250
box -6 -8 86 248
use OAI21X1  _13255_
timestamp 0
transform -1 0 14470 0 1 12250
box -6 -8 106 248
use OAI21X1  _13256_
timestamp 0
transform 1 0 13430 0 -1 13210
box -6 -8 106 248
use OAI21X1  _13257_
timestamp 0
transform 1 0 13510 0 1 12250
box -6 -8 106 248
use NOR2X1  _13258_
timestamp 0
transform -1 0 11270 0 1 12250
box -6 -8 86 248
use NAND2X1  _13259_
timestamp 0
transform 1 0 11310 0 1 12250
box -6 -8 86 248
use INVX1  _13260_
timestamp 0
transform -1 0 10970 0 1 12250
box -6 -8 66 248
use NOR2X1  _13261_
timestamp 0
transform -1 0 10850 0 1 12250
box -6 -8 86 248
use OAI21X1  _13262_
timestamp 0
transform -1 0 10710 0 -1 12730
box -6 -8 106 248
use AOI21X1  _13263_
timestamp 0
transform 1 0 10670 0 1 12730
box -6 -8 106 248
use NOR2X1  _13264_
timestamp 0
transform -1 0 11130 0 -1 13210
box -6 -8 86 248
use INVX1  _13265_
timestamp 0
transform -1 0 12110 0 -1 11770
box -6 -8 66 248
use AOI21X1  _13266_
timestamp 0
transform 1 0 13870 0 -1 12250
box -6 -8 106 248
use OAI21X1  _13267_
timestamp 0
transform -1 0 14130 0 -1 12250
box -6 -8 106 248
use OAI21X1  _13268_
timestamp 0
transform 1 0 13730 0 -1 12250
box -6 -8 106 248
use OR2X2  _13269_
timestamp 0
transform -1 0 11990 0 -1 11770
box -6 -8 106 248
use NAND2X1  _13270_
timestamp 0
transform 1 0 12070 0 1 11770
box -6 -8 86 248
use NAND2X1  _13271_
timestamp 0
transform -1 0 11870 0 1 11770
box -6 -8 86 248
use AOI21X1  _13272_
timestamp 0
transform 1 0 11030 0 1 12250
box -6 -8 106 248
use OAI21X1  _13273_
timestamp 0
transform -1 0 11350 0 1 11770
box -6 -8 106 248
use INVX1  _13274_
timestamp 0
transform 1 0 13470 0 1 11770
box -6 -8 66 248
use OAI21X1  _13275_
timestamp 0
transform -1 0 14030 0 -1 12730
box -6 -8 106 248
use OAI21X1  _13276_
timestamp 0
transform 1 0 13930 0 1 12250
box -6 -8 106 248
use OR2X2  _13277_
timestamp 0
transform -1 0 13890 0 1 12250
box -6 -8 106 248
use NAND2X1  _13278_
timestamp 0
transform -1 0 13730 0 1 12250
box -6 -8 86 248
use OR2X2  _13279_
timestamp 0
transform -1 0 12510 0 -1 11770
box -6 -8 106 248
use NAND2X1  _13280_
timestamp 0
transform 1 0 12550 0 -1 11770
box -6 -8 86 248
use NAND2X1  _13281_
timestamp 0
transform 1 0 11770 0 -1 11770
box -6 -8 86 248
use INVX1  _13282_
timestamp 0
transform -1 0 11570 0 -1 11770
box -6 -8 66 248
use NOR2X1  _13283_
timestamp 0
transform 1 0 11130 0 1 11770
box -6 -8 86 248
use NAND2X1  _13284_
timestamp 0
transform -1 0 10830 0 -1 11770
box -6 -8 86 248
use NAND2X1  _13285_
timestamp 0
transform 1 0 10610 0 -1 11770
box -6 -8 86 248
use OAI22X1  _13286_
timestamp 0
transform 1 0 10970 0 1 11770
box -6 -8 126 248
use INVX1  _13287_
timestamp 0
transform -1 0 11450 0 1 11770
box -6 -8 66 248
use NAND2X1  _13288_
timestamp 0
transform 1 0 10870 0 -1 11770
box -6 -8 86 248
use OAI21X1  _13289_
timestamp 0
transform 1 0 11630 0 -1 11770
box -6 -8 106 248
use INVX1  _13290_
timestamp 0
transform -1 0 11210 0 -1 11770
box -6 -8 66 248
use OAI21X1  _13291_
timestamp 0
transform 1 0 11010 0 -1 11770
box -6 -8 106 248
use OAI21X1  _13292_
timestamp 0
transform -1 0 14730 0 1 12250
box -6 -8 106 248
use NOR2X1  _13293_
timestamp 0
transform 1 0 14450 0 -1 12250
box -6 -8 86 248
use NAND2X1  _13294_
timestamp 0
transform 1 0 14310 0 -1 12250
box -6 -8 86 248
use OAI21X1  _13295_
timestamp 0
transform -1 0 14310 0 1 12250
box -6 -8 106 248
use NAND2X1  _13296_
timestamp 0
transform -1 0 14270 0 -1 12250
box -6 -8 86 248
use NAND2X1  _13297_
timestamp 0
transform 1 0 12450 0 -1 12250
box -6 -8 86 248
use OR2X2  _13298_
timestamp 0
transform -1 0 12410 0 -1 12250
box -6 -8 106 248
use NAND2X1  _13299_
timestamp 0
transform 1 0 12190 0 1 11770
box -6 -8 86 248
use INVX1  _13300_
timestamp 0
transform -1 0 11450 0 -1 11770
box -6 -8 66 248
use NAND2X1  _13301_
timestamp 0
transform -1 0 11350 0 -1 11770
box -6 -8 86 248
use INVX1  _13302_
timestamp 0
transform -1 0 11510 0 -1 12250
box -6 -8 66 248
use NAND2X1  _13303_
timestamp 0
transform -1 0 12250 0 -1 12250
box -6 -8 86 248
use INVX1  _13304_
timestamp 0
transform 1 0 12570 0 -1 12250
box -6 -8 66 248
use NAND2X1  _13305_
timestamp 0
transform -1 0 13310 0 -1 12250
box -6 -8 86 248
use OR2X2  _13306_
timestamp 0
transform -1 0 13170 0 -1 12250
box -6 -8 106 248
use NAND2X1  _13307_
timestamp 0
transform -1 0 13030 0 -1 12250
box -6 -8 86 248
use NOR2X1  _13308_
timestamp 0
transform 1 0 12830 0 -1 12250
box -6 -8 86 248
use INVX1  _13309_
timestamp 0
transform 1 0 12850 0 1 11770
box -6 -8 66 248
use NAND2X1  _13310_
timestamp 0
transform 1 0 12690 0 -1 12250
box -6 -8 86 248
use NAND2X1  _13311_
timestamp 0
transform 1 0 12730 0 1 11770
box -6 -8 86 248
use OR2X2  _13312_
timestamp 0
transform 1 0 12010 0 -1 12250
box -6 -8 106 248
use AOI21X1  _13313_
timestamp 0
transform -1 0 11970 0 -1 12250
box -6 -8 106 248
use AOI22X1  _13314_
timestamp 0
transform 1 0 11690 0 -1 12250
box -6 -8 126 248
use NOR2X1  _13315_
timestamp 0
transform 1 0 13110 0 -1 13210
box -6 -8 86 248
use INVX1  _13316_
timestamp 0
transform -1 0 12830 0 -1 13210
box -6 -8 66 248
use NAND3X1  _13317_
timestamp 0
transform -1 0 12730 0 -1 13210
box -6 -8 106 248
use INVX1  _13318_
timestamp 0
transform 1 0 12230 0 -1 13210
box -6 -8 66 248
use AOI21X1  _13319_
timestamp 0
transform -1 0 12570 0 -1 13210
box -6 -8 106 248
use NOR2X1  _13320_
timestamp 0
transform -1 0 12430 0 -1 13210
box -6 -8 86 248
use OAI21X1  _13321_
timestamp 0
transform 1 0 12310 0 1 11770
box -6 -8 106 248
use NOR2X1  _13322_
timestamp 0
transform 1 0 11930 0 1 11770
box -6 -8 86 248
use AOI21X1  _13323_
timestamp 0
transform 1 0 11650 0 1 11770
box -6 -8 106 248
use NAND3X1  _13324_
timestamp 0
transform 1 0 11510 0 1 11770
box -6 -8 106 248
use OAI21X1  _13325_
timestamp 0
transform 1 0 11550 0 -1 12250
box -6 -8 106 248
use AOI21X1  _13326_
timestamp 0
transform 1 0 11710 0 -1 13210
box -6 -8 106 248
use OR2X2  _13327_
timestamp 0
transform -1 0 12210 0 -1 13690
box -6 -8 106 248
use NAND2X1  _13328_
timestamp 0
transform 1 0 12250 0 -1 13690
box -6 -8 86 248
use NAND2X1  _13329_
timestamp 0
transform 1 0 11970 0 -1 13690
box -6 -8 86 248
use AND2X2  _13330_
timestamp 0
transform -1 0 11830 0 1 13210
box -6 -8 106 248
use OAI21X1  _13331_
timestamp 0
transform 1 0 11810 0 -1 13690
box -6 -8 106 248
use OAI22X1  _13332_
timestamp 0
transform 1 0 11650 0 -1 13690
box -6 -8 126 248
use OAI21X1  _13333_
timestamp 0
transform 1 0 11870 0 1 13210
box -6 -8 106 248
use NAND3X1  _13334_
timestamp 0
transform 1 0 12030 0 1 13210
box -6 -8 106 248
use INVX1  _13335_
timestamp 0
transform -1 0 12070 0 -1 13210
box -6 -8 66 248
use AOI21X1  _13336_
timestamp 0
transform 1 0 11870 0 -1 13210
box -6 -8 106 248
use INVX1  _13337_
timestamp 0
transform 1 0 12990 0 -1 13210
box -6 -8 66 248
use NAND2X1  _13338_
timestamp 0
transform -1 0 12950 0 -1 13210
box -6 -8 86 248
use NAND2X1  _13339_
timestamp 0
transform 1 0 12990 0 1 13210
box -6 -8 86 248
use NAND2X1  _13340_
timestamp 0
transform -1 0 12930 0 1 13210
box -6 -8 86 248
use NAND2X1  _13341_
timestamp 0
transform -1 0 11730 0 -1 14170
box -6 -8 86 248
use OAI21X1  _13342_
timestamp 0
transform -1 0 12270 0 1 13210
box -6 -8 106 248
use OAI21X1  _13343_
timestamp 0
transform -1 0 11910 0 1 13690
box -6 -8 106 248
use NAND2X1  _13344_
timestamp 0
transform 1 0 11970 0 1 14170
box -6 -8 86 248
use NAND2X1  _13345_
timestamp 0
transform 1 0 12230 0 1 14170
box -6 -8 86 248
use NOR2X1  _13346_
timestamp 0
transform 1 0 12110 0 1 14170
box -6 -8 86 248
use NAND2X1  _13347_
timestamp 0
transform -1 0 14790 0 1 12730
box -6 -8 86 248
use OAI21X1  _13348_
timestamp 0
transform 1 0 14970 0 -1 14170
box -6 -8 106 248
use NAND2X1  _13349_
timestamp 0
transform -1 0 15170 0 -1 13690
box -6 -8 86 248
use OAI21X1  _13350_
timestamp 0
transform -1 0 15290 0 -1 14650
box -6 -8 106 248
use INVX1  _13351_
timestamp 0
transform 1 0 15050 0 1 12250
box -6 -8 66 248
use OR2X2  _13352_
timestamp 0
transform 1 0 14750 0 1 13210
box -6 -8 106 248
use OAI21X1  _13353_
timestamp 0
transform 1 0 14910 0 1 13210
box -6 -8 106 248
use OAI21X1  _13354_
timestamp 0
transform -1 0 15090 0 -1 13210
box -6 -8 106 248
use INVX1  _13355_
timestamp 0
transform -1 0 15210 0 -1 13210
box -6 -8 66 248
use OAI21X1  _13356_
timestamp 0
transform 1 0 15050 0 1 13210
box -6 -8 106 248
use OAI21X1  _13357_
timestamp 0
transform 1 0 15190 0 1 13210
box -6 -8 106 248
use NAND2X1  _13358_
timestamp 0
transform -1 0 11750 0 1 13690
box -6 -8 86 248
use NAND2X1  _13359_
timestamp 0
transform -1 0 15390 0 1 12250
box -6 -8 86 248
use OAI21X1  _13360_
timestamp 0
transform 1 0 15170 0 1 12250
box -6 -8 106 248
use NAND2X1  _13361_
timestamp 0
transform -1 0 15350 0 1 12730
box -6 -8 86 248
use OAI21X1  _13362_
timestamp 0
transform 1 0 15130 0 1 12730
box -6 -8 106 248
use AND2X2  _13363_
timestamp 0
transform 1 0 12370 0 1 14170
box -6 -8 106 248
use NAND2X1  _13364_
timestamp 0
transform 1 0 16590 0 1 12250
box -6 -8 86 248
use OAI21X1  _13365_
timestamp 0
transform -1 0 16950 0 1 12250
box -6 -8 106 248
use NAND2X1  _13366_
timestamp 0
transform 1 0 16830 0 -1 12730
box -6 -8 86 248
use OAI21X1  _13367_
timestamp 0
transform 1 0 16810 0 1 12730
box -6 -8 106 248
use OAI21X1  _13368_
timestamp 0
transform 1 0 15270 0 -1 12730
box -6 -8 106 248
use OAI21X1  _13369_
timestamp 0
transform 1 0 15130 0 -1 12730
box -6 -8 106 248
use OAI21X1  _13370_
timestamp 0
transform 1 0 14850 0 1 12730
box -6 -8 106 248
use OAI21X1  _13371_
timestamp 0
transform -1 0 15090 0 1 12730
box -6 -8 106 248
use NAND2X1  _13372_
timestamp 0
transform -1 0 15770 0 1 12250
box -6 -8 86 248
use OAI21X1  _13373_
timestamp 0
transform -1 0 15910 0 1 12250
box -6 -8 106 248
use NAND2X1  _13374_
timestamp 0
transform -1 0 16170 0 1 12250
box -6 -8 86 248
use OAI21X1  _13375_
timestamp 0
transform 1 0 16210 0 1 12250
box -6 -8 106 248
use NAND2X1  _13376_
timestamp 0
transform 1 0 14130 0 -1 14650
box -6 -8 86 248
use OAI21X1  _13377_
timestamp 0
transform -1 0 14370 0 -1 14650
box -6 -8 106 248
use NAND2X1  _13378_
timestamp 0
transform -1 0 14750 0 -1 14650
box -6 -8 86 248
use OAI21X1  _13379_
timestamp 0
transform -1 0 14910 0 -1 14650
box -6 -8 106 248
use INVX1  _13380_
timestamp 0
transform 1 0 14070 0 1 12730
box -6 -8 66 248
use OAI21X1  _13381_
timestamp 0
transform 1 0 14950 0 -1 13690
box -6 -8 106 248
use OAI21X1  _13382_
timestamp 0
transform 1 0 14810 0 -1 13690
box -6 -8 106 248
use INVX1  _13383_
timestamp 0
transform 1 0 14270 0 -1 13210
box -6 -8 66 248
use OAI21X1  _13384_
timestamp 0
transform 1 0 14350 0 1 13690
box -6 -8 106 248
use OAI21X1  _13385_
timestamp 0
transform 1 0 14410 0 -1 13690
box -6 -8 106 248
use NAND2X1  _13386_
timestamp 0
transform -1 0 13930 0 1 13690
box -6 -8 86 248
use OAI21X1  _13387_
timestamp 0
transform -1 0 13970 0 -1 13690
box -6 -8 106 248
use NAND2X1  _13388_
timestamp 0
transform -1 0 14050 0 1 13690
box -6 -8 86 248
use OAI21X1  _13389_
timestamp 0
transform -1 0 14370 0 -1 13690
box -6 -8 106 248
use NAND2X1  _13390_
timestamp 0
transform 1 0 14190 0 -1 14170
box -6 -8 86 248
use OAI21X1  _13391_
timestamp 0
transform 1 0 14330 0 -1 14170
box -6 -8 106 248
use NAND2X1  _13392_
timestamp 0
transform -1 0 14710 0 1 14170
box -6 -8 86 248
use OAI21X1  _13393_
timestamp 0
transform 1 0 14490 0 1 14170
box -6 -8 106 248
use OAI21X1  _13394_
timestamp 0
transform -1 0 13650 0 1 12730
box -6 -8 106 248
use OAI21X1  _13395_
timestamp 0
transform -1 0 13790 0 1 12730
box -6 -8 106 248
use OAI21X1  _13396_
timestamp 0
transform 1 0 14570 0 1 12730
box -6 -8 106 248
use OAI21X1  _13397_
timestamp 0
transform 1 0 14370 0 -1 13210
box -6 -8 106 248
use NAND2X1  _13398_
timestamp 0
transform 1 0 13030 0 1 12730
box -6 -8 86 248
use OAI21X1  _13399_
timestamp 0
transform -1 0 13250 0 1 12730
box -6 -8 106 248
use NAND2X1  _13400_
timestamp 0
transform -1 0 14930 0 -1 12730
box -6 -8 86 248
use OAI21X1  _13401_
timestamp 0
transform -1 0 15090 0 -1 12730
box -6 -8 106 248
use NAND2X1  _13402_
timestamp 0
transform -1 0 12030 0 1 12730
box -6 -8 86 248
use OAI21X1  _13403_
timestamp 0
transform -1 0 12190 0 1 12730
box -6 -8 106 248
use NAND2X1  _13404_
timestamp 0
transform 1 0 12990 0 -1 12730
box -6 -8 86 248
use OAI21X1  _13405_
timestamp 0
transform -1 0 13230 0 -1 12730
box -6 -8 106 248
use INVX1  _13406_
timestamp 0
transform -1 0 12010 0 1 12250
box -6 -8 66 248
use OAI21X1  _13407_
timestamp 0
transform -1 0 12810 0 1 13210
box -6 -8 106 248
use OAI21X1  _13408_
timestamp 0
transform 1 0 12570 0 1 13210
box -6 -8 106 248
use INVX1  _13409_
timestamp 0
transform -1 0 12630 0 1 12250
box -6 -8 66 248
use OAI21X1  _13410_
timestamp 0
transform -1 0 12870 0 -1 13690
box -6 -8 106 248
use OAI21X1  _13411_
timestamp 0
transform 1 0 12610 0 -1 13690
box -6 -8 106 248
use NAND2X1  _13412_
timestamp 0
transform -1 0 11750 0 1 12250
box -6 -8 86 248
use OAI21X1  _13413_
timestamp 0
transform -1 0 11910 0 1 12250
box -6 -8 106 248
use NAND2X1  _13414_
timestamp 0
transform 1 0 12450 0 1 12250
box -6 -8 86 248
use OAI21X1  _13415_
timestamp 0
transform -1 0 12410 0 1 12250
box -6 -8 106 248
use NAND2X1  _13416_
timestamp 0
transform 1 0 12610 0 1 11770
box -6 -8 86 248
use OAI21X1  _13417_
timestamp 0
transform 1 0 12470 0 1 11770
box -6 -8 106 248
use NAND2X1  _13418_
timestamp 0
transform 1 0 12950 0 1 11770
box -6 -8 86 248
use OAI21X1  _13419_
timestamp 0
transform -1 0 13170 0 1 11770
box -6 -8 106 248
use OAI21X1  _13420_
timestamp 0
transform -1 0 11770 0 1 12730
box -6 -8 106 248
use OAI21X1  _13421_
timestamp 0
transform -1 0 11910 0 1 12730
box -6 -8 106 248
use OAI21X1  _13422_
timestamp 0
transform -1 0 12330 0 -1 12730
box -6 -8 106 248
use OAI21X1  _13423_
timestamp 0
transform -1 0 12470 0 -1 12730
box -6 -8 106 248
use NAND2X1  _13424_
timestamp 0
transform -1 0 12550 0 1 12730
box -6 -8 86 248
use OAI21X1  _13425_
timestamp 0
transform -1 0 12710 0 1 12730
box -6 -8 106 248
use NAND2X1  _13426_
timestamp 0
transform 1 0 11090 0 -1 12730
box -6 -8 86 248
use OAI21X1  _13427_
timestamp 0
transform -1 0 10930 0 1 12730
box -6 -8 106 248
use DFFPOSX1  _13428_
timestamp 0
transform -1 0 12330 0 -1 14170
box -6 -8 246 248
use DFFPOSX1  _13429_
timestamp 0
transform 1 0 11090 0 -1 14650
box -6 -8 246 248
use DFFPOSX1  _13430_
timestamp 0
transform -1 0 9730 0 -1 10810
box -6 -8 246 248
use DFFPOSX1  _13431_
timestamp 0
transform -1 0 12050 0 -1 15130
box -6 -8 246 248
use DFFPOSX1  _13432_
timestamp 0
transform -1 0 11790 0 1 14650
box -6 -8 246 248
use DFFPOSX1  _13433_
timestamp 0
transform -1 0 11950 0 1 15130
box -6 -8 246 248
use DFFPOSX1  _13434_
timestamp 0
transform -1 0 11470 0 -1 15610
box -6 -8 246 248
use DFFPOSX1  _13435_
timestamp 0
transform -1 0 12130 0 -1 15610
box -6 -8 246 248
use DFFPOSX1  _13436_
timestamp 0
transform -1 0 11850 0 1 15610
box -6 -8 246 248
use DFFPOSX1  _13437_
timestamp 0
transform -1 0 11750 0 -1 16090
box -6 -8 246 248
use DFFPOSX1  _13438_
timestamp 0
transform 1 0 10690 0 1 16570
box -6 -8 246 248
use DFFPOSX1  _13439_
timestamp 0
transform -1 0 11910 0 -1 16570
box -6 -8 246 248
use DFFPOSX1  _13440_
timestamp 0
transform -1 0 11670 0 -1 16570
box -6 -8 246 248
use DFFPOSX1  _13441_
timestamp 0
transform -1 0 14830 0 1 14650
box -6 -8 246 248
use DFFPOSX1  _13442_
timestamp 0
transform -1 0 12330 0 -1 14650
box -6 -8 246 248
use DFFPOSX1  _13443_
timestamp 0
transform -1 0 12730 0 1 14650
box -6 -8 246 248
use DFFPOSX1  _13444_
timestamp 0
transform -1 0 12830 0 1 14170
box -6 -8 246 248
use DFFPOSX1  _13445_
timestamp 0
transform -1 0 11790 0 1 16570
box -6 -8 246 248
use DFFPOSX1  _13446_
timestamp 0
transform -1 0 12570 0 1 16570
box -6 -8 246 248
use DFFPOSX1  _13447_
timestamp 0
transform 1 0 9270 0 -1 17050
box -6 -8 246 248
use DFFPOSX1  _13448_
timestamp 0
transform 1 0 11030 0 -1 17050
box -6 -8 246 248
use DFFPOSX1  _13449_
timestamp 0
transform -1 0 10750 0 -1 17050
box -6 -8 246 248
use DFFPOSX1  _13450_
timestamp 0
transform -1 0 13630 0 -1 16570
box -6 -8 246 248
use DFFPOSX1  _13451_
timestamp 0
transform 1 0 9890 0 -1 17050
box -6 -8 246 248
use DFFPOSX1  _13452_
timestamp 0
transform -1 0 13370 0 1 16570
box -6 -8 246 248
use DFFPOSX1  _13453_
timestamp 0
transform -1 0 11570 0 1 13210
box -6 -8 246 248
use DFFPOSX1  _13454_
timestamp 0
transform 1 0 10970 0 1 13210
box -6 -8 246 248
use DFFPOSX1  _13455_
timestamp 0
transform -1 0 10910 0 1 11770
box -6 -8 246 248
use DFFPOSX1  _13456_
timestamp 0
transform 1 0 11170 0 -1 12250
box -6 -8 246 248
use DFFPOSX1  _13457_
timestamp 0
transform 1 0 11350 0 -1 13690
box -6 -8 246 248
use DFFPOSX1  _13458_
timestamp 0
transform -1 0 11970 0 -1 14170
box -6 -8 246 248
use DFFPOSX1  _13459_
timestamp 0
transform 1 0 14970 0 1 14170
box -6 -8 246 248
use DFFPOSX1  _13460_
timestamp 0
transform 1 0 14910 0 -1 14650
box -6 -8 246 248
use DFFPOSX1  _13461_
timestamp 0
transform 1 0 14710 0 -1 13210
box -6 -8 246 248
use DFFPOSX1  _13462_
timestamp 0
transform 1 0 15290 0 1 13210
box -6 -8 246 248
use DFFPOSX1  _13463_
timestamp 0
transform 1 0 15390 0 1 12250
box -6 -8 246 248
use DFFPOSX1  _13464_
timestamp 0
transform 1 0 15350 0 1 12730
box -6 -8 246 248
use DFFPOSX1  _13465_
timestamp 0
transform 1 0 16910 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _13466_
timestamp 0
transform 1 0 16910 0 1 12730
box -6 -8 246 248
use DFFPOSX1  _13467_
timestamp 0
transform 1 0 15610 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _13468_
timestamp 0
transform 1 0 15370 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _13469_
timestamp 0
transform -1 0 16150 0 -1 12250
box -6 -8 246 248
use DFFPOSX1  _13470_
timestamp 0
transform 1 0 16310 0 1 12250
box -6 -8 246 248
use DFFPOSX1  _13471_
timestamp 0
transform 1 0 14190 0 1 14650
box -6 -8 246 248
use DFFPOSX1  _13472_
timestamp 0
transform 1 0 14830 0 1 14650
box -6 -8 246 248
use DFFPOSX1  _13473_
timestamp 0
transform -1 0 14750 0 -1 13690
box -6 -8 246 248
use DFFPOSX1  _13474_
timestamp 0
transform -1 0 14690 0 1 13690
box -6 -8 246 248
use DFFPOSX1  _13475_
timestamp 0
transform 1 0 13970 0 -1 13690
box -6 -8 246 248
use DFFPOSX1  _13476_
timestamp 0
transform -1 0 14290 0 1 13690
box -6 -8 246 248
use DFFPOSX1  _13477_
timestamp 0
transform 1 0 14670 0 -1 14170
box -6 -8 246 248
use DFFPOSX1  _13478_
timestamp 0
transform 1 0 14430 0 -1 14170
box -6 -8 246 248
use DFFPOSX1  _13479_
timestamp 0
transform 1 0 13790 0 1 12730
box -6 -8 246 248
use DFFPOSX1  _13480_
timestamp 0
transform 1 0 14470 0 -1 13210
box -6 -8 246 248
use DFFPOSX1  _13481_
timestamp 0
transform 1 0 13250 0 1 12730
box -6 -8 246 248
use DFFPOSX1  _13482_
timestamp 0
transform -1 0 14810 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _13483_
timestamp 0
transform 1 0 12190 0 1 12730
box -6 -8 246 248
use DFFPOSX1  _13484_
timestamp 0
transform 1 0 13370 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _13485_
timestamp 0
transform 1 0 12270 0 1 13210
box -6 -8 246 248
use DFFPOSX1  _13486_
timestamp 0
transform -1 0 12570 0 -1 13690
box -6 -8 246 248
use DFFPOSX1  _13487_
timestamp 0
transform 1 0 11390 0 1 12250
box -6 -8 246 248
use DFFPOSX1  _13488_
timestamp 0
transform 1 0 12010 0 1 12250
box -6 -8 246 248
use DFFPOSX1  _13489_
timestamp 0
transform -1 0 12350 0 -1 11770
box -6 -8 246 248
use DFFPOSX1  _13490_
timestamp 0
transform 1 0 13170 0 1 11770
box -6 -8 246 248
use DFFPOSX1  _13491_
timestamp 0
transform -1 0 11610 0 1 12730
box -6 -8 246 248
use DFFPOSX1  _13492_
timestamp 0
transform -1 0 12710 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _13493_
timestamp 0
transform 1 0 12710 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _13494_
timestamp 0
transform 1 0 10710 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _13495_
timestamp 0
transform -1 0 12870 0 1 12250
box -6 -8 246 248
use DFFPOSX1  _13496_
timestamp 0
transform -1 0 11510 0 1 14170
box -6 -8 246 248
use DFFPOSX1  _13497_
timestamp 0
transform 1 0 11030 0 1 14170
box -6 -8 246 248
use DFFPOSX1  _13498_
timestamp 0
transform 1 0 10630 0 -1 16090
box -6 -8 246 248
use DFFPOSX1  _13499_
timestamp 0
transform 1 0 10870 0 -1 16090
box -6 -8 246 248
use DFFPOSX1  _13500_
timestamp 0
transform -1 0 11390 0 1 14650
box -6 -8 246 248
use DFFPOSX1  _13501_
timestamp 0
transform -1 0 11090 0 -1 14650
box -6 -8 246 248
use INVX2  _13502_
timestamp 0
transform -1 0 7710 0 -1 12730
box -6 -8 66 248
use NOR2X1  _13503_
timestamp 0
transform -1 0 7610 0 -1 12730
box -6 -8 86 248
use INVX2  _13504_
timestamp 0
transform -1 0 7850 0 1 12730
box -6 -8 66 248
use INVX2  _13505_
timestamp 0
transform 1 0 7970 0 -1 11770
box -6 -8 66 248
use NOR2X1  _13506_
timestamp 0
transform 1 0 8390 0 1 11770
box -6 -8 86 248
use INVX1  _13507_
timestamp 0
transform 1 0 8610 0 -1 12250
box -6 -8 66 248
use AND2X2  _13508_
timestamp 0
transform 1 0 8470 0 -1 12250
box -6 -8 106 248
use NOR2X1  _13509_
timestamp 0
transform -1 0 7830 0 1 12250
box -6 -8 86 248
use INVX1  _13510_
timestamp 0
transform -1 0 7230 0 -1 12730
box -6 -8 66 248
use OAI21X1  _13511_
timestamp 0
transform 1 0 7210 0 1 12250
box -6 -8 106 248
use AOI21X1  _13512_
timestamp 0
transform -1 0 7170 0 1 12250
box -6 -8 106 248
use INVX1  _13513_
timestamp 0
transform 1 0 6410 0 -1 13210
box -6 -8 66 248
use NAND2X1  _13514_
timestamp 0
transform 1 0 7430 0 -1 12250
box -6 -8 86 248
use OAI21X1  _13515_
timestamp 0
transform -1 0 7790 0 -1 12250
box -6 -8 106 248
use OAI21X1  _13516_
timestamp 0
transform 1 0 7830 0 -1 12250
box -6 -8 106 248
use AOI22X1  _13517_
timestamp 0
transform -1 0 7270 0 -1 13210
box -6 -8 126 248
use NAND2X1  _13518_
timestamp 0
transform 1 0 7970 0 1 11770
box -6 -8 86 248
use INVX1  _13519_
timestamp 0
transform 1 0 7570 0 -1 11770
box -6 -8 66 248
use OAI21X1  _13520_
timestamp 0
transform 1 0 8110 0 1 11770
box -6 -8 106 248
use AOI21X1  _13521_
timestamp 0
transform -1 0 7930 0 -1 11770
box -6 -8 106 248
use INVX1  _13522_
timestamp 0
transform 1 0 7850 0 1 11770
box -6 -8 66 248
use NAND2X1  _13523_
timestamp 0
transform 1 0 7550 0 -1 12250
box -6 -8 86 248
use OAI21X1  _13524_
timestamp 0
transform -1 0 7790 0 1 11770
box -6 -8 106 248
use OAI21X1  _13525_
timestamp 0
transform -1 0 7790 0 -1 11770
box -6 -8 106 248
use AOI22X1  _13526_
timestamp 0
transform -1 0 7110 0 -1 12730
box -6 -8 126 248
use NAND2X1  _13527_
timestamp 0
transform 1 0 7610 0 1 11290
box -6 -8 86 248
use INVX1  _13528_
timestamp 0
transform -1 0 10170 0 -1 12250
box -6 -8 66 248
use OAI21X1  _13529_
timestamp 0
transform 1 0 9070 0 1 11770
box -6 -8 106 248
use AOI21X1  _13530_
timestamp 0
transform -1 0 9030 0 1 11770
box -6 -8 106 248
use INVX1  _13531_
timestamp 0
transform -1 0 9550 0 -1 12250
box -6 -8 66 248
use NAND2X1  _13532_
timestamp 0
transform -1 0 8830 0 1 12250
box -6 -8 86 248
use OAI21X1  _13533_
timestamp 0
transform 1 0 8710 0 -1 12250
box -6 -8 106 248
use OAI21X1  _13534_
timestamp 0
transform -1 0 8870 0 1 11770
box -6 -8 106 248
use AOI22X1  _13535_
timestamp 0
transform -1 0 8010 0 1 12730
box -6 -8 126 248
use NAND2X1  _13536_
timestamp 0
transform 1 0 8250 0 1 11770
box -6 -8 86 248
use INVX1  _13537_
timestamp 0
transform 1 0 8710 0 -1 12730
box -6 -8 66 248
use NOR2X1  _13538_
timestamp 0
transform 1 0 8930 0 -1 11770
box -6 -8 86 248
use OAI21X1  _13539_
timestamp 0
transform -1 0 9330 0 1 11770
box -6 -8 106 248
use AOI22X1  _13540_
timestamp 0
transform -1 0 8690 0 1 12250
box -6 -8 126 248
use OAI21X1  _13541_
timestamp 0
transform -1 0 8970 0 -1 12250
box -6 -8 106 248
use AOI22X1  _13542_
timestamp 0
transform 1 0 8290 0 1 12250
box -6 -8 126 248
use OAI21X1  _13543_
timestamp 0
transform -1 0 8410 0 -1 12730
box -6 -8 106 248
use INVX1  _13544_
timestamp 0
transform -1 0 7230 0 -1 13690
box -6 -8 66 248
use INVX1  _13545_
timestamp 0
transform 1 0 6730 0 -1 16090
box -6 -8 66 248
use INVX4  _13546_
timestamp 0
transform -1 0 7990 0 1 15130
box -6 -8 86 248
use INVX8  _13547_
timestamp 0
transform -1 0 7690 0 -1 15610
box -6 -8 126 248
use INVX1  _13548_
timestamp 0
transform 1 0 10270 0 -1 15610
box -6 -8 66 248
use NAND2X1  _13549_
timestamp 0
transform -1 0 9990 0 1 15130
box -6 -8 86 248
use OAI21X1  _13550_
timestamp 0
transform -1 0 10110 0 -1 15610
box -6 -8 106 248
use INVX1  _13551_
timestamp 0
transform 1 0 10250 0 -1 16090
box -6 -8 66 248
use NAND2X1  _13552_
timestamp 0
transform -1 0 9830 0 1 15610
box -6 -8 86 248
use OAI21X1  _13553_
timestamp 0
transform -1 0 10150 0 1 15610
box -6 -8 106 248
use MUX2X1  _13554_
timestamp 0
transform 1 0 9870 0 1 15610
box -6 -8 126 248
use INVX1  _13555_
timestamp 0
transform -1 0 7830 0 1 15610
box -6 -8 66 248
use NAND2X1  _13556_
timestamp 0
transform -1 0 8270 0 1 15610
box -6 -8 86 248
use OAI21X1  _13557_
timestamp 0
transform 1 0 7870 0 1 15610
box -6 -8 106 248
use INVX1  _13558_
timestamp 0
transform 1 0 8170 0 1 15130
box -6 -8 66 248
use NAND2X1  _13559_
timestamp 0
transform -1 0 8550 0 1 15610
box -6 -8 86 248
use OAI21X1  _13560_
timestamp 0
transform 1 0 8330 0 1 15610
box -6 -8 106 248
use MUX2X1  _13561_
timestamp 0
transform 1 0 8010 0 1 15610
box -6 -8 126 248
use MUX2X1  _13562_
timestamp 0
transform -1 0 7730 0 1 15610
box -6 -8 126 248
use NOR2X1  _13563_
timestamp 0
transform 1 0 7150 0 1 15610
box -6 -8 86 248
use NAND2X1  _13564_
timestamp 0
transform -1 0 6690 0 -1 16090
box -6 -8 86 248
use INVX1  _13565_
timestamp 0
transform 1 0 7330 0 -1 15610
box -6 -8 66 248
use NAND2X1  _13566_
timestamp 0
transform -1 0 8950 0 -1 15130
box -6 -8 86 248
use OAI21X1  _13567_
timestamp 0
transform 1 0 9410 0 1 14650
box -6 -8 106 248
use INVX2  _13568_
timestamp 0
transform 1 0 9950 0 1 14650
box -6 -8 66 248
use OAI21X1  _13569_
timestamp 0
transform 1 0 7430 0 -1 15610
box -6 -8 106 248
use OAI21X1  _13570_
timestamp 0
transform 1 0 7290 0 -1 13690
box -6 -8 106 248
use INVX4  _13571_
timestamp 0
transform -1 0 8270 0 1 12730
box -6 -8 86 248
use NAND2X1  _13572_
timestamp 0
transform -1 0 6310 0 1 12730
box -6 -8 86 248
use NOR2X1  _13573_
timestamp 0
transform 1 0 8470 0 1 14650
box -6 -8 86 248
use MUX2X1  _13574_
timestamp 0
transform -1 0 9390 0 -1 15130
box -6 -8 126 248
use MUX2X1  _13575_
timestamp 0
transform -1 0 9590 0 1 15610
box -6 -8 126 248
use MUX2X1  _13576_
timestamp 0
transform -1 0 8710 0 -1 15130
box -6 -8 126 248
use INVX1  _13577_
timestamp 0
transform -1 0 7510 0 -1 16090
box -6 -8 66 248
use NAND2X1  _13578_
timestamp 0
transform -1 0 7810 0 -1 15610
box -6 -8 86 248
use AOI21X1  _13579_
timestamp 0
transform 1 0 7850 0 -1 15610
box -6 -8 106 248
use NAND3X1  _13580_
timestamp 0
transform 1 0 8170 0 -1 15610
box -6 -8 106 248
use NAND3X1  _13581_
timestamp 0
transform -1 0 8570 0 -1 15610
box -6 -8 106 248
use NAND3X1  _13582_
timestamp 0
transform 1 0 8330 0 -1 15610
box -6 -8 106 248
use OAI22X1  _13583_
timestamp 0
transform 1 0 7990 0 -1 15610
box -6 -8 126 248
use INVX1  _13584_
timestamp 0
transform -1 0 7150 0 -1 16090
box -6 -8 66 248
use INVX8  _13585_
timestamp 0
transform 1 0 10350 0 -1 16090
box -6 -8 126 248
use INVX1  _13586_
timestamp 0
transform -1 0 9730 0 1 15130
box -6 -8 66 248
use NAND2X1  _13587_
timestamp 0
transform -1 0 9490 0 1 15130
box -6 -8 86 248
use OAI21X1  _13588_
timestamp 0
transform -1 0 9630 0 1 15130
box -6 -8 106 248
use INVX1  _13589_
timestamp 0
transform -1 0 9710 0 1 15610
box -6 -8 66 248
use NAND2X1  _13590_
timestamp 0
transform -1 0 9410 0 1 15610
box -6 -8 86 248
use OAI21X1  _13591_
timestamp 0
transform 1 0 9290 0 -1 16090
box -6 -8 106 248
use MUX2X1  _13592_
timestamp 0
transform -1 0 9090 0 -1 16090
box -6 -8 126 248
use INVX1  _13593_
timestamp 0
transform -1 0 8430 0 -1 16090
box -6 -8 66 248
use NAND2X1  _13594_
timestamp 0
transform 1 0 9350 0 1 16090
box -6 -8 86 248
use OAI21X1  _13595_
timestamp 0
transform 1 0 9190 0 1 16090
box -6 -8 106 248
use INVX1  _13596_
timestamp 0
transform 1 0 8930 0 -1 15610
box -6 -8 66 248
use NAND2X1  _13597_
timestamp 0
transform 1 0 8630 0 1 16090
box -6 -8 86 248
use OAI21X1  _13598_
timestamp 0
transform -1 0 8450 0 1 16090
box -6 -8 106 248
use MUX2X1  _13599_
timestamp 0
transform 1 0 7770 0 1 16090
box -6 -8 126 248
use MUX2X1  _13600_
timestamp 0
transform -1 0 7270 0 1 16090
box -6 -8 126 248
use NAND3X1  _13601_
timestamp 0
transform 1 0 6330 0 1 16090
box -6 -8 106 248
use MUX2X1  _13602_
timestamp 0
transform 1 0 9230 0 1 15130
box -6 -8 126 248
use MUX2X1  _13603_
timestamp 0
transform -1 0 9450 0 -1 15610
box -6 -8 126 248
use MUX2X1  _13604_
timestamp 0
transform 1 0 9070 0 1 15130
box -6 -8 126 248
use MUX2X1  _13605_
timestamp 0
transform 1 0 9170 0 1 15610
box -6 -8 126 248
use MUX2X1  _13606_
timestamp 0
transform 1 0 8850 0 1 15610
box -6 -8 126 248
use MUX2X1  _13607_
timestamp 0
transform -1 0 9130 0 1 15610
box -6 -8 126 248
use MUX2X1  _13608_
timestamp 0
transform -1 0 7570 0 1 15610
box -6 -8 126 248
use OAI21X1  _13609_
timestamp 0
transform 1 0 6830 0 -1 16570
box -6 -8 106 248
use AOI21X1  _13610_
timestamp 0
transform -1 0 6510 0 -1 16570
box -6 -8 106 248
use INVX1  _13611_
timestamp 0
transform -1 0 6230 0 1 16570
box -6 -8 66 248
use NAND3X1  _13612_
timestamp 0
transform 1 0 6550 0 -1 16570
box -6 -8 106 248
use AND2X2  _13613_
timestamp 0
transform 1 0 6270 0 -1 16570
box -6 -8 106 248
use OAI21X1  _13614_
timestamp 0
transform -1 0 6690 0 1 16090
box -6 -8 106 248
use OR2X2  _13615_
timestamp 0
transform 1 0 6330 0 -1 16090
box -6 -8 106 248
use AOI21X1  _13616_
timestamp 0
transform -1 0 6570 0 -1 16090
box -6 -8 106 248
use OAI21X1  _13617_
timestamp 0
transform -1 0 6450 0 1 12730
box -6 -8 106 248
use INVX1  _13618_
timestamp 0
transform 1 0 9150 0 -1 10810
box -6 -8 66 248
use NAND2X1  _13619_
timestamp 0
transform 1 0 9410 0 -1 10810
box -6 -8 86 248
use OAI21X1  _13620_
timestamp 0
transform 1 0 9270 0 -1 10810
box -6 -8 106 248
use NAND2X1  _13621_
timestamp 0
transform 1 0 7030 0 -1 13210
box -6 -8 86 248
use AOI21X1  _13622_
timestamp 0
transform -1 0 6210 0 -1 16570
box -6 -8 106 248
use MUX2X1  _13623_
timestamp 0
transform -1 0 9410 0 -1 14170
box -6 -8 126 248
use MUX2X1  _13624_
timestamp 0
transform 1 0 9250 0 1 14650
box -6 -8 126 248
use MUX2X1  _13625_
timestamp 0
transform -1 0 8550 0 -1 15130
box -6 -8 126 248
use NAND2X1  _13626_
timestamp 0
transform -1 0 8190 0 -1 15130
box -6 -8 86 248
use OAI22X1  _13627_
timestamp 0
transform 1 0 8250 0 -1 15130
box -6 -8 126 248
use AOI21X1  _13628_
timestamp 0
transform -1 0 8070 0 -1 15130
box -6 -8 106 248
use AOI21X1  _13629_
timestamp 0
transform -1 0 6790 0 -1 16570
box -6 -8 106 248
use NAND2X1  _13630_
timestamp 0
transform -1 0 5650 0 -1 17050
box -6 -8 86 248
use INVX1  _13631_
timestamp 0
transform -1 0 6110 0 1 16570
box -6 -8 66 248
use OAI21X1  _13632_
timestamp 0
transform -1 0 6270 0 1 16090
box -6 -8 106 248
use NAND2X1  _13633_
timestamp 0
transform -1 0 6010 0 1 16570
box -6 -8 86 248
use AOI21X1  _13634_
timestamp 0
transform -1 0 5370 0 -1 17050
box -6 -8 106 248
use NAND3X1  _13635_
timestamp 0
transform -1 0 5510 0 -1 17050
box -6 -8 106 248
use INVX1  _13636_
timestamp 0
transform -1 0 4830 0 -1 17050
box -6 -8 66 248
use OR2X2  _13637_
timestamp 0
transform -1 0 4730 0 -1 17050
box -6 -8 106 248
use NOR2X1  _13638_
timestamp 0
transform -1 0 5370 0 1 16570
box -6 -8 86 248
use INVX1  _13639_
timestamp 0
transform 1 0 5430 0 1 16570
box -6 -8 66 248
use OAI21X1  _13640_
timestamp 0
transform 1 0 4870 0 -1 17050
box -6 -8 106 248
use AOI21X1  _13641_
timestamp 0
transform 1 0 5530 0 1 16570
box -6 -8 106 248
use INVX2  _13642_
timestamp 0
transform 1 0 6790 0 1 13690
box -6 -8 66 248
use OAI21X1  _13643_
timestamp 0
transform 1 0 6590 0 1 13210
box -6 -8 106 248
use OAI21X1  _13644_
timestamp 0
transform 1 0 6750 0 1 13210
box -6 -8 106 248
use INVX1  _13645_
timestamp 0
transform 1 0 6890 0 -1 12730
box -6 -8 66 248
use INVX2  _13646_
timestamp 0
transform -1 0 6750 0 -1 13210
box -6 -8 66 248
use OAI21X1  _13647_
timestamp 0
transform -1 0 5210 0 -1 17050
box -6 -8 106 248
use INVX1  _13648_
timestamp 0
transform -1 0 5070 0 -1 17050
box -6 -8 66 248
use INVX1  _13649_
timestamp 0
transform -1 0 5890 0 1 16570
box -6 -8 66 248
use NAND3X1  _13650_
timestamp 0
transform 1 0 6830 0 1 15610
box -6 -8 106 248
use INVX1  _13651_
timestamp 0
transform 1 0 9930 0 -1 12730
box -6 -8 66 248
use NAND2X1  _13652_
timestamp 0
transform 1 0 10130 0 -1 13690
box -6 -8 86 248
use OAI21X1  _13653_
timestamp 0
transform 1 0 9990 0 -1 13690
box -6 -8 106 248
use NAND2X1  _13654_
timestamp 0
transform 1 0 9010 0 1 14650
box -6 -8 86 248
use OAI21X1  _13655_
timestamp 0
transform 1 0 8870 0 1 14650
box -6 -8 106 248
use NOR2X1  _13656_
timestamp 0
transform 1 0 7330 0 1 16090
box -6 -8 86 248
use NOR2X1  _13657_
timestamp 0
transform 1 0 6350 0 -1 17050
box -6 -8 86 248
use AOI22X1  _13658_
timestamp 0
transform -1 0 7710 0 1 16090
box -6 -8 126 248
use OAI21X1  _13659_
timestamp 0
transform 1 0 7670 0 -1 16090
box -6 -8 106 248
use NAND3X1  _13660_
timestamp 0
transform -1 0 6110 0 1 16090
box -6 -8 106 248
use INVX1  _13661_
timestamp 0
transform -1 0 5970 0 1 16090
box -6 -8 66 248
use INVX1  _13662_
timestamp 0
transform 1 0 6070 0 -1 16090
box -6 -8 66 248
use OAI21X1  _13663_
timestamp 0
transform -1 0 5850 0 1 16090
box -6 -8 106 248
use NAND3X1  _13664_
timestamp 0
transform -1 0 5750 0 -1 16570
box -6 -8 106 248
use AOI21X1  _13665_
timestamp 0
transform 1 0 5810 0 -1 16570
box -6 -8 106 248
use INVX1  _13666_
timestamp 0
transform -1 0 4450 0 -1 17050
box -6 -8 66 248
use NAND2X1  _13667_
timestamp 0
transform -1 0 4570 0 -1 17050
box -6 -8 86 248
use AOI21X1  _13668_
timestamp 0
transform 1 0 5010 0 1 16570
box -6 -8 106 248
use OAI21X1  _13669_
timestamp 0
transform 1 0 5150 0 1 16570
box -6 -8 106 248
use AOI22X1  _13670_
timestamp 0
transform -1 0 5750 0 1 12730
box -6 -8 126 248
use AOI21X1  _13671_
timestamp 0
transform 1 0 5670 0 1 16570
box -6 -8 106 248
use INVX1  _13672_
timestamp 0
transform -1 0 5690 0 1 16090
box -6 -8 66 248
use INVX1  _13673_
timestamp 0
transform 1 0 10270 0 -1 13210
box -6 -8 66 248
use NAND2X1  _13674_
timestamp 0
transform 1 0 9970 0 -1 14650
box -6 -8 86 248
use OAI21X1  _13675_
timestamp 0
transform 1 0 9830 0 -1 14650
box -6 -8 106 248
use NAND2X1  _13676_
timestamp 0
transform 1 0 9310 0 -1 14650
box -6 -8 86 248
use OAI21X1  _13677_
timestamp 0
transform 1 0 9170 0 -1 14650
box -6 -8 106 248
use NAND2X1  _13678_
timestamp 0
transform 1 0 7850 0 -1 15130
box -6 -8 86 248
use OAI21X1  _13679_
timestamp 0
transform -1 0 7810 0 -1 15130
box -6 -8 106 248
use INVX2  _13680_
timestamp 0
transform -1 0 7150 0 -1 15610
box -6 -8 66 248
use OAI21X1  _13681_
timestamp 0
transform 1 0 6290 0 1 15610
box -6 -8 106 248
use OR2X2  _13682_
timestamp 0
transform -1 0 6090 0 -1 15610
box -6 -8 106 248
use NOR2X1  _13683_
timestamp 0
transform -1 0 6650 0 -1 15610
box -6 -8 86 248
use OAI21X1  _13684_
timestamp 0
transform -1 0 6530 0 -1 15610
box -6 -8 106 248
use NAND3X1  _13685_
timestamp 0
transform -1 0 6230 0 -1 15610
box -6 -8 106 248
use NOR2X1  _13686_
timestamp 0
transform 1 0 6170 0 1 15610
box -6 -8 86 248
use AND2X2  _13687_
timestamp 0
transform -1 0 6130 0 1 15610
box -6 -8 106 248
use OAI21X1  _13688_
timestamp 0
transform -1 0 5970 0 1 15610
box -6 -8 106 248
use NAND2X1  _13689_
timestamp 0
transform 1 0 6070 0 -1 15130
box -6 -8 86 248
use AOI21X1  _13690_
timestamp 0
transform -1 0 6190 0 -1 14650
box -6 -8 106 248
use OAI21X1  _13691_
timestamp 0
transform 1 0 5950 0 -1 14650
box -6 -8 106 248
use AOI22X1  _13692_
timestamp 0
transform -1 0 6110 0 -1 13210
box -6 -8 126 248
use OAI21X1  _13693_
timestamp 0
transform -1 0 6330 0 -1 14650
box -6 -8 106 248
use INVX1  _13694_
timestamp 0
transform -1 0 7070 0 1 15130
box -6 -8 66 248
use NAND3X1  _13695_
timestamp 0
transform 1 0 6170 0 -1 16090
box -6 -8 106 248
use NAND2X1  _13696_
timestamp 0
transform 1 0 9690 0 -1 14650
box -6 -8 86 248
use INVX1  _13697_
timestamp 0
transform -1 0 9490 0 -1 14650
box -6 -8 66 248
use AOI21X1  _13698_
timestamp 0
transform -1 0 8830 0 -1 14650
box -6 -8 106 248
use NAND2X1  _13699_
timestamp 0
transform 1 0 7510 0 1 15130
box -6 -8 86 248
use OAI21X1  _13700_
timestamp 0
transform -1 0 7450 0 1 15130
box -6 -8 106 248
use NAND3X1  _13701_
timestamp 0
transform 1 0 6310 0 1 15130
box -6 -8 106 248
use NOR3X1  _13702_
timestamp 0
transform -1 0 7030 0 -1 15610
box -6 -8 186 248
use INVX1  _13703_
timestamp 0
transform 1 0 6630 0 1 15130
box -6 -8 66 248
use OAI21X1  _13704_
timestamp 0
transform -1 0 6850 0 -1 15130
box -6 -8 106 248
use NAND3X1  _13705_
timestamp 0
transform 1 0 6490 0 -1 15130
box -6 -8 106 248
use AOI21X1  _13706_
timestamp 0
transform -1 0 6570 0 1 15130
box -6 -8 106 248
use INVX1  _13707_
timestamp 0
transform -1 0 5830 0 1 15130
box -6 -8 66 248
use NAND2X1  _13708_
timestamp 0
transform 1 0 6890 0 1 14650
box -6 -8 86 248
use AND2X2  _13709_
timestamp 0
transform 1 0 6310 0 1 13210
box -6 -8 106 248
use OAI21X1  _13710_
timestamp 0
transform 1 0 6450 0 1 13210
box -6 -8 106 248
use OAI21X1  _13711_
timestamp 0
transform 1 0 6530 0 -1 13210
box -6 -8 106 248
use OAI21X1  _13712_
timestamp 0
transform -1 0 7410 0 1 11770
box -6 -8 106 248
use INVX1  _13713_
timestamp 0
transform -1 0 5870 0 1 12730
box -6 -8 66 248
use INVX1  _13714_
timestamp 0
transform 1 0 7690 0 1 14650
box -6 -8 66 248
use NAND3X1  _13715_
timestamp 0
transform 1 0 6710 0 -1 15610
box -6 -8 106 248
use AOI21X1  _13716_
timestamp 0
transform -1 0 9110 0 -1 14650
box -6 -8 106 248
use NAND2X1  _13717_
timestamp 0
transform 1 0 8350 0 1 14650
box -6 -8 86 248
use OAI21X1  _13718_
timestamp 0
transform 1 0 8210 0 1 14650
box -6 -8 106 248
use NAND3X1  _13719_
timestamp 0
transform -1 0 6770 0 -1 14650
box -6 -8 106 248
use INVX1  _13720_
timestamp 0
transform 1 0 7450 0 1 14650
box -6 -8 66 248
use OAI21X1  _13721_
timestamp 0
transform -1 0 6250 0 1 15130
box -6 -8 106 248
use NAND2X1  _13722_
timestamp 0
transform -1 0 6710 0 -1 15130
box -6 -8 86 248
use NAND3X1  _13723_
timestamp 0
transform -1 0 6490 0 -1 14650
box -6 -8 106 248
use NAND3X1  _13724_
timestamp 0
transform -1 0 7250 0 1 14650
box -6 -8 106 248
use NAND2X1  _13725_
timestamp 0
transform 1 0 7050 0 -1 15130
box -6 -8 86 248
use NAND3X1  _13726_
timestamp 0
transform -1 0 7110 0 1 14650
box -6 -8 106 248
use NAND2X1  _13727_
timestamp 0
transform -1 0 6310 0 1 13690
box -6 -8 86 248
use AOI21X1  _13728_
timestamp 0
transform 1 0 6270 0 -1 15610
box -6 -8 106 248
use NOR2X1  _13729_
timestamp 0
transform -1 0 5950 0 1 15130
box -6 -8 86 248
use OAI21X1  _13730_
timestamp 0
transform 1 0 6610 0 1 14650
box -6 -8 106 248
use NAND2X1  _13731_
timestamp 0
transform -1 0 6830 0 1 14650
box -6 -8 86 248
use AOI21X1  _13732_
timestamp 0
transform -1 0 6170 0 1 13690
box -6 -8 106 248
use OAI21X1  _13733_
timestamp 0
transform -1 0 6170 0 -1 13690
box -6 -8 106 248
use AOI22X1  _13734_
timestamp 0
transform 1 0 5930 0 1 12730
box -6 -8 126 248
use INVX1  _13735_
timestamp 0
transform -1 0 6910 0 1 12250
box -6 -8 66 248
use AOI21X1  _13736_
timestamp 0
transform -1 0 6630 0 -1 14650
box -6 -8 106 248
use AND2X2  _13737_
timestamp 0
transform 1 0 6210 0 -1 15130
box -6 -8 106 248
use NAND3X1  _13738_
timestamp 0
transform 1 0 6350 0 -1 15130
box -6 -8 106 248
use AOI21X1  _13739_
timestamp 0
transform -1 0 6110 0 1 15130
box -6 -8 106 248
use OAI21X1  _13740_
timestamp 0
transform 1 0 6450 0 1 14650
box -6 -8 106 248
use AOI21X1  _13741_
timestamp 0
transform 1 0 6470 0 -1 14170
box -6 -8 106 248
use INVX1  _13742_
timestamp 0
transform -1 0 7430 0 -1 14650
box -6 -8 66 248
use NAND3X1  _13743_
timestamp 0
transform 1 0 6890 0 -1 15130
box -6 -8 106 248
use INVX1  _13744_
timestamp 0
transform -1 0 9770 0 1 14170
box -6 -8 66 248
use NOR2X1  _13745_
timestamp 0
transform 1 0 9670 0 1 14650
box -6 -8 86 248
use INVX1  _13746_
timestamp 0
transform -1 0 9630 0 1 14650
box -6 -8 66 248
use OAI21X1  _13747_
timestamp 0
transform 1 0 8730 0 1 14650
box -6 -8 106 248
use NAND3X1  _13748_
timestamp 0
transform 1 0 7290 0 1 14650
box -6 -8 106 248
use INVX1  _13749_
timestamp 0
transform -1 0 7170 0 -1 14650
box -6 -8 66 248
use OAI21X1  _13750_
timestamp 0
transform 1 0 6810 0 -1 14650
box -6 -8 106 248
use NAND2X1  _13751_
timestamp 0
transform -1 0 7050 0 -1 14650
box -6 -8 86 248
use NAND3X1  _13752_
timestamp 0
transform -1 0 7310 0 -1 14650
box -6 -8 106 248
use NAND3X1  _13753_
timestamp 0
transform 1 0 7190 0 1 14170
box -6 -8 106 248
use NAND2X1  _13754_
timestamp 0
transform -1 0 7010 0 1 14170
box -6 -8 86 248
use NAND3X1  _13755_
timestamp 0
transform -1 0 7150 0 1 14170
box -6 -8 106 248
use NAND2X1  _13756_
timestamp 0
transform -1 0 6850 0 -1 14170
box -6 -8 86 248
use INVX1  _13757_
timestamp 0
transform 1 0 7050 0 -1 13690
box -6 -8 66 248
use NOR2X1  _13758_
timestamp 0
transform -1 0 7010 0 -1 13690
box -6 -8 86 248
use OAI21X1  _13759_
timestamp 0
transform 1 0 6470 0 -1 13690
box -6 -8 106 248
use OAI21X1  _13760_
timestamp 0
transform 1 0 6610 0 -1 13690
box -6 -8 106 248
use OAI21X1  _13761_
timestamp 0
transform -1 0 7010 0 -1 14170
box -6 -8 106 248
use INVX1  _13762_
timestamp 0
transform -1 0 6950 0 1 13690
box -6 -8 66 248
use OAI21X1  _13763_
timestamp 0
transform 1 0 6770 0 -1 13690
box -6 -8 106 248
use OAI21X1  _13764_
timestamp 0
transform -1 0 6810 0 1 12250
box -6 -8 106 248
use INVX1  _13765_
timestamp 0
transform -1 0 7030 0 1 12250
box -6 -8 66 248
use OAI21X1  _13766_
timestamp 0
transform 1 0 6630 0 1 13690
box -6 -8 106 248
use NOR2X1  _13767_
timestamp 0
transform 1 0 6350 0 1 13690
box -6 -8 86 248
use AOI21X1  _13768_
timestamp 0
transform 1 0 6490 0 1 13690
box -6 -8 106 248
use INVX1  _13769_
timestamp 0
transform -1 0 8170 0 -1 14170
box -6 -8 66 248
use OR2X2  _13770_
timestamp 0
transform 1 0 7930 0 -1 14650
box -6 -8 106 248
use OAI21X1  _13771_
timestamp 0
transform 1 0 8590 0 1 14650
box -6 -8 106 248
use NAND3X1  _13772_
timestamp 0
transform -1 0 8470 0 -1 14170
box -6 -8 106 248
use NOR2X1  _13773_
timestamp 0
transform -1 0 8170 0 -1 14650
box -6 -8 86 248
use INVX1  _13774_
timestamp 0
transform 1 0 8350 0 1 14170
box -6 -8 66 248
use OAI21X1  _13775_
timestamp 0
transform -1 0 8170 0 1 14170
box -6 -8 106 248
use NAND3X1  _13776_
timestamp 0
transform -1 0 8070 0 -1 14170
box -6 -8 106 248
use NAND3X1  _13777_
timestamp 0
transform -1 0 8330 0 -1 14170
box -6 -8 106 248
use OAI21X1  _13778_
timestamp 0
transform 1 0 8210 0 1 14170
box -6 -8 106 248
use NAND3X1  _13779_
timestamp 0
transform -1 0 7890 0 1 13690
box -6 -8 106 248
use AND2X2  _13780_
timestamp 0
transform 1 0 7550 0 1 13690
box -6 -8 106 248
use INVX1  _13781_
timestamp 0
transform -1 0 7350 0 1 13690
box -6 -8 66 248
use AOI21X1  _13782_
timestamp 0
transform -1 0 7250 0 1 13690
box -6 -8 106 248
use OAI21X1  _13783_
timestamp 0
transform -1 0 7090 0 1 13690
box -6 -8 106 248
use AOI22X1  _13784_
timestamp 0
transform -1 0 7030 0 1 13210
box -6 -8 126 248
use NAND2X1  _13785_
timestamp 0
transform 1 0 6790 0 1 14170
box -6 -8 86 248
use AND2X2  _13786_
timestamp 0
transform -1 0 6750 0 1 14170
box -6 -8 106 248
use AND2X2  _13787_
timestamp 0
transform 1 0 6330 0 -1 14170
box -6 -8 106 248
use NAND3X1  _13788_
timestamp 0
transform -1 0 6710 0 -1 14170
box -6 -8 106 248
use OAI21X1  _13789_
timestamp 0
transform 1 0 6510 0 1 14170
box -6 -8 106 248
use INVX1  _13790_
timestamp 0
transform -1 0 7750 0 1 13690
box -6 -8 66 248
use AOI21X1  _13791_
timestamp 0
transform -1 0 7490 0 1 13690
box -6 -8 106 248
use INVX1  _13792_
timestamp 0
transform -1 0 9050 0 -1 13690
box -6 -8 66 248
use NOR3X1  _13793_
timestamp 0
transform 1 0 8210 0 -1 14650
box -6 -8 186 248
use INVX1  _13794_
timestamp 0
transform -1 0 8630 0 1 13690
box -6 -8 66 248
use OAI21X1  _13795_
timestamp 0
transform 1 0 8590 0 -1 14650
box -6 -8 106 248
use NAND3X1  _13796_
timestamp 0
transform -1 0 8510 0 1 13690
box -6 -8 106 248
use INVX1  _13797_
timestamp 0
transform 1 0 8650 0 -1 14170
box -6 -8 66 248
use OAI21X1  _13798_
timestamp 0
transform 1 0 8510 0 -1 14170
box -6 -8 106 248
use NAND3X1  _13799_
timestamp 0
transform -1 0 8210 0 1 13690
box -6 -8 106 248
use NAND3X1  _13800_
timestamp 0
transform 1 0 8670 0 1 13690
box -6 -8 106 248
use OAI21X1  _13801_
timestamp 0
transform -1 0 8870 0 -1 14170
box -6 -8 106 248
use NAND3X1  _13802_
timestamp 0
transform -1 0 8930 0 -1 13690
box -6 -8 106 248
use AND2X2  _13803_
timestamp 0
transform -1 0 7910 0 -1 13690
box -6 -8 106 248
use AND2X2  _13804_
timestamp 0
transform -1 0 7430 0 1 13210
box -6 -8 106 248
use OAI21X1  _13805_
timestamp 0
transform 1 0 7470 0 1 13210
box -6 -8 106 248
use OAI21X1  _13806_
timestamp 0
transform -1 0 7430 0 -1 13210
box -6 -8 106 248
use OAI21X1  _13807_
timestamp 0
transform -1 0 7530 0 -1 11770
box -6 -8 106 248
use INVX1  _13808_
timestamp 0
transform -1 0 9890 0 1 13690
box -6 -8 66 248
use OAI21X1  _13809_
timestamp 0
transform -1 0 8970 0 -1 14650
box -6 -8 106 248
use INVX1  _13810_
timestamp 0
transform 1 0 9030 0 -1 14170
box -6 -8 66 248
use AOI21X1  _13811_
timestamp 0
transform 1 0 9150 0 -1 14170
box -6 -8 106 248
use NAND3X1  _13812_
timestamp 0
transform 1 0 9090 0 1 13690
box -6 -8 106 248
use NAND2X1  _13813_
timestamp 0
transform 1 0 9250 0 1 13690
box -6 -8 86 248
use NAND2X1  _13814_
timestamp 0
transform -1 0 8990 0 -1 14170
box -6 -8 86 248
use OAI21X1  _13815_
timestamp 0
transform -1 0 9050 0 1 13690
box -6 -8 106 248
use NAND2X1  _13816_
timestamp 0
transform -1 0 8890 0 1 13690
box -6 -8 86 248
use INVX1  _13817_
timestamp 0
transform 1 0 9250 0 -1 13690
box -6 -8 66 248
use AND2X2  _13818_
timestamp 0
transform 1 0 9390 0 1 13690
box -6 -8 106 248
use NAND2X1  _13819_
timestamp 0
transform -1 0 9430 0 -1 13690
box -6 -8 86 248
use NAND3X1  _13820_
timestamp 0
transform 1 0 9110 0 -1 13690
box -6 -8 106 248
use NAND2X1  _13821_
timestamp 0
transform 1 0 8550 0 -1 13690
box -6 -8 86 248
use AOI21X1  _13822_
timestamp 0
transform -1 0 8350 0 1 13690
box -6 -8 106 248
use AOI21X1  _13823_
timestamp 0
transform 1 0 7950 0 1 13690
box -6 -8 106 248
use NAND3X1  _13824_
timestamp 0
transform 1 0 7670 0 -1 13690
box -6 -8 106 248
use AOI21X1  _13825_
timestamp 0
transform 1 0 8270 0 -1 13690
box -6 -8 106 248
use AND2X2  _13826_
timestamp 0
transform -1 0 8510 0 -1 13690
box -6 -8 106 248
use NAND3X1  _13827_
timestamp 0
transform 1 0 7970 0 -1 13690
box -6 -8 106 248
use OAI21X1  _13828_
timestamp 0
transform 1 0 8110 0 -1 13690
box -6 -8 106 248
use OAI21X1  _13829_
timestamp 0
transform -1 0 8150 0 1 13210
box -6 -8 106 248
use OR2X2  _13830_
timestamp 0
transform -1 0 7750 0 -1 13210
box -6 -8 106 248
use AOI22X1  _13831_
timestamp 0
transform 1 0 7110 0 1 12730
box -6 -8 126 248
use NAND2X1  _13832_
timestamp 0
transform -1 0 7450 0 1 12250
box -6 -8 86 248
use INVX1  _13833_
timestamp 0
transform -1 0 8410 0 1 13210
box -6 -8 66 248
use NAND2X1  _13834_
timestamp 0
transform -1 0 10190 0 -1 14170
box -6 -8 86 248
use INVX1  _13835_
timestamp 0
transform 1 0 10470 0 1 14170
box -6 -8 66 248
use NAND2X1  _13836_
timestamp 0
transform 1 0 10050 0 1 14170
box -6 -8 86 248
use NAND2X1  _13837_
timestamp 0
transform -1 0 10070 0 -1 14170
box -6 -8 86 248
use INVX1  _13838_
timestamp 0
transform 1 0 9790 0 -1 13210
box -6 -8 66 248
use NAND2X1  _13839_
timestamp 0
transform -1 0 9570 0 1 13210
box -6 -8 86 248
use NAND2X1  _13840_
timestamp 0
transform -1 0 9550 0 -1 13690
box -6 -8 86 248
use NAND2X1  _13841_
timestamp 0
transform 1 0 9350 0 1 13210
box -6 -8 86 248
use INVX1  _13842_
timestamp 0
transform -1 0 8090 0 -1 13210
box -6 -8 66 248
use NOR3X1  _13843_
timestamp 0
transform -1 0 7970 0 -1 13210
box -6 -8 186 248
use AOI21X1  _13844_
timestamp 0
transform 1 0 8210 0 1 13210
box -6 -8 106 248
use OAI21X1  _13845_
timestamp 0
transform -1 0 8010 0 1 13210
box -6 -8 106 248
use OAI21X1  _13846_
timestamp 0
transform -1 0 7590 0 -1 13210
box -6 -8 106 248
use NAND2X1  _13847_
timestamp 0
transform 1 0 7490 0 1 12250
box -6 -8 86 248
use NAND2X1  _13848_
timestamp 0
transform -1 0 8530 0 1 13210
box -6 -8 86 248
use INVX1  _13849_
timestamp 0
transform -1 0 5890 0 -1 17050
box -6 -8 66 248
use NAND2X1  _13850_
timestamp 0
transform -1 0 5770 0 -1 17050
box -6 -8 86 248
use OAI21X1  _13851_
timestamp 0
transform -1 0 6050 0 -1 17050
box -6 -8 106 248
use NAND2X1  _13852_
timestamp 0
transform -1 0 6170 0 -1 17050
box -6 -8 86 248
use NOR2X1  _13853_
timestamp 0
transform -1 0 6810 0 1 16090
box -6 -8 86 248
use NOR2X1  _13854_
timestamp 0
transform 1 0 7030 0 1 16090
box -6 -8 86 248
use AOI22X1  _13855_
timestamp 0
transform 1 0 6850 0 1 16090
box -6 -8 126 248
use NAND3X1  _13856_
timestamp 0
transform -1 0 6850 0 1 16570
box -6 -8 106 248
use NAND2X1  _13857_
timestamp 0
transform -1 0 7870 0 1 14650
box -6 -8 86 248
use OAI21X1  _13858_
timestamp 0
transform -1 0 8030 0 1 14650
box -6 -8 106 248
use NAND2X1  _13859_
timestamp 0
transform 1 0 6730 0 1 15130
box -6 -8 86 248
use OAI21X1  _13860_
timestamp 0
transform 1 0 6690 0 1 15610
box -6 -8 106 248
use MUX2X1  _13861_
timestamp 0
transform -1 0 8070 0 -1 16090
box -6 -8 126 248
use NAND2X1  _13862_
timestamp 0
transform 1 0 7990 0 1 16570
box -6 -8 86 248
use AND2X2  _13863_
timestamp 0
transform 1 0 7850 0 1 16570
box -6 -8 106 248
use NOR2X1  _13864_
timestamp 0
transform -1 0 8110 0 1 15130
box -6 -8 86 248
use NAND2X1  _13865_
timestamp 0
transform -1 0 7510 0 1 16570
box -6 -8 86 248
use NAND2X1  _13866_
timestamp 0
transform 1 0 7950 0 -1 16570
box -6 -8 86 248
use NAND2X1  _13867_
timestamp 0
transform 1 0 7550 0 1 16570
box -6 -8 86 248
use OAI21X1  _13868_
timestamp 0
transform 1 0 7690 0 1 16570
box -6 -8 106 248
use OAI21X1  _13869_
timestamp 0
transform 1 0 8610 0 -1 15610
box -6 -8 106 248
use OAI21X1  _13870_
timestamp 0
transform 1 0 8690 0 -1 13690
box -6 -8 106 248
use NAND2X1  _13871_
timestamp 0
transform -1 0 8250 0 1 12250
box -6 -8 86 248
use NOR2X1  _13872_
timestamp 0
transform -1 0 8330 0 -1 16090
box -6 -8 86 248
use NAND2X1  _13873_
timestamp 0
transform 1 0 5530 0 -1 16570
box -6 -8 86 248
use OAI21X1  _13874_
timestamp 0
transform -1 0 6050 0 -1 16570
box -6 -8 106 248
use NAND2X1  _13875_
timestamp 0
transform -1 0 6370 0 1 16570
box -6 -8 86 248
use OAI21X1  _13876_
timestamp 0
transform -1 0 6510 0 1 16570
box -6 -8 106 248
use MUX2X1  _13877_
timestamp 0
transform -1 0 6690 0 1 16570
box -6 -8 126 248
use NAND2X1  _13878_
timestamp 0
transform -1 0 7250 0 1 16570
box -6 -8 86 248
use NAND2X1  _13879_
timestamp 0
transform 1 0 7790 0 -1 14650
box -6 -8 86 248
use OAI21X1  _13880_
timestamp 0
transform 1 0 7650 0 -1 14650
box -6 -8 106 248
use INVX1  _13881_
timestamp 0
transform -1 0 7170 0 -1 16570
box -6 -8 66 248
use NAND2X1  _13882_
timestamp 0
transform 1 0 7570 0 1 14650
box -6 -8 86 248
use OAI21X1  _13883_
timestamp 0
transform 1 0 7310 0 -1 15130
box -6 -8 106 248
use NAND2X1  _13884_
timestamp 0
transform -1 0 6970 0 1 16570
box -6 -8 86 248
use OAI21X1  _13885_
timestamp 0
transform -1 0 7130 0 1 16570
box -6 -8 106 248
use OAI21X1  _13886_
timestamp 0
transform -1 0 7390 0 1 16570
box -6 -8 106 248
use NAND3X1  _13887_
timestamp 0
transform -1 0 8230 0 1 16570
box -6 -8 106 248
use MUX2X1  _13888_
timestamp 0
transform -1 0 7510 0 -1 16570
box -6 -8 126 248
use MUX2X1  _13889_
timestamp 0
transform 1 0 7230 0 -1 16570
box -6 -8 126 248
use OAI21X1  _13890_
timestamp 0
transform -1 0 8310 0 -1 16570
box -6 -8 106 248
use AOI21X1  _13891_
timestamp 0
transform 1 0 8490 0 -1 16570
box -6 -8 106 248
use INVX1  _13892_
timestamp 0
transform 1 0 8810 0 -1 16570
box -6 -8 66 248
use NAND3X1  _13893_
timestamp 0
transform 1 0 8350 0 -1 16570
box -6 -8 106 248
use AND2X2  _13894_
timestamp 0
transform -1 0 8750 0 -1 16570
box -6 -8 106 248
use NAND2X1  _13895_
timestamp 0
transform 1 0 8230 0 1 16090
box -6 -8 86 248
use OR2X2  _13896_
timestamp 0
transform -1 0 8190 0 1 16090
box -6 -8 106 248
use AOI21X1  _13897_
timestamp 0
transform -1 0 8030 0 1 16090
box -6 -8 106 248
use OAI21X1  _13898_
timestamp 0
transform 1 0 8030 0 1 12250
box -6 -8 106 248
use NAND2X1  _13899_
timestamp 0
transform -1 0 7610 0 1 12730
box -6 -8 86 248
use AOI21X1  _13900_
timestamp 0
transform 1 0 8490 0 1 16090
box -6 -8 106 248
use NAND2X1  _13901_
timestamp 0
transform 1 0 8450 0 1 16570
box -6 -8 86 248
use NAND2X1  _13902_
timestamp 0
transform 1 0 9570 0 1 14170
box -6 -8 86 248
use OAI21X1  _13903_
timestamp 0
transform 1 0 9530 0 -1 14650
box -6 -8 106 248
use NAND2X1  _13904_
timestamp 0
transform -1 0 8890 0 1 15130
box -6 -8 86 248
use OAI21X1  _13905_
timestamp 0
transform -1 0 9230 0 -1 15130
box -6 -8 106 248
use NAND2X1  _13906_
timestamp 0
transform -1 0 6310 0 -1 17050
box -6 -8 86 248
use NAND2X1  _13907_
timestamp 0
transform -1 0 6690 0 -1 17050
box -6 -8 86 248
use NAND2X1  _13908_
timestamp 0
transform 1 0 6490 0 -1 17050
box -6 -8 86 248
use AOI21X1  _13909_
timestamp 0
transform -1 0 7350 0 -1 17050
box -6 -8 106 248
use INVX1  _13910_
timestamp 0
transform 1 0 8570 0 1 16570
box -6 -8 66 248
use NAND3X1  _13911_
timestamp 0
transform 1 0 8690 0 1 16570
box -6 -8 106 248
use AOI21X1  _13912_
timestamp 0
transform 1 0 8070 0 -1 16570
box -6 -8 106 248
use OAI21X1  _13913_
timestamp 0
transform 1 0 8930 0 -1 16570
box -6 -8 106 248
use NAND3X1  _13914_
timestamp 0
transform 1 0 9050 0 1 16090
box -6 -8 106 248
use INVX1  _13915_
timestamp 0
transform 1 0 8870 0 -1 16090
box -6 -8 66 248
use AOI21X1  _13916_
timestamp 0
transform -1 0 9010 0 1 16090
box -6 -8 106 248
use NOR2X1  _13917_
timestamp 0
transform 1 0 8750 0 -1 16090
box -6 -8 86 248
use AND2X2  _13918_
timestamp 0
transform -1 0 8590 0 -1 16090
box -6 -8 106 248
use NOR2X1  _13919_
timestamp 0
transform -1 0 8710 0 -1 16090
box -6 -8 86 248
use OAI21X1  _13920_
timestamp 0
transform 1 0 8770 0 -1 15610
box -6 -8 106 248
use OAI21X1  _13921_
timestamp 0
transform -1 0 7750 0 1 12730
box -6 -8 106 248
use OAI21X1  _13922_
timestamp 0
transform 1 0 8750 0 1 16090
box -6 -8 106 248
use INVX1  _13923_
timestamp 0
transform -1 0 7210 0 -1 17050
box -6 -8 66 248
use NAND2X1  _13924_
timestamp 0
transform -1 0 9610 0 1 13690
box -6 -8 86 248
use OAI21X1  _13925_
timestamp 0
transform -1 0 9770 0 1 13690
box -6 -8 106 248
use MUX2X1  _13926_
timestamp 0
transform 1 0 10050 0 1 14650
box -6 -8 126 248
use NOR2X1  _13927_
timestamp 0
transform 1 0 9450 0 -1 16090
box -6 -8 86 248
use NAND2X1  _13928_
timestamp 0
transform 1 0 7670 0 -1 16570
box -6 -8 86 248
use NAND2X1  _13929_
timestamp 0
transform 1 0 7550 0 -1 16570
box -6 -8 86 248
use NAND2X1  _13930_
timestamp 0
transform 1 0 7810 0 -1 16570
box -6 -8 86 248
use OR2X2  _13931_
timestamp 0
transform 1 0 9490 0 -1 16570
box -6 -8 106 248
use OAI21X1  _13932_
timestamp 0
transform 1 0 8850 0 1 16570
box -6 -8 106 248
use OR2X2  _13933_
timestamp 0
transform -1 0 9090 0 1 16570
box -6 -8 106 248
use OAI21X1  _13934_
timestamp 0
transform -1 0 9170 0 -1 16570
box -6 -8 106 248
use AOI21X1  _13935_
timestamp 0
transform -1 0 8030 0 -1 17050
box -6 -8 106 248
use INVX1  _13936_
timestamp 0
transform -1 0 7570 0 -1 17050
box -6 -8 66 248
use NAND3X1  _13937_
timestamp 0
transform -1 0 7870 0 -1 17050
box -6 -8 106 248
use NAND2X1  _13938_
timestamp 0
transform -1 0 7470 0 -1 17050
box -6 -8 86 248
use OR2X2  _13939_
timestamp 0
transform -1 0 6850 0 -1 17050
box -6 -8 106 248
use NAND2X1  _13940_
timestamp 0
transform -1 0 7090 0 -1 17050
box -6 -8 86 248
use NAND2X1  _13941_
timestamp 0
transform -1 0 6970 0 -1 17050
box -6 -8 86 248
use AOI22X1  _13942_
timestamp 0
transform -1 0 8270 0 -1 12730
box -6 -8 126 248
use AOI21X1  _13943_
timestamp 0
transform 1 0 7610 0 -1 17050
box -6 -8 106 248
use NAND2X1  _13944_
timestamp 0
transform 1 0 10330 0 1 14170
box -6 -8 86 248
use OAI21X1  _13945_
timestamp 0
transform 1 0 10170 0 1 14170
box -6 -8 106 248
use NAND2X1  _13946_
timestamp 0
transform -1 0 10410 0 1 14650
box -6 -8 86 248
use OAI21X1  _13947_
timestamp 0
transform 1 0 10470 0 1 14650
box -6 -8 106 248
use NAND2X1  _13948_
timestamp 0
transform 1 0 10610 0 1 14650
box -6 -8 86 248
use OAI21X1  _13949_
timestamp 0
transform 1 0 10530 0 -1 16090
box -6 -8 106 248
use INVX1  _13950_
timestamp 0
transform 1 0 10230 0 1 16570
box -6 -8 66 248
use NAND3X1  _13951_
timestamp 0
transform 1 0 8290 0 1 16570
box -6 -8 106 248
use OAI21X1  _13952_
timestamp 0
transform 1 0 9530 0 1 16570
box -6 -8 106 248
use OR2X2  _13953_
timestamp 0
transform 1 0 9990 0 1 16090
box -6 -8 106 248
use NOR2X1  _13954_
timestamp 0
transform 1 0 9410 0 1 16570
box -6 -8 86 248
use OAI21X1  _13955_
timestamp 0
transform -1 0 10390 0 1 16090
box -6 -8 106 248
use NAND3X1  _13956_
timestamp 0
transform -1 0 10250 0 1 16090
box -6 -8 106 248
use OR2X2  _13957_
timestamp 0
transform 1 0 10750 0 -1 16570
box -6 -8 106 248
use OAI21X1  _13958_
timestamp 0
transform 1 0 10450 0 1 16090
box -6 -8 106 248
use NAND3X1  _13959_
timestamp 0
transform 1 0 10610 0 -1 16570
box -6 -8 106 248
use NAND2X1  _13960_
timestamp 0
transform 1 0 9790 0 -1 16570
box -6 -8 86 248
use OR2X2  _13961_
timestamp 0
transform -1 0 8190 0 -1 17050
box -6 -8 106 248
use NAND2X1  _13962_
timestamp 0
transform 1 0 9270 0 1 16570
box -6 -8 86 248
use NAND2X1  _13963_
timestamp 0
transform -1 0 9230 0 1 16570
box -6 -8 86 248
use AOI22X1  _13964_
timestamp 0
transform -1 0 9490 0 1 12250
box -6 -8 126 248
use INVX1  _13965_
timestamp 0
transform 1 0 9110 0 1 12250
box -6 -8 66 248
use OAI21X1  _13966_
timestamp 0
transform 1 0 9650 0 -1 16570
box -6 -8 106 248
use NAND2X1  _13967_
timestamp 0
transform -1 0 9270 0 -1 17050
box -6 -8 86 248
use NOR2X1  _13968_
timestamp 0
transform 1 0 10250 0 -1 14650
box -6 -8 86 248
use AOI21X1  _13969_
timestamp 0
transform 1 0 10090 0 -1 14650
box -6 -8 106 248
use NAND2X1  _13970_
timestamp 0
transform -1 0 9230 0 -1 16090
box -6 -8 86 248
use OAI21X1  _13971_
timestamp 0
transform 1 0 9850 0 -1 16090
box -6 -8 106 248
use INVX1  _13972_
timestamp 0
transform -1 0 8890 0 -1 17050
box -6 -8 66 248
use NAND3X1  _13973_
timestamp 0
transform -1 0 8670 0 -1 17050
box -6 -8 106 248
use NOR2X1  _13974_
timestamp 0
transform 1 0 9370 0 -1 16570
box -6 -8 86 248
use NAND3X1  _13975_
timestamp 0
transform 1 0 9230 0 -1 16570
box -6 -8 106 248
use OAI21X1  _13976_
timestamp 0
transform -1 0 9770 0 1 16570
box -6 -8 106 248
use NAND2X1  _13977_
timestamp 0
transform -1 0 8790 0 -1 17050
box -6 -8 86 248
use AOI21X1  _13978_
timestamp 0
transform -1 0 8350 0 -1 17050
box -6 -8 106 248
use INVX1  _13979_
timestamp 0
transform -1 0 9970 0 -1 16570
box -6 -8 66 248
use NAND3X1  _13980_
timestamp 0
transform 1 0 8410 0 -1 17050
box -6 -8 106 248
use NAND2X1  _13981_
timestamp 0
transform 1 0 9870 0 1 16090
box -6 -8 86 248
use NOR2X1  _13982_
timestamp 0
transform -1 0 9710 0 1 16090
box -6 -8 86 248
use AND2X2  _13983_
timestamp 0
transform 1 0 9710 0 -1 16090
box -6 -8 106 248
use OAI21X1  _13984_
timestamp 0
transform -1 0 9670 0 -1 16090
box -6 -8 106 248
use OAI21X1  _13985_
timestamp 0
transform 1 0 9230 0 1 12250
box -6 -8 106 248
use INVX1  _13986_
timestamp 0
transform 1 0 9530 0 -1 12730
box -6 -8 66 248
use NAND3X1  _13987_
timestamp 0
transform 1 0 10350 0 1 16570
box -6 -8 106 248
use AOI21X1  _13988_
timestamp 0
transform 1 0 10370 0 -1 14650
box -6 -8 106 248
use NAND2X1  _13989_
timestamp 0
transform 1 0 10530 0 -1 14650
box -6 -8 86 248
use OAI21X1  _13990_
timestamp 0
transform 1 0 10390 0 -1 15130
box -6 -8 106 248
use NAND3X1  _13991_
timestamp 0
transform -1 0 10870 0 -1 15610
box -6 -8 106 248
use NOR3X1  _13992_
timestamp 0
transform 1 0 10010 0 -1 16090
box -6 -8 186 248
use INVX1  _13993_
timestamp 0
transform 1 0 10910 0 -1 15610
box -6 -8 66 248
use OAI21X1  _13994_
timestamp 0
transform 1 0 10710 0 1 15610
box -6 -8 106 248
use NAND2X1  _13995_
timestamp 0
transform 1 0 10650 0 -1 15610
box -6 -8 86 248
use NAND2X1  _13996_
timestamp 0
transform 1 0 10370 0 -1 15610
box -6 -8 86 248
use NAND3X1  _13997_
timestamp 0
transform -1 0 10610 0 -1 15610
box -6 -8 106 248
use NAND2X1  _13998_
timestamp 0
transform -1 0 10230 0 1 15130
box -6 -8 86 248
use AOI21X1  _13999_
timestamp 0
transform -1 0 10570 0 -1 16570
box -6 -8 106 248
use NOR2X1  _14000_
timestamp 0
transform -1 0 10050 0 1 16570
box -6 -8 86 248
use OAI21X1  _14001_
timestamp 0
transform 1 0 9830 0 1 16570
box -6 -8 106 248
use NAND2X1  _14002_
timestamp 0
transform -1 0 9830 0 1 16090
box -6 -8 86 248
use NOR2X1  _14003_
timestamp 0
transform -1 0 9850 0 1 15130
box -6 -8 86 248
use AND2X2  _14004_
timestamp 0
transform -1 0 10390 0 1 15130
box -6 -8 106 248
use AND2X2  _14005_
timestamp 0
transform -1 0 10410 0 -1 16570
box -6 -8 106 248
use NAND3X1  _14006_
timestamp 0
transform -1 0 10270 0 -1 16570
box -6 -8 106 248
use AOI21X1  _14007_
timestamp 0
transform -1 0 10190 0 1 16570
box -6 -8 106 248
use OAI21X1  _14008_
timestamp 0
transform 1 0 10010 0 -1 16570
box -6 -8 106 248
use NOR2X1  _14009_
timestamp 0
transform -1 0 10050 0 -1 15130
box -6 -8 86 248
use OAI21X1  _14010_
timestamp 0
transform -1 0 9690 0 -1 15130
box -6 -8 106 248
use NAND2X1  _14011_
timestamp 0
transform -1 0 9750 0 -1 13210
box -6 -8 86 248
use OAI21X1  _14012_
timestamp 0
transform 1 0 9630 0 -1 12730
box -6 -8 106 248
use INVX1  _14013_
timestamp 0
transform -1 0 8750 0 1 12730
box -6 -8 66 248
use INVX1  _14014_
timestamp 0
transform -1 0 9910 0 -1 15130
box -6 -8 66 248
use NAND2X1  _14015_
timestamp 0
transform -1 0 10610 0 -1 15130
box -6 -8 86 248
use NOR2X1  _14016_
timestamp 0
transform 1 0 10750 0 1 14650
box -6 -8 86 248
use INVX1  _14017_
timestamp 0
transform -1 0 10710 0 -1 14650
box -6 -8 66 248
use OAI21X1  _14018_
timestamp 0
transform 1 0 10890 0 1 14650
box -6 -8 106 248
use NAND3X1  _14019_
timestamp 0
transform -1 0 10810 0 1 15130
box -6 -8 106 248
use INVX1  _14020_
timestamp 0
transform -1 0 10890 0 -1 15130
box -6 -8 66 248
use OAI21X1  _14021_
timestamp 0
transform 1 0 11010 0 -1 15610
box -6 -8 106 248
use NAND2X1  _14022_
timestamp 0
transform 1 0 11130 0 1 15130
box -6 -8 86 248
use NAND3X1  _14023_
timestamp 0
transform -1 0 10670 0 1 15130
box -6 -8 106 248
use NAND3X1  _14024_
timestamp 0
transform -1 0 11090 0 1 15130
box -6 -8 106 248
use NAND2X1  _14025_
timestamp 0
transform 1 0 11270 0 1 15130
box -6 -8 86 248
use NAND3X1  _14026_
timestamp 0
transform -1 0 10950 0 1 15130
box -6 -8 106 248
use NAND2X1  _14027_
timestamp 0
transform 1 0 10430 0 1 15130
box -6 -8 86 248
use OAI21X1  _14028_
timestamp 0
transform -1 0 9550 0 -1 15130
box -6 -8 106 248
use NOR2X1  _14029_
timestamp 0
transform -1 0 9810 0 -1 15130
box -6 -8 86 248
use INVX1  _14030_
timestamp 0
transform 1 0 10230 0 1 14650
box -6 -8 66 248
use AOI21X1  _14031_
timestamp 0
transform -1 0 9890 0 1 14650
box -6 -8 106 248
use AOI22X1  _14032_
timestamp 0
transform 1 0 8950 0 1 12730
box -6 -8 126 248
use OAI21X1  _14033_
timestamp 0
transform 1 0 10250 0 -1 15130
box -6 -8 106 248
use NOR2X1  _14034_
timestamp 0
transform -1 0 10110 0 1 15130
box -6 -8 86 248
use AOI21X1  _14035_
timestamp 0
transform 1 0 10110 0 -1 15130
box -6 -8 106 248
use INVX1  _14036_
timestamp 0
transform 1 0 10510 0 -1 13210
box -6 -8 66 248
use NAND3X1  _14037_
timestamp 0
transform -1 0 10770 0 -1 15130
box -6 -8 106 248
use INVX1  _14038_
timestamp 0
transform -1 0 10670 0 -1 14170
box -6 -8 66 248
use OAI21X1  _14039_
timestamp 0
transform 1 0 10650 0 1 13690
box -6 -8 106 248
use INVX1  _14040_
timestamp 0
transform -1 0 10910 0 -1 13690
box -6 -8 66 248
use NAND3X1  _14041_
timestamp 0
transform 1 0 10870 0 1 13210
box -6 -8 106 248
use OAI21X1  _14042_
timestamp 0
transform 1 0 11050 0 1 14650
box -6 -8 106 248
use NAND2X1  _14043_
timestamp 0
transform 1 0 10950 0 -1 13690
box -6 -8 86 248
use AOI21X1  _14044_
timestamp 0
transform -1 0 11010 0 -1 13210
box -6 -8 106 248
use NAND3X1  _14045_
timestamp 0
transform -1 0 10710 0 1 13210
box -6 -8 106 248
use NAND2X1  _14046_
timestamp 0
transform 1 0 10750 0 1 13210
box -6 -8 86 248
use AOI21X1  _14047_
timestamp 0
transform -1 0 10570 0 1 13210
box -6 -8 106 248
use OAI21X1  _14048_
timestamp 0
transform -1 0 10050 0 1 12250
box -6 -8 106 248
use INVX1  _14049_
timestamp 0
transform 1 0 10010 0 -1 12250
box -6 -8 66 248
use OR2X2  _14050_
timestamp 0
transform -1 0 9870 0 -1 12730
box -6 -8 106 248
use OAI21X1  _14051_
timestamp 0
transform -1 0 9650 0 1 12250
box -6 -8 106 248
use OAI22X1  _14052_
timestamp 0
transform -1 0 9950 0 -1 12250
box -6 -8 126 248
use NAND2X1  _14053_
timestamp 0
transform -1 0 9730 0 1 11770
box -6 -8 86 248
use NOR2X1  _14054_
timestamp 0
transform 1 0 9710 0 1 12250
box -6 -8 86 248
use NOR2X1  _14055_
timestamp 0
transform -1 0 9910 0 1 12250
box -6 -8 86 248
use OAI21X1  _14056_
timestamp 0
transform 1 0 10490 0 1 13690
box -6 -8 106 248
use INVX1  _14057_
timestamp 0
transform -1 0 9890 0 1 12730
box -6 -8 66 248
use OAI21X1  _14058_
timestamp 0
transform 1 0 10750 0 -1 13210
box -6 -8 106 248
use NAND2X1  _14059_
timestamp 0
transform -1 0 10030 0 1 12730
box -6 -8 86 248
use OR2X2  _14060_
timestamp 0
transform -1 0 10550 0 -1 12730
box -6 -8 106 248
use NAND3X1  _14061_
timestamp 0
transform 1 0 10310 0 -1 12730
box -6 -8 106 248
use NAND2X1  _14062_
timestamp 0
transform 1 0 10170 0 -1 12730
box -6 -8 86 248
use NAND2X1  _14063_
timestamp 0
transform 1 0 10050 0 -1 12730
box -6 -8 86 248
use NAND2X1  _14064_
timestamp 0
transform -1 0 10810 0 -1 12250
box -6 -8 86 248
use AND2X2  _14065_
timestamp 0
transform 1 0 10470 0 1 11770
box -6 -8 106 248
use OAI21X1  _14066_
timestamp 0
transform -1 0 10430 0 1 11770
box -6 -8 106 248
use OAI21X1  _14067_
timestamp 0
transform -1 0 10270 0 1 11770
box -6 -8 106 248
use INVX1  _14068_
timestamp 0
transform 1 0 9390 0 1 11770
box -6 -8 66 248
use INVX1  _14069_
timestamp 0
transform 1 0 10850 0 -1 12250
box -6 -8 66 248
use AOI21X1  _14070_
timestamp 0
transform -1 0 10730 0 1 12250
box -6 -8 106 248
use NOR2X1  _14071_
timestamp 0
transform -1 0 10170 0 1 12250
box -6 -8 86 248
use NAND3X1  _14072_
timestamp 0
transform -1 0 10310 0 1 12250
box -6 -8 106 248
use OAI21X1  _14073_
timestamp 0
transform 1 0 10590 0 -1 12250
box -6 -8 106 248
use OAI21X1  _14074_
timestamp 0
transform 1 0 10470 0 -1 14170
box -6 -8 106 248
use INVX1  _14075_
timestamp 0
transform 1 0 10510 0 -1 13690
box -6 -8 66 248
use OR2X2  _14076_
timestamp 0
transform -1 0 10710 0 -1 13210
box -6 -8 106 248
use OAI21X1  _14077_
timestamp 0
transform -1 0 10470 0 -1 13210
box -6 -8 106 248
use NAND2X1  _14078_
timestamp 0
transform 1 0 10150 0 -1 13210
box -6 -8 86 248
use OR2X2  _14079_
timestamp 0
transform -1 0 9210 0 1 12730
box -6 -8 106 248
use NAND3X1  _14080_
timestamp 0
transform -1 0 9790 0 1 12730
box -6 -8 106 248
use AND2X2  _14081_
timestamp 0
transform 1 0 9390 0 1 12730
box -6 -8 106 248
use NOR2X1  _14082_
timestamp 0
transform -1 0 9350 0 1 12730
box -6 -8 86 248
use OAI21X1  _14083_
timestamp 0
transform 1 0 9530 0 1 12730
box -6 -8 106 248
use NAND2X1  _14084_
timestamp 0
transform 1 0 10450 0 -1 12250
box -6 -8 86 248
use AND2X2  _14085_
timestamp 0
transform -1 0 10190 0 -1 11770
box -6 -8 106 248
use NOR2X1  _14086_
timestamp 0
transform 1 0 10230 0 -1 11770
box -6 -8 86 248
use NOR2X1  _14087_
timestamp 0
transform -1 0 10030 0 -1 11770
box -6 -8 86 248
use AOI22X1  _14088_
timestamp 0
transform 1 0 9490 0 1 11770
box -6 -8 126 248
use NAND2X1  _14089_
timestamp 0
transform 1 0 9290 0 -1 11770
box -6 -8 86 248
use INVX1  _14090_
timestamp 0
transform 1 0 11110 0 -1 12250
box -6 -8 66 248
use AOI21X1  _14091_
timestamp 0
transform 1 0 10950 0 -1 12250
box -6 -8 106 248
use NAND2X1  _14092_
timestamp 0
transform 1 0 10090 0 1 13210
box -6 -8 86 248
use NOR2X1  _14093_
timestamp 0
transform 1 0 10010 0 -1 13210
box -6 -8 86 248
use AOI21X1  _14094_
timestamp 0
transform -1 0 10030 0 1 13210
box -6 -8 106 248
use NOR2X1  _14095_
timestamp 0
transform 1 0 9890 0 -1 13210
box -6 -8 86 248
use AND2X2  _14096_
timestamp 0
transform -1 0 9890 0 -1 11770
box -6 -8 106 248
use OAI21X1  _14097_
timestamp 0
transform -1 0 9890 0 1 11770
box -6 -8 106 248
use OAI21X1  _14098_
timestamp 0
transform -1 0 9750 0 -1 11770
box -6 -8 106 248
use NAND2X1  _14099_
timestamp 0
transform 1 0 8810 0 -1 11770
box -6 -8 86 248
use NAND2X1  _14100_
timestamp 0
transform 1 0 8450 0 1 12250
box -6 -8 86 248
use NOR2X1  _14101_
timestamp 0
transform 1 0 8810 0 1 12730
box -6 -8 86 248
use NAND2X1  _14102_
timestamp 0
transform -1 0 10430 0 -1 14170
box -6 -8 86 248
use OAI21X1  _14103_
timestamp 0
transform 1 0 10330 0 1 13690
box -6 -8 106 248
use NAND2X1  _14104_
timestamp 0
transform -1 0 9790 0 -1 14170
box -6 -8 86 248
use OAI21X1  _14105_
timestamp 0
transform -1 0 9930 0 -1 14170
box -6 -8 106 248
use INVX1  _14106_
timestamp 0
transform -1 0 9650 0 -1 14170
box -6 -8 66 248
use OR2X2  _14107_
timestamp 0
transform -1 0 9610 0 -1 13210
box -6 -8 106 248
use OAI21X1  _14108_
timestamp 0
transform 1 0 9610 0 1 13210
box -6 -8 106 248
use OAI21X1  _14109_
timestamp 0
transform 1 0 9770 0 1 13210
box -6 -8 106 248
use INVX1  _14110_
timestamp 0
transform -1 0 9930 0 -1 13690
box -6 -8 66 248
use OAI21X1  _14111_
timestamp 0
transform 1 0 9370 0 -1 13210
box -6 -8 106 248
use OAI21X1  _14112_
timestamp 0
transform 1 0 9210 0 -1 13210
box -6 -8 106 248
use NAND2X1  _14113_
timestamp 0
transform 1 0 7630 0 1 12250
box -6 -8 86 248
use NAND2X1  _14114_
timestamp 0
transform 1 0 9450 0 1 14170
box -6 -8 86 248
use OAI21X1  _14115_
timestamp 0
transform 1 0 9310 0 1 14170
box -6 -8 106 248
use NAND2X1  _14116_
timestamp 0
transform -1 0 9690 0 -1 13690
box -6 -8 86 248
use OAI21X1  _14117_
timestamp 0
transform 1 0 9730 0 -1 13690
box -6 -8 106 248
use AND2X2  _14118_
timestamp 0
transform -1 0 7990 0 1 12250
box -6 -8 106 248
use NAND2X1  _14119_
timestamp 0
transform -1 0 10230 0 -1 15610
box -6 -8 86 248
use OAI21X1  _14120_
timestamp 0
transform -1 0 10290 0 1 15610
box -6 -8 106 248
use NAND2X1  _14121_
timestamp 0
transform 1 0 9890 0 -1 15610
box -6 -8 86 248
use OAI21X1  _14122_
timestamp 0
transform 1 0 9730 0 -1 15610
box -6 -8 106 248
use OAI21X1  _14123_
timestamp 0
transform -1 0 8550 0 -1 14650
box -6 -8 106 248
use OAI21X1  _14124_
timestamp 0
transform -1 0 8670 0 1 14170
box -6 -8 106 248
use OAI21X1  _14125_
timestamp 0
transform 1 0 8150 0 -1 13210
box -6 -8 106 248
use OAI21X1  _14126_
timestamp 0
transform -1 0 8630 0 -1 13210
box -6 -8 106 248
use NAND2X1  _14127_
timestamp 0
transform 1 0 8670 0 1 15130
box -6 -8 86 248
use OAI21X1  _14128_
timestamp 0
transform -1 0 8630 0 1 15130
box -6 -8 106 248
use NAND2X1  _14129_
timestamp 0
transform 1 0 9190 0 -1 15610
box -6 -8 86 248
use OAI21X1  _14130_
timestamp 0
transform 1 0 9050 0 -1 15610
box -6 -8 106 248
use NAND2X1  _14131_
timestamp 0
transform -1 0 10310 0 -1 14170
box -6 -8 86 248
use OAI21X1  _14132_
timestamp 0
transform 1 0 10190 0 1 13690
box -6 -8 106 248
use NAND2X1  _14133_
timestamp 0
transform -1 0 11030 0 1 14170
box -6 -8 86 248
use OAI21X1  _14134_
timestamp 0
transform 1 0 10810 0 1 14170
box -6 -8 106 248
use INVX1  _14135_
timestamp 0
transform -1 0 8530 0 1 14170
box -6 -8 66 248
use OAI21X1  _14136_
timestamp 0
transform -1 0 9310 0 1 13210
box -6 -8 106 248
use OAI21X1  _14137_
timestamp 0
transform 1 0 9070 0 1 13210
box -6 -8 106 248
use INVX1  _14138_
timestamp 0
transform 1 0 7950 0 1 14170
box -6 -8 66 248
use OAI21X1  _14139_
timestamp 0
transform -1 0 9170 0 -1 13210
box -6 -8 106 248
use OAI21X1  _14140_
timestamp 0
transform 1 0 8930 0 -1 13210
box -6 -8 106 248
use NAND2X1  _14141_
timestamp 0
transform 1 0 7710 0 1 14170
box -6 -8 86 248
use OAI21X1  _14142_
timestamp 0
transform 1 0 7670 0 -1 14170
box -6 -8 106 248
use NAND2X1  _14143_
timestamp 0
transform 1 0 7830 0 1 14170
box -6 -8 86 248
use OAI21X1  _14144_
timestamp 0
transform -1 0 7930 0 -1 14170
box -6 -8 106 248
use NAND2X1  _14145_
timestamp 0
transform -1 0 6650 0 1 15610
box -6 -8 86 248
use OAI21X1  _14146_
timestamp 0
transform 1 0 6430 0 1 15610
box -6 -8 106 248
use NAND2X1  _14147_
timestamp 0
transform 1 0 7590 0 -1 15130
box -6 -8 86 248
use OAI21X1  _14148_
timestamp 0
transform 1 0 7170 0 -1 15130
box -6 -8 106 248
use OAI21X1  _14149_
timestamp 0
transform -1 0 7590 0 -1 14650
box -6 -8 106 248
use OAI21X1  _14150_
timestamp 0
transform -1 0 7670 0 1 14170
box -6 -8 106 248
use OAI21X1  _14151_
timestamp 0
transform -1 0 7730 0 1 13210
box -6 -8 106 248
use OAI21X1  _14152_
timestamp 0
transform -1 0 7870 0 1 13210
box -6 -8 106 248
use NAND2X1  _14153_
timestamp 0
transform 1 0 7190 0 -1 15610
box -6 -8 86 248
use OAI21X1  _14154_
timestamp 0
transform -1 0 7090 0 1 15610
box -6 -8 106 248
use NAND2X1  _14155_
timestamp 0
transform 1 0 7450 0 -1 15130
box -6 -8 86 248
use OAI21X1  _14156_
timestamp 0
transform 1 0 7290 0 1 15610
box -6 -8 106 248
use NAND2X1  _14157_
timestamp 0
transform -1 0 11170 0 -1 14170
box -6 -8 86 248
use OAI21X1  _14158_
timestamp 0
transform 1 0 10950 0 -1 14170
box -6 -8 106 248
use DFFPOSX1  _14159_
timestamp 0
transform -1 0 7630 0 -1 13690
box -6 -8 246 248
use DFFPOSX1  _14160_
timestamp 0
transform 1 0 6370 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _14161_
timestamp 0
transform 1 0 8730 0 1 10810
box -6 -8 246 248
use DFFPOSX1  _14162_
timestamp 0
transform 1 0 6750 0 -1 13210
box -6 -8 246 248
use DFFPOSX1  _14163_
timestamp 0
transform 1 0 6610 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _14164_
timestamp 0
transform 1 0 6110 0 -1 13210
box -6 -8 246 248
use DFFPOSX1  _14165_
timestamp 0
transform 1 0 7410 0 1 11770
box -6 -8 246 248
use DFFPOSX1  _14166_
timestamp 0
transform 1 0 6130 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _14167_
timestamp 0
transform 1 0 7150 0 -1 12250
box -6 -8 246 248
use DFFPOSX1  _14168_
timestamp 0
transform 1 0 6830 0 1 12730
box -6 -8 246 248
use DFFPOSX1  _14169_
timestamp 0
transform 1 0 7310 0 1 11290
box -6 -8 246 248
use DFFPOSX1  _14170_
timestamp 0
transform -1 0 7470 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _14171_
timestamp 0
transform 1 0 7930 0 -1 12250
box -6 -8 246 248
use DFFPOSX1  _14172_
timestamp 0
transform -1 0 8770 0 1 13210
box -6 -8 246 248
use DFFPOSX1  _14173_
timestamp 0
transform -1 0 9210 0 -1 12250
box -6 -8 246 248
use DFFPOSX1  _14174_
timestamp 0
transform 1 0 7230 0 1 12730
box -6 -8 246 248
use DFFPOSX1  _14175_
timestamp 0
transform 1 0 8410 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _14176_
timestamp 0
transform -1 0 9790 0 -1 12250
box -6 -8 246 248
use DFFPOSX1  _14177_
timestamp 0
transform -1 0 9070 0 1 12250
box -6 -8 246 248
use DFFPOSX1  _14178_
timestamp 0
transform -1 0 9490 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _14179_
timestamp 0
transform -1 0 9010 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _14180_
timestamp 0
transform -1 0 10410 0 -1 12250
box -6 -8 246 248
use DFFPOSX1  _14181_
timestamp 0
transform -1 0 10130 0 1 11770
box -6 -8 246 248
use DFFPOSX1  _14182_
timestamp 0
transform -1 0 9250 0 -1 11770
box -6 -8 246 248
use DFFPOSX1  _14183_
timestamp 0
transform -1 0 9610 0 -1 11770
box -6 -8 246 248
use DFFPOSX1  _14184_
timestamp 0
transform -1 0 10810 0 -1 13690
box -6 -8 246 248
use DFFPOSX1  _14185_
timestamp 0
transform 1 0 9770 0 1 14170
box -6 -8 246 248
use DFFPOSX1  _14186_
timestamp 0
transform 1 0 10170 0 1 13210
box -6 -8 246 248
use DFFPOSX1  _14187_
timestamp 0
transform 1 0 8390 0 1 12730
box -6 -8 246 248
use DFFPOSX1  _14188_
timestamp 0
transform 1 0 9030 0 1 14170
box -6 -8 246 248
use DFFPOSX1  _14189_
timestamp 0
transform 1 0 10210 0 -1 13690
box -6 -8 246 248
use DFFPOSX1  _14190_
timestamp 0
transform -1 0 10530 0 1 15610
box -6 -8 246 248
use DFFPOSX1  _14191_
timestamp 0
transform -1 0 9690 0 -1 15610
box -6 -8 246 248
use DFFPOSX1  _14192_
timestamp 0
transform 1 0 8670 0 1 14170
box -6 -8 246 248
use DFFPOSX1  _14193_
timestamp 0
transform -1 0 8490 0 -1 13210
box -6 -8 246 248
use DFFPOSX1  _14194_
timestamp 0
transform -1 0 8470 0 1 15130
box -6 -8 246 248
use DFFPOSX1  _14195_
timestamp 0
transform -1 0 8790 0 1 15610
box -6 -8 246 248
use DFFPOSX1  _14196_
timestamp 0
transform -1 0 10130 0 1 13690
box -6 -8 246 248
use DFFPOSX1  _14197_
timestamp 0
transform -1 0 10770 0 1 14170
box -6 -8 246 248
use DFFPOSX1  _14198_
timestamp 0
transform -1 0 9010 0 1 13210
box -6 -8 246 248
use DFFPOSX1  _14199_
timestamp 0
transform 1 0 8630 0 -1 13210
box -6 -8 246 248
use DFFPOSX1  _14200_
timestamp 0
transform -1 0 7370 0 -1 14170
box -6 -8 246 248
use DFFPOSX1  _14201_
timestamp 0
transform -1 0 7610 0 -1 14170
box -6 -8 246 248
use DFFPOSX1  _14202_
timestamp 0
transform -1 0 6030 0 -1 16090
box -6 -8 246 248
use DFFPOSX1  _14203_
timestamp 0
transform -1 0 7310 0 1 15130
box -6 -8 246 248
use DFFPOSX1  _14204_
timestamp 0
transform -1 0 7530 0 1 14170
box -6 -8 246 248
use DFFPOSX1  _14205_
timestamp 0
transform -1 0 7270 0 1 13210
box -6 -8 246 248
use DFFPOSX1  _14206_
timestamp 0
transform -1 0 7030 0 -1 16090
box -6 -8 246 248
use DFFPOSX1  _14207_
timestamp 0
transform -1 0 7390 0 -1 16090
box -6 -8 246 248
use DFFPOSX1  _14208_
timestamp 0
transform -1 0 10910 0 -1 14170
box -6 -8 246 248
use DFFPOSX1  _14209_
timestamp 0
transform -1 0 9250 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _14210_
timestamp 0
transform 1 0 7710 0 -1 12730
box -6 -8 246 248
use DFFPOSX1  _14211_
timestamp 0
transform 1 0 8170 0 -1 12250
box -6 -8 246 248
use DFFPOSX1  _14212_
timestamp 0
transform -1 0 8710 0 1 11770
box -6 -8 246 248
use DFFPOSX1  _14213_
timestamp 0
transform -1 0 8510 0 -1 11770
box -6 -8 246 248
use DFFPOSX1  _14214_
timestamp 0
transform 1 0 8030 0 -1 11770
box -6 -8 246 248
use DFFPOSX1  _14215_
timestamp 0
transform 1 0 8510 0 -1 11770
box -6 -8 246 248
use INVX1  _14216_
timestamp 0
transform 1 0 7510 0 -1 6970
box -6 -8 66 248
use NAND2X1  _14217_
timestamp 0
transform 1 0 7710 0 -1 7450
box -6 -8 86 248
use OAI21X1  _14218_
timestamp 0
transform -1 0 7830 0 1 6970
box -6 -8 106 248
use INVX1  _14219_
timestamp 0
transform -1 0 7590 0 1 8410
box -6 -8 66 248
use NAND2X1  _14220_
timestamp 0
transform 1 0 7690 0 1 7930
box -6 -8 86 248
use OAI21X1  _14221_
timestamp 0
transform 1 0 7530 0 1 7930
box -6 -8 106 248
use INVX1  _14222_
timestamp 0
transform -1 0 7490 0 1 7450
box -6 -8 66 248
use NAND2X1  _14223_
timestamp 0
transform -1 0 7010 0 1 6970
box -6 -8 86 248
use OAI21X1  _14224_
timestamp 0
transform 1 0 7050 0 1 6970
box -6 -8 106 248
use INVX1  _14225_
timestamp 0
transform 1 0 6870 0 -1 6970
box -6 -8 66 248
use NAND2X1  _14226_
timestamp 0
transform -1 0 7290 0 -1 7450
box -6 -8 86 248
use OAI21X1  _14227_
timestamp 0
transform 1 0 7190 0 1 6970
box -6 -8 106 248
use INVX1  _14228_
timestamp 0
transform -1 0 8610 0 -1 6490
box -6 -8 66 248
use NAND2X1  _14229_
timestamp 0
transform 1 0 7970 0 -1 6970
box -6 -8 86 248
use OAI21X1  _14230_
timestamp 0
transform -1 0 8490 0 -1 6490
box -6 -8 106 248
use INVX1  _14231_
timestamp 0
transform -1 0 10290 0 -1 7450
box -6 -8 66 248
use NAND2X1  _14232_
timestamp 0
transform -1 0 10050 0 -1 7450
box -6 -8 86 248
use OAI21X1  _14233_
timestamp 0
transform -1 0 10190 0 -1 7450
box -6 -8 106 248
use INVX1  _14234_
timestamp 0
transform -1 0 9050 0 1 6490
box -6 -8 66 248
use NAND2X1  _14235_
timestamp 0
transform 1 0 8570 0 -1 6970
box -6 -8 86 248
use OAI21X1  _14236_
timestamp 0
transform 1 0 8450 0 1 6490
box -6 -8 106 248
use INVX1  _14237_
timestamp 0
transform -1 0 8950 0 1 6490
box -6 -8 66 248
use NAND2X1  _14238_
timestamp 0
transform -1 0 7970 0 1 6490
box -6 -8 86 248
use OAI21X1  _14239_
timestamp 0
transform -1 0 8130 0 1 6490
box -6 -8 106 248
use INVX1  _14240_
timestamp 0
transform -1 0 8510 0 -1 6970
box -6 -8 66 248
use NAND2X1  _14241_
timestamp 0
transform -1 0 8410 0 -1 6970
box -6 -8 86 248
use OAI21X1  _14242_
timestamp 0
transform -1 0 8410 0 1 6490
box -6 -8 106 248
use INVX1  _14243_
timestamp 0
transform -1 0 8430 0 1 7450
box -6 -8 66 248
use NAND2X1  _14244_
timestamp 0
transform 1 0 6930 0 1 7450
box -6 -8 86 248
use OAI21X1  _14245_
timestamp 0
transform -1 0 6870 0 1 7450
box -6 -8 106 248
use INVX1  _14246_
timestamp 0
transform 1 0 9490 0 1 6970
box -6 -8 66 248
use NAND2X1  _14247_
timestamp 0
transform 1 0 8750 0 1 6490
box -6 -8 86 248
use OAI21X1  _14248_
timestamp 0
transform 1 0 8590 0 1 6490
box -6 -8 106 248
use INVX1  _14249_
timestamp 0
transform 1 0 9850 0 -1 7450
box -6 -8 66 248
use NAND2X1  _14250_
timestamp 0
transform 1 0 10010 0 1 6970
box -6 -8 86 248
use OAI21X1  _14251_
timestamp 0
transform 1 0 9870 0 1 6970
box -6 -8 106 248
use INVX1  _14252_
timestamp 0
transform 1 0 7610 0 -1 10330
box -6 -8 66 248
use INVX8  _14253_
timestamp 0
transform 1 0 7830 0 -1 7450
box -6 -8 126 248
use NAND2X1  _14254_
timestamp 0
transform 1 0 7690 0 1 7450
box -6 -8 86 248
use OAI21X1  _14255_
timestamp 0
transform 1 0 7530 0 1 7450
box -6 -8 106 248
use NAND3X1  _14256_
timestamp 0
transform 1 0 7190 0 1 8890
box -6 -8 106 248
use INVX4  _14257_
timestamp 0
transform -1 0 8190 0 -1 8890
box -6 -8 86 248
use INVX1  _14258_
timestamp 0
transform 1 0 7070 0 -1 9370
box -6 -8 66 248
use OAI21X1  _14259_
timestamp 0
transform -1 0 7290 0 -1 9370
box -6 -8 106 248
use NAND2X1  _14260_
timestamp 0
transform 1 0 7330 0 1 8890
box -6 -8 86 248
use NAND2X1  _14261_
timestamp 0
transform 1 0 7770 0 -1 8410
box -6 -8 86 248
use OAI21X1  _14262_
timestamp 0
transform 1 0 7610 0 -1 8410
box -6 -8 106 248
use INVX1  _14263_
timestamp 0
transform -1 0 7890 0 1 8890
box -6 -8 66 248
use OAI21X1  _14264_
timestamp 0
transform 1 0 7030 0 1 8890
box -6 -8 106 248
use OR2X2  _14265_
timestamp 0
transform -1 0 7130 0 -1 8890
box -6 -8 106 248
use NOR2X1  _14266_
timestamp 0
transform -1 0 7030 0 -1 9370
box -6 -8 86 248
use OAI21X1  _14267_
timestamp 0
transform -1 0 7270 0 -1 8890
box -6 -8 106 248
use NAND2X1  _14268_
timestamp 0
transform -1 0 6990 0 -1 8890
box -6 -8 86 248
use NAND2X1  _14269_
timestamp 0
transform 1 0 7090 0 -1 7450
box -6 -8 86 248
use OAI21X1  _14270_
timestamp 0
transform 1 0 6950 0 -1 7450
box -6 -8 106 248
use OAI21X1  _14271_
timestamp 0
transform -1 0 7410 0 -1 8890
box -6 -8 106 248
use NAND2X1  _14272_
timestamp 0
transform -1 0 7530 0 -1 8890
box -6 -8 86 248
use OR2X2  _14273_
timestamp 0
transform 1 0 7590 0 -1 8890
box -6 -8 106 248
use NAND2X1  _14274_
timestamp 0
transform -1 0 7810 0 -1 8890
box -6 -8 86 248
use NAND2X1  _14275_
timestamp 0
transform 1 0 7310 0 1 7450
box -6 -8 86 248
use OAI21X1  _14276_
timestamp 0
transform -1 0 7810 0 -1 7930
box -6 -8 106 248
use NOR2X1  _14277_
timestamp 0
transform -1 0 8010 0 1 8890
box -6 -8 86 248
use NAND2X1  _14278_
timestamp 0
transform -1 0 8070 0 -1 8890
box -6 -8 86 248
use NAND3X1  _14279_
timestamp 0
transform 1 0 9330 0 -1 7930
box -6 -8 106 248
use INVX1  _14280_
timestamp 0
transform -1 0 9330 0 1 7930
box -6 -8 66 248
use AND2X2  _14281_
timestamp 0
transform 1 0 8050 0 1 8890
box -6 -8 106 248
use OAI21X1  _14282_
timestamp 0
transform -1 0 9490 0 1 7930
box -6 -8 106 248
use NAND2X1  _14283_
timestamp 0
transform 1 0 9470 0 -1 7930
box -6 -8 86 248
use NAND2X1  _14284_
timestamp 0
transform 1 0 8290 0 1 6970
box -6 -8 86 248
use OAI21X1  _14285_
timestamp 0
transform -1 0 8530 0 1 6970
box -6 -8 106 248
use INVX1  _14286_
timestamp 0
transform 1 0 8230 0 -1 7450
box -6 -8 66 248
use OAI21X1  _14287_
timestamp 0
transform -1 0 9290 0 -1 7930
box -6 -8 106 248
use NAND2X1  _14288_
timestamp 0
transform 1 0 8250 0 1 7450
box -6 -8 86 248
use NOR2X1  _14289_
timestamp 0
transform 1 0 8090 0 -1 7930
box -6 -8 86 248
use NOR2X1  _14290_
timestamp 0
transform 1 0 7970 0 1 7450
box -6 -8 86 248
use AOI22X1  _14291_
timestamp 0
transform -1 0 8210 0 1 7450
box -6 -8 126 248
use NOR2X1  _14292_
timestamp 0
transform -1 0 8290 0 1 8890
box -6 -8 86 248
use NAND2X1  _14293_
timestamp 0
transform 1 0 9230 0 1 8410
box -6 -8 86 248
use NAND3X1  _14294_
timestamp 0
transform -1 0 9350 0 -1 8410
box -6 -8 106 248
use INVX1  _14295_
timestamp 0
transform 1 0 8990 0 -1 8410
box -6 -8 66 248
use NAND2X1  _14296_
timestamp 0
transform 1 0 9110 0 1 8410
box -6 -8 86 248
use NAND2X1  _14297_
timestamp 0
transform 1 0 9110 0 -1 8410
box -6 -8 86 248
use NAND2X1  _14298_
timestamp 0
transform -1 0 9210 0 1 7930
box -6 -8 86 248
use NAND2X1  _14299_
timestamp 0
transform -1 0 8930 0 1 6970
box -6 -8 86 248
use OAI21X1  _14300_
timestamp 0
transform -1 0 9210 0 1 6970
box -6 -8 106 248
use INVX1  _14301_
timestamp 0
transform 1 0 7870 0 -1 6970
box -6 -8 66 248
use NAND3X1  _14302_
timestamp 0
transform -1 0 8950 0 -1 8410
box -6 -8 106 248
use NAND3X1  _14303_
timestamp 0
transform -1 0 8990 0 1 7930
box -6 -8 106 248
use INVX1  _14304_
timestamp 0
transform -1 0 9070 0 1 8410
box -6 -8 66 248
use NAND2X1  _14305_
timestamp 0
transform 1 0 8710 0 1 8410
box -6 -8 86 248
use NAND3X1  _14306_
timestamp 0
transform -1 0 8950 0 1 8410
box -6 -8 106 248
use NAND3X1  _14307_
timestamp 0
transform 1 0 8750 0 1 7930
box -6 -8 106 248
use OAI21X1  _14308_
timestamp 0
transform 1 0 8150 0 1 6970
box -6 -8 106 248
use INVX1  _14309_
timestamp 0
transform 1 0 9410 0 -1 8410
box -6 -8 66 248
use NOR2X1  _14310_
timestamp 0
transform -1 0 8410 0 1 8890
box -6 -8 86 248
use NAND2X1  _14311_
timestamp 0
transform -1 0 8450 0 -1 8890
box -6 -8 86 248
use OAI21X1  _14312_
timestamp 0
transform 1 0 8490 0 -1 8890
box -6 -8 106 248
use OR2X2  _14313_
timestamp 0
transform -1 0 9770 0 1 7930
box -6 -8 106 248
use NAND2X1  _14314_
timestamp 0
transform -1 0 9610 0 1 7930
box -6 -8 86 248
use NAND2X1  _14315_
timestamp 0
transform 1 0 9590 0 -1 7930
box -6 -8 86 248
use NAND2X1  _14316_
timestamp 0
transform 1 0 8710 0 1 6970
box -6 -8 86 248
use OAI21X1  _14317_
timestamp 0
transform -1 0 8790 0 -1 7450
box -6 -8 106 248
use INVX1  _14318_
timestamp 0
transform 1 0 8470 0 -1 7930
box -6 -8 66 248
use INVX1  _14319_
timestamp 0
transform -1 0 9090 0 1 7930
box -6 -8 66 248
use OAI21X1  _14320_
timestamp 0
transform -1 0 9830 0 -1 7930
box -6 -8 106 248
use OR2X2  _14321_
timestamp 0
transform -1 0 8850 0 -1 7930
box -6 -8 106 248
use AOI21X1  _14322_
timestamp 0
transform -1 0 8990 0 -1 7930
box -6 -8 106 248
use AOI22X1  _14323_
timestamp 0
transform 1 0 8590 0 -1 7930
box -6 -8 126 248
use INVX1  _14324_
timestamp 0
transform 1 0 8930 0 -1 6970
box -6 -8 66 248
use AND2X2  _14325_
timestamp 0
transform 1 0 8470 0 1 8890
box -6 -8 106 248
use NOR2X1  _14326_
timestamp 0
transform -1 0 8710 0 -1 8890
box -6 -8 86 248
use NAND3X1  _14327_
timestamp 0
transform 1 0 8730 0 1 8890
box -6 -8 106 248
use NAND3X1  _14328_
timestamp 0
transform 1 0 8890 0 1 8890
box -6 -8 106 248
use INVX1  _14329_
timestamp 0
transform -1 0 8870 0 1 9370
box -6 -8 66 248
use NAND2X1  _14330_
timestamp 0
transform 1 0 9050 0 1 8890
box -6 -8 86 248
use NAND2X1  _14331_
timestamp 0
transform -1 0 9250 0 1 8890
box -6 -8 86 248
use NAND3X1  _14332_
timestamp 0
transform -1 0 9410 0 1 8890
box -6 -8 106 248
use OAI21X1  _14333_
timestamp 0
transform 1 0 8970 0 1 6970
box -6 -8 106 248
use NAND2X1  _14334_
timestamp 0
transform -1 0 9790 0 -1 7450
box -6 -8 86 248
use INVX1  _14335_
timestamp 0
transform -1 0 8730 0 1 10810
box -6 -8 66 248
use NAND2X1  _14336_
timestamp 0
transform 1 0 8530 0 1 10810
box -6 -8 86 248
use INVX1  _14337_
timestamp 0
transform -1 0 8490 0 1 10810
box -6 -8 66 248
use NAND2X1  _14338_
timestamp 0
transform 1 0 8870 0 -1 10810
box -6 -8 86 248
use NAND2X1  _14339_
timestamp 0
transform 1 0 9030 0 1 10330
box -6 -8 86 248
use INVX1  _14340_
timestamp 0
transform -1 0 9090 0 1 9370
box -6 -8 66 248
use NAND2X1  _14341_
timestamp 0
transform -1 0 8950 0 -1 9370
box -6 -8 86 248
use NAND3X1  _14342_
timestamp 0
transform 1 0 9170 0 -1 9370
box -6 -8 106 248
use OAI21X1  _14343_
timestamp 0
transform 1 0 8730 0 -1 9370
box -6 -8 106 248
use NAND3X1  _14344_
timestamp 0
transform 1 0 9010 0 -1 9370
box -6 -8 106 248
use NAND2X1  _14345_
timestamp 0
transform 1 0 9310 0 -1 9370
box -6 -8 86 248
use NAND3X1  _14346_
timestamp 0
transform 1 0 9430 0 -1 9370
box -6 -8 106 248
use NAND2X1  _14347_
timestamp 0
transform -1 0 9670 0 -1 7450
box -6 -8 86 248
use NAND2X1  _14348_
timestamp 0
transform 1 0 8030 0 1 6970
box -6 -8 86 248
use OAI21X1  _14349_
timestamp 0
transform 1 0 7890 0 1 6970
box -6 -8 106 248
use NAND3X1  _14350_
timestamp 0
transform -1 0 8270 0 1 8410
box -6 -8 106 248
use INVX1  _14351_
timestamp 0
transform -1 0 7770 0 1 8890
box -6 -8 66 248
use INVX1  _14352_
timestamp 0
transform -1 0 7510 0 1 8890
box -6 -8 66 248
use OAI21X1  _14353_
timestamp 0
transform -1 0 7650 0 1 8890
box -6 -8 106 248
use NAND3X1  _14354_
timestamp 0
transform -1 0 8130 0 1 8410
box -6 -8 106 248
use OAI21X1  _14355_
timestamp 0
transform 1 0 7870 0 1 8410
box -6 -8 106 248
use INVX1  _14356_
timestamp 0
transform 1 0 8330 0 -1 8410
box -6 -8 66 248
use OAI21X1  _14357_
timestamp 0
transform -1 0 8410 0 1 8410
box -6 -8 106 248
use OR2X2  _14358_
timestamp 0
transform 1 0 8330 0 1 7930
box -6 -8 106 248
use NOR2X1  _14359_
timestamp 0
transform 1 0 8470 0 1 8410
box -6 -8 86 248
use OAI21X1  _14360_
timestamp 0
transform -1 0 8530 0 -1 8410
box -6 -8 106 248
use NAND3X1  _14361_
timestamp 0
transform 1 0 8490 0 1 7930
box -6 -8 106 248
use OAI21X1  _14362_
timestamp 0
transform 1 0 7570 0 -1 7450
box -6 -8 106 248
use OAI21X1  _14363_
timestamp 0
transform 1 0 8170 0 -1 8410
box -6 -8 106 248
use NAND2X1  _14364_
timestamp 0
transform -1 0 8110 0 -1 8410
box -6 -8 86 248
use OR2X2  _14365_
timestamp 0
transform -1 0 7990 0 -1 8410
box -6 -8 106 248
use NAND3X1  _14366_
timestamp 0
transform 1 0 8070 0 1 7930
box -6 -8 106 248
use OAI21X1  _14367_
timestamp 0
transform 1 0 7330 0 1 6970
box -6 -8 106 248
use INVX1  _14368_
timestamp 0
transform -1 0 9490 0 -1 8890
box -6 -8 66 248
use NOR2X1  _14369_
timestamp 0
transform 1 0 8590 0 1 8410
box -6 -8 86 248
use NAND2X1  _14370_
timestamp 0
transform 1 0 8570 0 -1 8410
box -6 -8 86 248
use NAND2X1  _14371_
timestamp 0
transform -1 0 9750 0 -1 8410
box -6 -8 86 248
use OR2X2  _14372_
timestamp 0
transform -1 0 10930 0 -1 7930
box -6 -8 106 248
use AND2X2  _14373_
timestamp 0
transform 1 0 8710 0 -1 8410
box -6 -8 106 248
use OAI21X1  _14374_
timestamp 0
transform 1 0 10370 0 1 7930
box -6 -8 106 248
use NAND3X1  _14375_
timestamp 0
transform 1 0 10410 0 -1 7930
box -6 -8 106 248
use OAI21X1  _14376_
timestamp 0
transform 1 0 8890 0 -1 6490
box -6 -8 106 248
use INVX1  _14377_
timestamp 0
transform 1 0 10010 0 -1 8890
box -6 -8 66 248
use OAI21X1  _14378_
timestamp 0
transform 1 0 10990 0 -1 7930
box -6 -8 106 248
use OR2X2  _14379_
timestamp 0
transform 1 0 11290 0 -1 7930
box -6 -8 106 248
use AOI21X1  _14380_
timestamp 0
transform -1 0 11250 0 -1 7930
box -6 -8 106 248
use AOI22X1  _14381_
timestamp 0
transform 1 0 11050 0 1 7450
box -6 -8 126 248
use NOR2X1  _14382_
timestamp 0
transform 1 0 9550 0 -1 8890
box -6 -8 86 248
use NAND2X1  _14383_
timestamp 0
transform -1 0 10290 0 -1 8410
box -6 -8 86 248
use NAND3X1  _14384_
timestamp 0
transform 1 0 10510 0 1 7930
box -6 -8 106 248
use INVX1  _14385_
timestamp 0
transform 1 0 10750 0 1 8410
box -6 -8 66 248
use NAND2X1  _14386_
timestamp 0
transform -1 0 10870 0 1 7930
box -6 -8 86 248
use NAND2X1  _14387_
timestamp 0
transform 1 0 10670 0 1 7930
box -6 -8 86 248
use NAND3X1  _14388_
timestamp 0
transform -1 0 10650 0 -1 7930
box -6 -8 106 248
use OAI21X1  _14389_
timestamp 0
transform 1 0 9090 0 1 6490
box -6 -8 106 248
use NAND3X1  _14390_
timestamp 0
transform -1 0 10450 0 -1 8410
box -6 -8 106 248
use NAND3X1  _14391_
timestamp 0
transform 1 0 10490 0 -1 8410
box -6 -8 106 248
use INVX1  _14392_
timestamp 0
transform 1 0 10650 0 -1 8410
box -6 -8 66 248
use NAND2X1  _14393_
timestamp 0
transform 1 0 11070 0 1 7930
box -6 -8 86 248
use NAND3X1  _14394_
timestamp 0
transform -1 0 11030 0 1 7930
box -6 -8 106 248
use NAND3X1  _14395_
timestamp 0
transform 1 0 10690 0 -1 7930
box -6 -8 106 248
use OAI21X1  _14396_
timestamp 0
transform 1 0 9590 0 1 6970
box -6 -8 106 248
use INVX1  _14397_
timestamp 0
transform 1 0 9810 0 -1 8410
box -6 -8 66 248
use NOR2X1  _14398_
timestamp 0
transform -1 0 10050 0 1 8890
box -6 -8 86 248
use NAND2X1  _14399_
timestamp 0
transform 1 0 10610 0 1 8410
box -6 -8 86 248
use OAI21X1  _14400_
timestamp 0
transform -1 0 10110 0 1 8410
box -6 -8 106 248
use OR2X2  _14401_
timestamp 0
transform 1 0 10010 0 -1 7930
box -6 -8 106 248
use NAND2X1  _14402_
timestamp 0
transform 1 0 10110 0 1 7930
box -6 -8 86 248
use NAND2X1  _14403_
timestamp 0
transform 1 0 10150 0 -1 7930
box -6 -8 86 248
use NAND2X1  _14404_
timestamp 0
transform -1 0 9050 0 -1 7450
box -6 -8 86 248
use OAI21X1  _14405_
timestamp 0
transform -1 0 9270 0 1 7450
box -6 -8 106 248
use INVX1  _14406_
timestamp 0
transform 1 0 10290 0 -1 7930
box -6 -8 66 248
use OAI21X1  _14407_
timestamp 0
transform 1 0 9870 0 -1 7930
box -6 -8 106 248
use OR2X2  _14408_
timestamp 0
transform -1 0 8970 0 1 7450
box -6 -8 106 248
use AOI21X1  _14409_
timestamp 0
transform -1 0 9130 0 1 7450
box -6 -8 106 248
use AOI22X1  _14410_
timestamp 0
transform 1 0 8710 0 1 7450
box -6 -8 126 248
use AND2X2  _14411_
timestamp 0
transform -1 0 10550 0 1 8410
box -6 -8 106 248
use NOR2X1  _14412_
timestamp 0
transform 1 0 10150 0 1 8410
box -6 -8 86 248
use NAND3X1  _14413_
timestamp 0
transform 1 0 10290 0 1 8410
box -6 -8 106 248
use NAND3X1  _14414_
timestamp 0
transform 1 0 9110 0 -1 8890
box -6 -8 106 248
use INVX1  _14415_
timestamp 0
transform 1 0 8910 0 1 9370
box -6 -8 66 248
use NAND2X1  _14416_
timestamp 0
transform 1 0 9890 0 1 8410
box -6 -8 86 248
use NAND2X1  _14417_
timestamp 0
transform 1 0 9450 0 1 8890
box -6 -8 86 248
use NAND3X1  _14418_
timestamp 0
transform -1 0 9370 0 -1 8890
box -6 -8 106 248
use OAI21X1  _14419_
timestamp 0
transform -1 0 9530 0 1 7450
box -6 -8 106 248
use NAND2X1  _14420_
timestamp 0
transform 1 0 9810 0 1 7450
box -6 -8 86 248
use INVX1  _14421_
timestamp 0
transform -1 0 8250 0 1 10810
box -6 -8 66 248
use NAND2X1  _14422_
timestamp 0
transform -1 0 8370 0 1 10810
box -6 -8 86 248
use NAND2X1  _14423_
timestamp 0
transform 1 0 9010 0 -1 10810
box -6 -8 86 248
use NAND2X1  _14424_
timestamp 0
transform 1 0 9290 0 1 10330
box -6 -8 86 248
use INVX1  _14425_
timestamp 0
transform 1 0 9630 0 1 8410
box -6 -8 66 248
use NAND2X1  _14426_
timestamp 0
transform -1 0 9070 0 -1 8890
box -6 -8 86 248
use NAND3X1  _14427_
timestamp 0
transform 1 0 9730 0 1 8410
box -6 -8 106 248
use OAI21X1  _14428_
timestamp 0
transform -1 0 10170 0 -1 8410
box -6 -8 106 248
use NAND3X1  _14429_
timestamp 0
transform -1 0 10010 0 -1 8410
box -6 -8 106 248
use NAND2X1  _14430_
timestamp 0
transform 1 0 9830 0 1 7930
box -6 -8 86 248
use NAND3X1  _14431_
timestamp 0
transform -1 0 10050 0 1 7930
box -6 -8 106 248
use NAND2X1  _14432_
timestamp 0
transform 1 0 9930 0 1 7450
box -6 -8 86 248
use INVX2  _14433_
timestamp 0
transform 1 0 8070 0 1 10330
box -6 -8 66 248
use NOR2X1  _14434_
timestamp 0
transform -1 0 8490 0 1 10330
box -6 -8 86 248
use AND2X2  _14435_
timestamp 0
transform 1 0 8530 0 -1 10330
box -6 -8 106 248
use INVX1  _14436_
timestamp 0
transform 1 0 7910 0 1 10810
box -6 -8 66 248
use NAND2X1  _14437_
timestamp 0
transform -1 0 8230 0 -1 10810
box -6 -8 86 248
use NOR2X1  _14438_
timestamp 0
transform -1 0 8450 0 -1 10810
box -6 -8 86 248
use AND2X2  _14439_
timestamp 0
transform 1 0 8490 0 -1 10810
box -6 -8 106 248
use NAND2X1  _14440_
timestamp 0
transform 1 0 9170 0 1 10330
box -6 -8 86 248
use OAI21X1  _14441_
timestamp 0
transform -1 0 9250 0 -1 10330
box -6 -8 106 248
use NAND2X1  _14442_
timestamp 0
transform 1 0 8350 0 -1 11290
box -6 -8 86 248
use OAI21X1  _14443_
timestamp 0
transform -1 0 8570 0 -1 11290
box -6 -8 106 248
use INVX1  _14444_
timestamp 0
transform 1 0 9050 0 -1 10330
box -6 -8 66 248
use NOR2X1  _14445_
timestamp 0
transform -1 0 8850 0 1 10330
box -6 -8 86 248
use NAND2X1  _14446_
timestamp 0
transform 1 0 8910 0 -1 10330
box -6 -8 86 248
use NAND2X1  _14447_
timestamp 0
transform 1 0 8690 0 1 9370
box -6 -8 86 248
use OAI21X1  _14448_
timestamp 0
transform 1 0 8530 0 1 9370
box -6 -8 106 248
use INVX1  _14449_
timestamp 0
transform 1 0 8050 0 1 9850
box -6 -8 66 248
use NAND2X1  _14450_
timestamp 0
transform 1 0 9090 0 -1 9850
box -6 -8 86 248
use OAI21X1  _14451_
timestamp 0
transform 1 0 8950 0 -1 9850
box -6 -8 106 248
use NAND2X1  _14452_
timestamp 0
transform 1 0 8910 0 1 10330
box -6 -8 86 248
use NAND2X1  _14453_
timestamp 0
transform 1 0 8310 0 1 9850
box -6 -8 86 248
use OAI21X1  _14454_
timestamp 0
transform 1 0 8170 0 1 9850
box -6 -8 106 248
use NAND2X1  _14455_
timestamp 0
transform 1 0 8610 0 1 8890
box -6 -8 86 248
use OAI21X1  _14456_
timestamp 0
transform 1 0 8590 0 -1 9370
box -6 -8 106 248
use INVX1  _14457_
timestamp 0
transform 1 0 8270 0 -1 10810
box -6 -8 66 248
use NAND3X1  _14458_
timestamp 0
transform 1 0 8370 0 -1 10330
box -6 -8 106 248
use NAND2X1  _14459_
timestamp 0
transform 1 0 8170 0 1 9370
box -6 -8 86 248
use OAI21X1  _14460_
timestamp 0
transform -1 0 8110 0 1 9370
box -6 -8 106 248
use NAND2X1  _14461_
timestamp 0
transform 1 0 8210 0 -1 9370
box -6 -8 86 248
use OAI21X1  _14462_
timestamp 0
transform 1 0 8050 0 -1 9370
box -6 -8 106 248
use NAND2X1  _14463_
timestamp 0
transform 1 0 8250 0 -1 10330
box -6 -8 86 248
use OAI21X1  _14464_
timestamp 0
transform -1 0 8050 0 -1 10330
box -6 -8 106 248
use OAI21X1  _14465_
timestamp 0
transform -1 0 8190 0 -1 10330
box -6 -8 106 248
use OAI21X1  _14466_
timestamp 0
transform -1 0 7850 0 1 9850
box -6 -8 106 248
use OAI21X1  _14467_
timestamp 0
transform -1 0 7990 0 1 9850
box -6 -8 106 248
use NAND2X1  _14468_
timestamp 0
transform 1 0 7930 0 1 10330
box -6 -8 86 248
use OAI21X1  _14469_
timestamp 0
transform 1 0 7770 0 1 10330
box -6 -8 106 248
use NAND2X1  _14470_
timestamp 0
transform -1 0 7450 0 1 9850
box -6 -8 86 248
use OAI21X1  _14471_
timestamp 0
transform 1 0 7190 0 1 9370
box -6 -8 106 248
use NAND2X1  _14472_
timestamp 0
transform 1 0 9370 0 -1 9850
box -6 -8 86 248
use OAI21X1  _14473_
timestamp 0
transform 1 0 9230 0 -1 9850
box -6 -8 106 248
use NAND2X1  _14474_
timestamp 0
transform 1 0 7790 0 1 10810
box -6 -8 86 248
use OAI21X1  _14475_
timestamp 0
transform -1 0 8130 0 1 10810
box -6 -8 106 248
use INVX1  _14476_
timestamp 0
transform 1 0 9490 0 -1 9850
box -6 -8 66 248
use NAND2X1  _14477_
timestamp 0
transform -1 0 9210 0 1 9370
box -6 -8 86 248
use OAI21X1  _14478_
timestamp 0
transform -1 0 9370 0 1 9370
box -6 -8 106 248
use INVX1  _14479_
timestamp 0
transform -1 0 7850 0 -1 10810
box -6 -8 66 248
use NAND2X1  _14480_
timestamp 0
transform 1 0 9750 0 -1 9850
box -6 -8 86 248
use OAI21X1  _14481_
timestamp 0
transform 1 0 9590 0 -1 9850
box -6 -8 106 248
use NAND2X1  _14482_
timestamp 0
transform 1 0 9990 0 -1 9370
box -6 -8 86 248
use OAI21X1  _14483_
timestamp 0
transform 1 0 9850 0 -1 9370
box -6 -8 106 248
use NAND2X1  _14484_
timestamp 0
transform 1 0 9930 0 -1 10330
box -6 -8 86 248
use OAI21X1  _14485_
timestamp 0
transform 1 0 9550 0 -1 10330
box -6 -8 106 248
use NAND2X1  _14486_
timestamp 0
transform 1 0 9870 0 -1 9850
box -6 -8 86 248
use OAI21X1  _14487_
timestamp 0
transform 1 0 9910 0 1 9370
box -6 -8 106 248
use NAND2X1  _14488_
timestamp 0
transform -1 0 9610 0 1 9850
box -6 -8 86 248
use OAI21X1  _14489_
timestamp 0
transform 1 0 9390 0 1 9850
box -6 -8 106 248
use OAI21X1  _14490_
timestamp 0
transform 1 0 8430 0 -1 9850
box -6 -8 106 248
use OAI21X1  _14491_
timestamp 0
transform -1 0 8670 0 -1 9850
box -6 -8 106 248
use OAI21X1  _14492_
timestamp 0
transform 1 0 8270 0 -1 9850
box -6 -8 106 248
use OAI21X1  _14493_
timestamp 0
transform 1 0 8110 0 -1 9850
box -6 -8 106 248
use NAND2X1  _14494_
timestamp 0
transform -1 0 7590 0 1 9370
box -6 -8 86 248
use OAI21X1  _14495_
timestamp 0
transform -1 0 7730 0 1 9370
box -6 -8 106 248
use NAND2X1  _14496_
timestamp 0
transform 1 0 7430 0 -1 10810
box -6 -8 86 248
use OAI21X1  _14497_
timestamp 0
transform -1 0 7450 0 1 9370
box -6 -8 106 248
use NAND2X1  _14498_
timestamp 0
transform 1 0 9570 0 -1 9370
box -6 -8 86 248
use OAI21X1  _14499_
timestamp 0
transform -1 0 9690 0 1 8890
box -6 -8 106 248
use DFFPOSX1  _14500_
timestamp 0
transform 1 0 7290 0 -1 7450
box -6 -8 246 248
use DFFPOSX1  _14501_
timestamp 0
transform -1 0 8010 0 1 7930
box -6 -8 246 248
use DFFPOSX1  _14502_
timestamp 0
transform 1 0 6650 0 -1 7450
box -6 -8 246 248
use DFFPOSX1  _14503_
timestamp 0
transform 1 0 7010 0 1 7450
box -6 -8 246 248
use DFFPOSX1  _14504_
timestamp 0
transform -1 0 8290 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _14505_
timestamp 0
transform 1 0 7950 0 -1 7450
box -6 -8 246 248
use DFFPOSX1  _14506_
timestamp 0
transform -1 0 9450 0 1 6970
box -6 -8 246 248
use DFFPOSX1  _14507_
timestamp 0
transform 1 0 7610 0 1 6490
box -6 -8 246 248
use DFFPOSX1  _14508_
timestamp 0
transform -1 0 8650 0 -1 7450
box -6 -8 246 248
use DFFPOSX1  _14509_
timestamp 0
transform -1 0 8410 0 -1 7930
box -6 -8 246 248
use DFFPOSX1  _14510_
timestamp 0
transform 1 0 8650 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _14511_
timestamp 0
transform 1 0 9590 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _14512_
timestamp 0
transform 1 0 7210 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _14513_
timestamp 0
transform -1 0 7830 0 1 8410
box -6 -8 246 248
use DFFPOSX1  _14514_
timestamp 0
transform -1 0 7670 0 1 6970
box -6 -8 246 248
use DFFPOSX1  _14515_
timestamp 0
transform 1 0 6570 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _14516_
timestamp 0
transform -1 0 8850 0 -1 6490
box -6 -8 246 248
use DFFPOSX1  _14517_
timestamp 0
transform -1 0 10510 0 1 7450
box -6 -8 246 248
use DFFPOSX1  _14518_
timestamp 0
transform -1 0 9230 0 -1 6490
box -6 -8 246 248
use DFFPOSX1  _14519_
timestamp 0
transform -1 0 9230 0 -1 6970
box -6 -8 246 248
use DFFPOSX1  _14520_
timestamp 0
transform -1 0 9290 0 -1 7450
box -6 -8 246 248
use DFFPOSX1  _14521_
timestamp 0
transform -1 0 8670 0 1 7450
box -6 -8 246 248
use DFFPOSX1  _14522_
timestamp 0
transform 1 0 9290 0 -1 7450
box -6 -8 246 248
use DFFPOSX1  _14523_
timestamp 0
transform 1 0 9530 0 1 7450
box -6 -8 246 248
use DFFPOSX1  _14524_
timestamp 0
transform 1 0 8630 0 1 9850
box -6 -8 246 248
use DFFPOSX1  _14525_
timestamp 0
transform 1 0 8570 0 -1 11290
box -6 -8 246 248
use DFFPOSX1  _14526_
timestamp 0
transform 1 0 8250 0 1 9370
box -6 -8 246 248
use DFFPOSX1  _14527_
timestamp 0
transform -1 0 8910 0 -1 9850
box -6 -8 246 248
use DFFPOSX1  _14528_
timestamp 0
transform 1 0 8390 0 1 9850
box -6 -8 246 248
use DFFPOSX1  _14529_
timestamp 0
transform -1 0 8530 0 -1 9370
box -6 -8 246 248
use DFFPOSX1  _14530_
timestamp 0
transform 1 0 7730 0 1 9370
box -6 -8 246 248
use DFFPOSX1  _14531_
timestamp 0
transform 1 0 7770 0 -1 9370
box -6 -8 246 248
use DFFPOSX1  _14532_
timestamp 0
transform 1 0 7670 0 -1 10330
box -6 -8 246 248
use DFFPOSX1  _14533_
timestamp 0
transform -1 0 7830 0 -1 9850
box -6 -8 246 248
use DFFPOSX1  _14534_
timestamp 0
transform -1 0 7730 0 1 10330
box -6 -8 246 248
use DFFPOSX1  _14535_
timestamp 0
transform -1 0 7130 0 1 9370
box -6 -8 246 248
use DFFPOSX1  _14536_
timestamp 0
transform -1 0 9110 0 1 9850
box -6 -8 246 248
use DFFPOSX1  _14537_
timestamp 0
transform 1 0 8590 0 -1 10810
box -6 -8 246 248
use DFFPOSX1  _14538_
timestamp 0
transform 1 0 9370 0 1 9370
box -6 -8 246 248
use DFFPOSX1  _14539_
timestamp 0
transform 1 0 9110 0 1 9850
box -6 -8 246 248
use DFFPOSX1  _14540_
timestamp 0
transform 1 0 9690 0 1 8890
box -6 -8 246 248
use DFFPOSX1  _14541_
timestamp 0
transform 1 0 9650 0 -1 10330
box -6 -8 246 248
use DFFPOSX1  _14542_
timestamp 0
transform -1 0 9850 0 1 9370
box -6 -8 246 248
use DFFPOSX1  _14543_
timestamp 0
transform -1 0 10570 0 -1 9850
box -6 -8 246 248
use DFFPOSX1  _14544_
timestamp 0
transform 1 0 7450 0 1 9850
box -6 -8 246 248
use DFFPOSX1  _14545_
timestamp 0
transform 1 0 7830 0 -1 9850
box -6 -8 246 248
use DFFPOSX1  _14546_
timestamp 0
transform 1 0 7530 0 -1 9370
box -6 -8 246 248
use DFFPOSX1  _14547_
timestamp 0
transform 1 0 7290 0 -1 9370
box -6 -8 246 248
use DFFPOSX1  _14548_
timestamp 0
transform 1 0 7150 0 -1 10810
box -6 -8 246 248
use DFFPOSX1  _14549_
timestamp 0
transform 1 0 7510 0 -1 10810
box -6 -8 246 248
use DFFPOSX1  _14550_
timestamp 0
transform 1 0 8130 0 1 10330
box -6 -8 246 248
use DFFPOSX1  _14551_
timestamp 0
transform 1 0 8490 0 1 10330
box -6 -8 246 248
use DFFPOSX1  _14552_
timestamp 0
transform 1 0 7510 0 1 10810
box -6 -8 246 248
use DFFPOSX1  _14553_
timestamp 0
transform 1 0 7850 0 -1 10810
box -6 -8 246 248
use DFFPOSX1  _14554_
timestamp 0
transform 1 0 8630 0 -1 10330
box -6 -8 246 248
use DFFPOSX1  _14555_
timestamp 0
transform -1 0 8950 0 -1 8890
box -6 -8 246 248
use INVX1  _14556_
timestamp 0
transform -1 0 14810 0 -1 2170
box -6 -8 66 248
use INVX1  _14557_
timestamp 0
transform -1 0 14550 0 -1 2170
box -6 -8 66 248
use INVX1  _14558_
timestamp 0
transform -1 0 14130 0 1 1690
box -6 -8 66 248
use INVX1  _14559_
timestamp 0
transform -1 0 12990 0 -1 1690
box -6 -8 66 248
use INVX1  _14560_
timestamp 0
transform -1 0 12230 0 1 1210
box -6 -8 66 248
use INVX1  _14561_
timestamp 0
transform -1 0 13130 0 1 1690
box -6 -8 66 248
use NAND2X1  _14562_
timestamp 0
transform 1 0 11750 0 1 1210
box -6 -8 86 248
use OAI21X1  _14563_
timestamp 0
transform -1 0 12110 0 1 1210
box -6 -8 106 248
use NAND2X1  _14564_
timestamp 0
transform -1 0 12610 0 -1 1690
box -6 -8 86 248
use OAI21X1  _14565_
timestamp 0
transform -1 0 12770 0 -1 1690
box -6 -8 106 248
use NAND2X1  _14566_
timestamp 0
transform -1 0 14650 0 1 1690
box -6 -8 86 248
use OAI21X1  _14567_
timestamp 0
transform -1 0 14710 0 -1 2170
box -6 -8 106 248
use INVX1  _14568_
timestamp 0
transform -1 0 15530 0 -1 2170
box -6 -8 66 248
use NAND2X1  _14569_
timestamp 0
transform 1 0 15090 0 -1 2170
box -6 -8 86 248
use OAI21X1  _14570_
timestamp 0
transform 1 0 15090 0 1 2170
box -6 -8 106 248
use NAND2X1  _14571_
timestamp 0
transform 1 0 14090 0 -1 2170
box -6 -8 86 248
use OAI21X1  _14572_
timestamp 0
transform -1 0 14250 0 1 2170
box -6 -8 106 248
use INVX1  _14573_
timestamp 0
transform -1 0 12570 0 1 1210
box -6 -8 66 248
use INVX1  _14574_
timestamp 0
transform 1 0 11690 0 1 730
box -6 -8 66 248
use OAI21X1  _14575_
timestamp 0
transform 1 0 11870 0 1 1210
box -6 -8 106 248
use INVX1  _14576_
timestamp 0
transform -1 0 13390 0 -1 1690
box -6 -8 66 248
use AOI21X1  _14577_
timestamp 0
transform -1 0 13290 0 -1 1690
box -6 -8 106 248
use OAI21X1  _14578_
timestamp 0
transform 1 0 13030 0 -1 1690
box -6 -8 106 248
use OAI21X1  _14579_
timestamp 0
transform -1 0 13530 0 1 1690
box -6 -8 106 248
use INVX1  _14580_
timestamp 0
transform -1 0 13050 0 1 1210
box -6 -8 66 248
use NAND2X1  _14581_
timestamp 0
transform 1 0 14370 0 -1 2170
box -6 -8 86 248
use OAI21X1  _14582_
timestamp 0
transform -1 0 14310 0 -1 2170
box -6 -8 106 248
use NAND2X1  _14583_
timestamp 0
transform -1 0 13890 0 -1 2170
box -6 -8 86 248
use OAI21X1  _14584_
timestamp 0
transform -1 0 14050 0 -1 2170
box -6 -8 106 248
use INVX1  _14585_
timestamp 0
transform -1 0 12430 0 1 1690
box -6 -8 66 248
use NAND2X1  _14586_
timestamp 0
transform -1 0 9850 0 -1 730
box -6 -8 86 248
use INVX1  _14587_
timestamp 0
transform -1 0 10070 0 -1 730
box -6 -8 66 248
use INVX1  _14588_
timestamp 0
transform 1 0 10050 0 1 250
box -6 -8 66 248
use NAND2X1  _14589_
timestamp 0
transform -1 0 10010 0 1 250
box -6 -8 86 248
use NAND2X1  _14590_
timestamp 0
transform 1 0 9890 0 -1 730
box -6 -8 86 248
use NAND2X1  _14591_
timestamp 0
transform -1 0 12090 0 1 1690
box -6 -8 86 248
use OAI21X1  _14592_
timestamp 0
transform 1 0 11990 0 -1 1690
box -6 -8 106 248
use INVX8  _14593_
timestamp 0
transform 1 0 13070 0 1 730
box -6 -8 126 248
use INVX2  _14594_
timestamp 0
transform -1 0 14010 0 1 1690
box -6 -8 66 248
use NOR2X1  _14595_
timestamp 0
transform 1 0 11310 0 -1 1210
box -6 -8 86 248
use AND2X2  _14596_
timestamp 0
transform 1 0 14310 0 1 2170
box -6 -8 106 248
use AND2X2  _14597_
timestamp 0
transform -1 0 15030 0 1 2170
box -6 -8 106 248
use NOR2X1  _14598_
timestamp 0
transform 1 0 13830 0 1 1690
box -6 -8 86 248
use NOR2X1  _14599_
timestamp 0
transform -1 0 12890 0 -1 1690
box -6 -8 86 248
use NAND2X1  _14600_
timestamp 0
transform -1 0 13030 0 1 1690
box -6 -8 86 248
use NOR2X1  _14601_
timestamp 0
transform -1 0 11950 0 -1 1690
box -6 -8 86 248
use INVX1  _14602_
timestamp 0
transform 1 0 14930 0 1 1690
box -6 -8 66 248
use NAND2X1  _14603_
timestamp 0
transform 1 0 15350 0 1 1690
box -6 -8 86 248
use OAI21X1  _14604_
timestamp 0
transform 1 0 15190 0 1 1690
box -6 -8 106 248
use AOI21X1  _14605_
timestamp 0
transform -1 0 15150 0 1 1690
box -6 -8 106 248
use NAND2X1  _14606_
timestamp 0
transform -1 0 14650 0 -1 1690
box -6 -8 86 248
use NAND2X1  _14607_
timestamp 0
transform -1 0 15050 0 -1 1690
box -6 -8 86 248
use INVX1  _14608_
timestamp 0
transform -1 0 14930 0 -1 1690
box -6 -8 66 248
use NOR2X1  _14609_
timestamp 0
transform 1 0 15090 0 -1 1690
box -6 -8 86 248
use OAI21X1  _14610_
timestamp 0
transform -1 0 15890 0 1 1690
box -6 -8 106 248
use OR2X2  _14611_
timestamp 0
transform 1 0 16050 0 1 1690
box -6 -8 106 248
use NOR2X1  _14612_
timestamp 0
transform 1 0 16210 0 1 1690
box -6 -8 86 248
use INVX1  _14613_
timestamp 0
transform 1 0 16330 0 1 1690
box -6 -8 66 248
use NAND2X1  _14614_
timestamp 0
transform 1 0 15930 0 1 1690
box -6 -8 86 248
use OAI21X1  _14615_
timestamp 0
transform 1 0 15230 0 -1 1690
box -6 -8 106 248
use AOI21X1  _14616_
timestamp 0
transform -1 0 15730 0 1 1690
box -6 -8 106 248
use OAI21X1  _14617_
timestamp 0
transform -1 0 14810 0 -1 1690
box -6 -8 106 248
use AND2X2  _14618_
timestamp 0
transform 1 0 13750 0 -1 1210
box -6 -8 106 248
use NOR2X1  _14619_
timestamp 0
transform -1 0 13710 0 -1 1210
box -6 -8 86 248
use NOR2X1  _14620_
timestamp 0
transform 1 0 14370 0 1 1210
box -6 -8 86 248
use AND2X2  _14621_
timestamp 0
transform -1 0 14310 0 1 1210
box -6 -8 106 248
use NOR2X1  _14622_
timestamp 0
transform 1 0 13950 0 1 1210
box -6 -8 86 248
use OAI21X1  _14623_
timestamp 0
transform -1 0 14170 0 1 1210
box -6 -8 106 248
use NAND2X1  _14624_
timestamp 0
transform -1 0 13890 0 1 1210
box -6 -8 86 248
use AOI21X1  _14625_
timestamp 0
transform -1 0 14050 0 -1 1690
box -6 -8 106 248
use OAI21X1  _14626_
timestamp 0
transform 1 0 13890 0 1 730
box -6 -8 106 248
use AND2X2  _14627_
timestamp 0
transform 1 0 14710 0 -1 1210
box -6 -8 106 248
use NOR2X1  _14628_
timestamp 0
transform -1 0 14650 0 -1 1210
box -6 -8 86 248
use NOR2X1  _14629_
timestamp 0
transform 1 0 14450 0 -1 1210
box -6 -8 86 248
use OAI21X1  _14630_
timestamp 0
transform 1 0 14010 0 -1 1210
box -6 -8 106 248
use NOR2X1  _14631_
timestamp 0
transform -1 0 14250 0 -1 1210
box -6 -8 86 248
use OAI21X1  _14632_
timestamp 0
transform -1 0 14390 0 -1 1210
box -6 -8 106 248
use NAND2X1  _14633_
timestamp 0
transform -1 0 13970 0 -1 1210
box -6 -8 86 248
use AOI21X1  _14634_
timestamp 0
transform -1 0 13850 0 1 730
box -6 -8 106 248
use NAND3X1  _14635_
timestamp 0
transform 1 0 14490 0 1 1210
box -6 -8 106 248
use INVX1  _14636_
timestamp 0
transform 1 0 14650 0 1 1210
box -6 -8 66 248
use AOI21X1  _14637_
timestamp 0
transform 1 0 14750 0 1 1210
box -6 -8 106 248
use AND2X2  _14638_
timestamp 0
transform 1 0 15010 0 1 1210
box -6 -8 106 248
use AND2X2  _14639_
timestamp 0
transform 1 0 15550 0 1 1210
box -6 -8 106 248
use NOR2X1  _14640_
timestamp 0
transform -1 0 15490 0 1 1210
box -6 -8 86 248
use OAI21X1  _14641_
timestamp 0
transform -1 0 15810 0 1 1210
box -6 -8 106 248
use NAND2X1  _14642_
timestamp 0
transform -1 0 14970 0 1 1210
box -6 -8 86 248
use NOR2X1  _14643_
timestamp 0
transform 1 0 15870 0 1 1210
box -6 -8 86 248
use NAND2X1  _14644_
timestamp 0
transform 1 0 16030 0 -1 1690
box -6 -8 86 248
use NAND2X1  _14645_
timestamp 0
transform -1 0 15990 0 -1 1690
box -6 -8 86 248
use OAI21X1  _14646_
timestamp 0
transform -1 0 15730 0 -1 1690
box -6 -8 106 248
use AOI21X1  _14647_
timestamp 0
transform 1 0 15770 0 -1 1690
box -6 -8 106 248
use AOI21X1  _14648_
timestamp 0
transform 1 0 16170 0 -1 1690
box -6 -8 106 248
use AND2X2  _14649_
timestamp 0
transform -1 0 17150 0 1 1690
box -6 -8 106 248
use NOR2X1  _14650_
timestamp 0
transform 1 0 16890 0 1 16570
box -6 -8 86 248
use NOR2X1  _14651_
timestamp 0
transform 1 0 16990 0 -1 1690
box -6 -8 86 248
use NAND2X1  _14652_
timestamp 0
transform -1 0 16650 0 -1 1690
box -6 -8 86 248
use NOR2X1  _14653_
timestamp 0
transform 1 0 16450 0 -1 1690
box -6 -8 86 248
use NOR2X1  _14654_
timestamp 0
transform 1 0 16310 0 -1 1690
box -6 -8 86 248
use OAI21X1  _14655_
timestamp 0
transform -1 0 16930 0 -1 1690
box -6 -8 106 248
use AOI21X1  _14656_
timestamp 0
transform 1 0 16670 0 1 1690
box -6 -8 106 248
use INVX1  _14657_
timestamp 0
transform 1 0 16410 0 1 1210
box -6 -8 66 248
use INVX1  _14658_
timestamp 0
transform 1 0 16710 0 -1 1690
box -6 -8 66 248
use OAI21X1  _14659_
timestamp 0
transform -1 0 16610 0 1 1210
box -6 -8 106 248
use AND2X2  _14660_
timestamp 0
transform 1 0 16130 0 1 1210
box -6 -8 106 248
use AOI21X1  _14661_
timestamp 0
transform 1 0 16270 0 1 1210
box -6 -8 106 248
use NAND2X1  _14662_
timestamp 0
transform -1 0 16990 0 1 730
box -6 -8 86 248
use OR2X2  _14663_
timestamp 0
transform 1 0 17030 0 1 730
box -6 -8 106 248
use NAND2X1  _14664_
timestamp 0
transform 1 0 16670 0 1 730
box -6 -8 86 248
use OR2X2  _14665_
timestamp 0
transform 1 0 17070 0 -1 1210
box -6 -8 106 248
use INVX1  _14666_
timestamp 0
transform 1 0 16790 0 1 730
box -6 -8 66 248
use INVX1  _14667_
timestamp 0
transform 1 0 17050 0 -1 730
box -6 -8 66 248
use OAI21X1  _14668_
timestamp 0
transform 1 0 16890 0 -1 730
box -6 -8 106 248
use NAND2X1  _14669_
timestamp 0
transform 1 0 16930 0 -1 1210
box -6 -8 86 248
use OAI21X1  _14670_
timestamp 0
transform -1 0 16750 0 -1 1210
box -6 -8 106 248
use AOI21X1  _14671_
timestamp 0
transform -1 0 16890 0 -1 1210
box -6 -8 106 248
use OAI21X1  _14672_
timestamp 0
transform -1 0 16850 0 -1 730
box -6 -8 106 248
use NAND2X1  _14673_
timestamp 0
transform -1 0 16170 0 -1 250
box -6 -8 86 248
use OR2X2  _14674_
timestamp 0
transform -1 0 16470 0 1 250
box -6 -8 106 248
use NAND2X1  _14675_
timestamp 0
transform 1 0 16230 0 1 250
box -6 -8 86 248
use OR2X2  _14676_
timestamp 0
transform 1 0 16130 0 -1 730
box -6 -8 106 248
use AOI21X1  _14677_
timestamp 0
transform -1 0 16090 0 -1 730
box -6 -8 106 248
use OAI21X1  _14678_
timestamp 0
transform 1 0 16290 0 1 730
box -6 -8 106 248
use AOI21X1  _14679_
timestamp 0
transform 1 0 16290 0 -1 730
box -6 -8 106 248
use NAND2X1  _14680_
timestamp 0
transform -1 0 16070 0 1 1210
box -6 -8 86 248
use AND2X2  _14681_
timestamp 0
transform 1 0 16510 0 1 250
box -6 -8 106 248
use NOR2X1  _14682_
timestamp 0
transform -1 0 16050 0 -1 250
box -6 -8 86 248
use NOR2X1  _14683_
timestamp 0
transform 1 0 16650 0 1 250
box -6 -8 86 248
use NAND3X1  _14684_
timestamp 0
transform -1 0 16690 0 -1 730
box -6 -8 106 248
use NOR2X1  _14685_
timestamp 0
transform 1 0 15970 0 -1 1210
box -6 -8 86 248
use INVX1  _14686_
timestamp 0
transform -1 0 16870 0 1 1210
box -6 -8 66 248
use AOI21X1  _14687_
timestamp 0
transform -1 0 16750 0 1 1210
box -6 -8 106 248
use OAI21X1  _14688_
timestamp 0
transform -1 0 16530 0 -1 730
box -6 -8 106 248
use INVX1  _14689_
timestamp 0
transform 1 0 16390 0 -1 1210
box -6 -8 66 248
use OAI21X1  _14690_
timestamp 0
transform -1 0 16590 0 -1 1210
box -6 -8 106 248
use AOI21X1  _14691_
timestamp 0
transform -1 0 15930 0 -1 1210
box -6 -8 106 248
use NAND2X1  _14692_
timestamp 0
transform -1 0 14430 0 -1 730
box -6 -8 86 248
use OR2X2  _14693_
timestamp 0
transform 1 0 14490 0 -1 730
box -6 -8 106 248
use NAND2X1  _14694_
timestamp 0
transform -1 0 14850 0 -1 730
box -6 -8 86 248
use OR2X2  _14695_
timestamp 0
transform -1 0 15050 0 1 730
box -6 -8 106 248
use NAND2X1  _14696_
timestamp 0
transform 1 0 14710 0 1 730
box -6 -8 86 248
use NAND2X1  _14697_
timestamp 0
transform 1 0 14830 0 1 730
box -6 -8 86 248
use OAI21X1  _14698_
timestamp 0
transform -1 0 14970 0 -1 1210
box -6 -8 106 248
use AOI21X1  _14699_
timestamp 0
transform 1 0 15010 0 -1 1210
box -6 -8 106 248
use OAI21X1  _14700_
timestamp 0
transform -1 0 14730 0 -1 730
box -6 -8 106 248
use NAND2X1  _14701_
timestamp 0
transform 1 0 14870 0 1 250
box -6 -8 86 248
use INVX1  _14702_
timestamp 0
transform -1 0 14610 0 -1 250
box -6 -8 66 248
use INVX1  _14703_
timestamp 0
transform -1 0 14390 0 -1 250
box -6 -8 66 248
use NAND2X1  _14704_
timestamp 0
transform -1 0 14510 0 -1 250
box -6 -8 86 248
use NAND2X1  _14705_
timestamp 0
transform 1 0 15010 0 1 250
box -6 -8 86 248
use NAND2X1  _14706_
timestamp 0
transform 1 0 14230 0 -1 730
box -6 -8 86 248
use NOR2X1  _14707_
timestamp 0
transform -1 0 14190 0 -1 730
box -6 -8 86 248
use NOR2X1  _14708_
timestamp 0
transform -1 0 14070 0 -1 730
box -6 -8 86 248
use OAI21X1  _14709_
timestamp 0
transform 1 0 14030 0 1 730
box -6 -8 106 248
use AOI21X1  _14710_
timestamp 0
transform 1 0 14190 0 1 730
box -6 -8 106 248
use NOR2X1  _14711_
timestamp 0
transform -1 0 14730 0 -1 250
box -6 -8 86 248
use OAI21X1  _14712_
timestamp 0
transform 1 0 15130 0 1 250
box -6 -8 106 248
use INVX1  _14713_
timestamp 0
transform 1 0 15290 0 1 250
box -6 -8 66 248
use OR2X2  _14714_
timestamp 0
transform 1 0 15010 0 -1 730
box -6 -8 106 248
use OAI21X1  _14715_
timestamp 0
transform 1 0 15170 0 -1 730
box -6 -8 106 248
use AND2X2  _14716_
timestamp 0
transform -1 0 15650 0 1 250
box -6 -8 106 248
use NOR2X1  _14717_
timestamp 0
transform 1 0 15710 0 1 250
box -6 -8 86 248
use NOR2X1  _14718_
timestamp 0
transform -1 0 15630 0 -1 250
box -6 -8 86 248
use NAND2X1  _14719_
timestamp 0
transform -1 0 15390 0 -1 730
box -6 -8 86 248
use OR2X2  _14720_
timestamp 0
transform 1 0 15570 0 -1 730
box -6 -8 106 248
use NAND2X1  _14721_
timestamp 0
transform 1 0 15430 0 -1 730
box -6 -8 86 248
use OAI21X1  _14722_
timestamp 0
transform 1 0 15490 0 1 730
box -6 -8 106 248
use AOI21X1  _14723_
timestamp 0
transform -1 0 15430 0 1 730
box -6 -8 106 248
use NAND2X1  _14724_
timestamp 0
transform -1 0 15930 0 1 250
box -6 -8 86 248
use NAND2X1  _14725_
timestamp 0
transform -1 0 15790 0 -1 730
box -6 -8 86 248
use AND2X2  _14726_
timestamp 0
transform -1 0 15770 0 -1 250
box -6 -8 106 248
use NOR2X1  _14727_
timestamp 0
transform 1 0 15830 0 -1 250
box -6 -8 86 248
use NOR2X1  _14728_
timestamp 0
transform 1 0 15430 0 -1 250
box -6 -8 86 248
use INVX1  _14729_
timestamp 0
transform 1 0 16130 0 1 250
box -6 -8 66 248
use OR2X2  _14730_
timestamp 0
transform 1 0 15970 0 1 250
box -6 -8 106 248
use AOI21X1  _14731_
timestamp 0
transform 1 0 15830 0 -1 730
box -6 -8 106 248
use OAI21X1  _14732_
timestamp 0
transform 1 0 16030 0 1 730
box -6 -8 106 248
use AOI21X1  _14733_
timestamp 0
transform -1 0 15970 0 1 730
box -6 -8 106 248
use NAND2X1  _14734_
timestamp 0
transform 1 0 12790 0 -1 1210
box -6 -8 86 248
use NOR2X1  _14735_
timestamp 0
transform 1 0 14890 0 -1 730
box -6 -8 86 248
use NAND3X1  _14736_
timestamp 0
transform -1 0 15510 0 1 250
box -6 -8 106 248
use NAND3X1  _14737_
timestamp 0
transform -1 0 15130 0 -1 250
box -6 -8 106 248
use INVX1  _14738_
timestamp 0
transform -1 0 15390 0 -1 250
box -6 -8 66 248
use AOI21X1  _14739_
timestamp 0
transform -1 0 15290 0 -1 250
box -6 -8 106 248
use AND2X2  _14740_
timestamp 0
transform -1 0 14870 0 -1 250
box -6 -8 106 248
use OAI21X1  _14741_
timestamp 0
transform 1 0 14710 0 1 250
box -6 -8 106 248
use NAND2X1  _14742_
timestamp 0
transform 1 0 12190 0 -1 250
box -6 -8 86 248
use OR2X2  _14743_
timestamp 0
transform -1 0 12150 0 -1 250
box -6 -8 106 248
use NAND2X1  _14744_
timestamp 0
transform 1 0 11910 0 -1 250
box -6 -8 86 248
use NOR2X1  _14745_
timestamp 0
transform -1 0 12530 0 1 250
box -6 -8 86 248
use AND2X2  _14746_
timestamp 0
transform -1 0 12690 0 1 250
box -6 -8 106 248
use OAI21X1  _14747_
timestamp 0
transform -1 0 12510 0 -1 730
box -6 -8 106 248
use AOI21X1  _14748_
timestamp 0
transform -1 0 12730 0 -1 1210
box -6 -8 106 248
use INVX1  _14749_
timestamp 0
transform -1 0 11730 0 -1 250
box -6 -8 66 248
use OAI21X1  _14750_
timestamp 0
transform -1 0 11870 0 -1 250
box -6 -8 106 248
use NAND2X1  _14751_
timestamp 0
transform -1 0 11350 0 -1 250
box -6 -8 86 248
use OR2X2  _14752_
timestamp 0
transform 1 0 12170 0 1 250
box -6 -8 106 248
use NAND2X1  _14753_
timestamp 0
transform 1 0 12330 0 1 250
box -6 -8 86 248
use OR2X2  _14754_
timestamp 0
transform -1 0 12210 0 -1 730
box -6 -8 106 248
use AOI21X1  _14755_
timestamp 0
transform 1 0 12270 0 -1 730
box -6 -8 106 248
use OAI21X1  _14756_
timestamp 0
transform -1 0 11930 0 -1 730
box -6 -8 106 248
use AOI21X1  _14757_
timestamp 0
transform -1 0 12070 0 -1 730
box -6 -8 106 248
use NOR2X1  _14758_
timestamp 0
transform 1 0 12750 0 1 250
box -6 -8 86 248
use NOR2X1  _14759_
timestamp 0
transform -1 0 11470 0 -1 250
box -6 -8 86 248
use OAI21X1  _14760_
timestamp 0
transform -1 0 11630 0 -1 250
box -6 -8 106 248
use AOI21X1  _14761_
timestamp 0
transform 1 0 12730 0 -1 250
box -6 -8 106 248
use AND2X2  _14762_
timestamp 0
transform 1 0 12450 0 -1 250
box -6 -8 106 248
use NOR2X1  _14763_
timestamp 0
transform -1 0 12410 0 -1 250
box -6 -8 86 248
use OR2X2  _14764_
timestamp 0
transform 1 0 12590 0 -1 250
box -6 -8 106 248
use OR2X2  _14765_
timestamp 0
transform 1 0 13450 0 1 250
box -6 -8 106 248
use OAI21X1  _14766_
timestamp 0
transform 1 0 12870 0 -1 250
box -6 -8 106 248
use NAND2X1  _14767_
timestamp 0
transform 1 0 13030 0 1 250
box -6 -8 86 248
use OAI21X1  _14768_
timestamp 0
transform 1 0 12790 0 1 730
box -6 -8 106 248
use AOI21X1  _14769_
timestamp 0
transform -1 0 12890 0 -1 730
box -6 -8 106 248
use NAND2X1  _14770_
timestamp 0
transform 1 0 12890 0 1 250
box -6 -8 86 248
use NAND2X1  _14771_
timestamp 0
transform -1 0 13690 0 -1 730
box -6 -8 86 248
use INVX1  _14772_
timestamp 0
transform 1 0 13510 0 -1 730
box -6 -8 66 248
use NOR2X1  _14773_
timestamp 0
transform -1 0 13950 0 1 250
box -6 -8 86 248
use NOR2X1  _14774_
timestamp 0
transform -1 0 13830 0 1 250
box -6 -8 86 248
use NAND3X1  _14775_
timestamp 0
transform -1 0 13250 0 1 250
box -6 -8 106 248
use OAI21X1  _14776_
timestamp 0
transform -1 0 13390 0 1 250
box -6 -8 106 248
use INVX1  _14777_
timestamp 0
transform 1 0 14010 0 1 250
box -6 -8 66 248
use NAND2X1  _14778_
timestamp 0
transform -1 0 13450 0 -1 730
box -6 -8 86 248
use AOI21X1  _14779_
timestamp 0
transform -1 0 13330 0 -1 730
box -6 -8 106 248
use OAI21X1  _14780_
timestamp 0
transform -1 0 13030 0 -1 730
box -6 -8 106 248
use AOI21X1  _14781_
timestamp 0
transform -1 0 13170 0 -1 730
box -6 -8 106 248
use NOR2X1  _14782_
timestamp 0
transform 1 0 13030 0 -1 250
box -6 -8 86 248
use NAND3X1  _14783_
timestamp 0
transform 1 0 13290 0 -1 250
box -6 -8 106 248
use OR2X2  _14784_
timestamp 0
transform -1 0 14510 0 1 250
box -6 -8 106 248
use NAND2X1  _14785_
timestamp 0
transform 1 0 14910 0 -1 250
box -6 -8 86 248
use NOR2X1  _14786_
timestamp 0
transform 1 0 13610 0 1 250
box -6 -8 86 248
use AND2X2  _14787_
timestamp 0
transform 1 0 13590 0 -1 250
box -6 -8 106 248
use NAND3X1  _14788_
timestamp 0
transform 1 0 13150 0 -1 250
box -6 -8 106 248
use AOI21X1  _14789_
timestamp 0
transform 1 0 13450 0 -1 250
box -6 -8 106 248
use NAND2X1  _14790_
timestamp 0
transform -1 0 13810 0 -1 250
box -6 -8 86 248
use AOI21X1  _14791_
timestamp 0
transform 1 0 14010 0 -1 250
box -6 -8 106 248
use OAI21X1  _14792_
timestamp 0
transform -1 0 14210 0 1 250
box -6 -8 106 248
use AND2X2  _14793_
timestamp 0
transform -1 0 11070 0 -1 250
box -6 -8 106 248
use NOR2X1  _14794_
timestamp 0
transform 1 0 11130 0 -1 250
box -6 -8 86 248
use NOR2X1  _14795_
timestamp 0
transform 1 0 11510 0 1 250
box -6 -8 86 248
use NAND2X1  _14796_
timestamp 0
transform 1 0 11650 0 1 250
box -6 -8 86 248
use NOR2X1  _14797_
timestamp 0
transform 1 0 16170 0 1 730
box -6 -8 86 248
use NAND2X1  _14798_
timestamp 0
transform 1 0 16110 0 -1 1210
box -6 -8 86 248
use AOI21X1  _14799_
timestamp 0
transform 1 0 16230 0 -1 1210
box -6 -8 106 248
use OAI21X1  _14800_
timestamp 0
transform -1 0 15770 0 -1 1210
box -6 -8 106 248
use NOR2X1  _14801_
timestamp 0
transform 1 0 14570 0 1 250
box -6 -8 86 248
use AND2X2  _14802_
timestamp 0
transform 1 0 13850 0 -1 250
box -6 -8 106 248
use OAI21X1  _14803_
timestamp 0
transform -1 0 14270 0 -1 250
box -6 -8 106 248
use AOI21X1  _14804_
timestamp 0
transform -1 0 14350 0 1 250
box -6 -8 106 248
use OAI21X1  _14805_
timestamp 0
transform 1 0 11910 0 1 250
box -6 -8 106 248
use NAND2X1  _14806_
timestamp 0
transform -1 0 11850 0 1 250
box -6 -8 86 248
use OAI21X1  _14807_
timestamp 0
transform -1 0 11630 0 -1 730
box -6 -8 106 248
use AOI21X1  _14808_
timestamp 0
transform -1 0 11790 0 -1 730
box -6 -8 106 248
use AOI21X1  _14809_
timestamp 0
transform 1 0 11210 0 1 250
box -6 -8 106 248
use AND2X2  _14810_
timestamp 0
transform 1 0 10830 0 -1 250
box -6 -8 106 248
use NOR2X1  _14811_
timestamp 0
transform 1 0 10690 0 -1 250
box -6 -8 86 248
use NOR2X1  _14812_
timestamp 0
transform -1 0 10650 0 -1 250
box -6 -8 86 248
use OR2X2  _14813_
timestamp 0
transform 1 0 11370 0 1 250
box -6 -8 106 248
use AOI21X1  _14814_
timestamp 0
transform 1 0 11250 0 -1 730
box -6 -8 106 248
use OAI21X1  _14815_
timestamp 0
transform -1 0 11210 0 -1 730
box -6 -8 106 248
use AOI21X1  _14816_
timestamp 0
transform 1 0 11390 0 -1 730
box -6 -8 106 248
use NAND2X1  _14817_
timestamp 0
transform -1 0 11170 0 1 250
box -6 -8 86 248
use AOI21X1  _14818_
timestamp 0
transform -1 0 10530 0 -1 250
box -6 -8 106 248
use OAI21X1  _14819_
timestamp 0
transform -1 0 11030 0 1 250
box -6 -8 106 248
use INVX1  _14820_
timestamp 0
transform -1 0 10350 0 1 250
box -6 -8 66 248
use NOR2X1  _14821_
timestamp 0
transform 1 0 10150 0 1 250
box -6 -8 86 248
use NOR2X1  _14822_
timestamp 0
transform 1 0 10410 0 1 250
box -6 -8 86 248
use NOR2X1  _14823_
timestamp 0
transform -1 0 10010 0 -1 250
box -6 -8 86 248
use NAND2X1  _14824_
timestamp 0
transform 1 0 10810 0 1 250
box -6 -8 86 248
use INVX1  _14825_
timestamp 0
transform -1 0 10290 0 -1 250
box -6 -8 66 248
use INVX1  _14826_
timestamp 0
transform -1 0 10390 0 -1 250
box -6 -8 66 248
use AOI21X1  _14827_
timestamp 0
transform -1 0 10170 0 -1 250
box -6 -8 106 248
use OAI21X1  _14828_
timestamp 0
transform 1 0 9790 0 -1 250
box -6 -8 106 248
use NAND2X1  _14829_
timestamp 0
transform -1 0 10210 0 -1 730
box -6 -8 86 248
use OAI21X1  _14830_
timestamp 0
transform 1 0 10650 0 -1 730
box -6 -8 106 248
use AOI21X1  _14831_
timestamp 0
transform 1 0 10370 0 -1 730
box -6 -8 106 248
use INVX1  _14832_
timestamp 0
transform -1 0 10990 0 -1 1210
box -6 -8 66 248
use NAND2X1  _14833_
timestamp 0
transform 1 0 10670 0 -1 1210
box -6 -8 86 248
use INVX1  _14834_
timestamp 0
transform -1 0 9610 0 -1 250
box -6 -8 66 248
use OAI21X1  _14835_
timestamp 0
transform -1 0 9750 0 -1 250
box -6 -8 106 248
use NAND2X1  _14836_
timestamp 0
transform -1 0 9230 0 -1 250
box -6 -8 86 248
use OR2X2  _14837_
timestamp 0
transform 1 0 9270 0 -1 250
box -6 -8 106 248
use NAND2X1  _14838_
timestamp 0
transform -1 0 9490 0 -1 250
box -6 -8 86 248
use NAND2X1  _14839_
timestamp 0
transform 1 0 10550 0 1 250
box -6 -8 86 248
use AOI21X1  _14840_
timestamp 0
transform -1 0 10770 0 1 250
box -6 -8 106 248
use INVX1  _14841_
timestamp 0
transform 1 0 10270 0 -1 730
box -6 -8 66 248
use AOI21X1  _14842_
timestamp 0
transform 1 0 10510 0 -1 730
box -6 -8 106 248
use AOI22X1  _14843_
timestamp 0
transform -1 0 10670 0 1 730
box -6 -8 126 248
use NOR2X1  _14844_
timestamp 0
transform -1 0 12350 0 -1 1690
box -6 -8 86 248
use OAI21X1  _14845_
timestamp 0
transform -1 0 12430 0 -1 1210
box -6 -8 106 248
use NOR2X1  _14846_
timestamp 0
transform 1 0 12410 0 -1 1690
box -6 -8 86 248
use NOR2X1  _14847_
timestamp 0
transform -1 0 11750 0 -1 1210
box -6 -8 86 248
use OAI21X1  _14848_
timestamp 0
transform -1 0 13590 0 -1 1210
box -6 -8 106 248
use NOR2X1  _14849_
timestamp 0
transform 1 0 11790 0 -1 1210
box -6 -8 86 248
use OAI21X1  _14850_
timestamp 0
transform -1 0 15370 0 1 1210
box -6 -8 106 248
use AOI21X1  _14851_
timestamp 0
transform 1 0 15490 0 1 1690
box -6 -8 106 248
use OAI21X1  _14852_
timestamp 0
transform -1 0 13750 0 1 1210
box -6 -8 106 248
use AOI21X1  _14853_
timestamp 0
transform -1 0 13450 0 1 1210
box -6 -8 106 248
use OAI21X1  _14854_
timestamp 0
transform 1 0 12850 0 1 1210
box -6 -8 106 248
use AOI21X1  _14855_
timestamp 0
transform 1 0 14430 0 1 1690
box -6 -8 106 248
use OAI21X1  _14856_
timestamp 0
transform -1 0 12270 0 1 730
box -6 -8 106 248
use AOI21X1  _14857_
timestamp 0
transform 1 0 12470 0 -1 1210
box -6 -8 106 248
use OAI21X1  _14858_
timestamp 0
transform 1 0 13070 0 -1 1210
box -6 -8 106 248
use AOI21X1  _14859_
timestamp 0
transform 1 0 13810 0 -1 1690
box -6 -8 106 248
use OAI21X1  _14860_
timestamp 0
transform -1 0 13610 0 1 1210
box -6 -8 106 248
use AOI21X1  _14861_
timestamp 0
transform 1 0 13430 0 -1 1690
box -6 -8 106 248
use OAI21X1  _14862_
timestamp 0
transform 1 0 12030 0 1 730
box -6 -8 106 248
use AOI21X1  _14863_
timestamp 0
transform 1 0 12190 0 -1 1210
box -6 -8 106 248
use OAI21X1  _14864_
timestamp 0
transform 1 0 10790 0 -1 730
box -6 -8 106 248
use AOI21X1  _14865_
timestamp 0
transform -1 0 11050 0 -1 730
box -6 -8 106 248
use NOR2X1  _14866_
timestamp 0
transform 1 0 11610 0 1 1210
box -6 -8 86 248
use OAI21X1  _14867_
timestamp 0
transform 1 0 11050 0 -1 1210
box -6 -8 106 248
use NOR2X1  _14868_
timestamp 0
transform -1 0 11330 0 1 1210
box -6 -8 86 248
use DFFPOSX1  _14869_
timestamp 0
transform 1 0 13530 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _14870_
timestamp 0
transform 1 0 14410 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _14871_
timestamp 0
transform -1 0 14890 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _14872_
timestamp 0
transform -1 0 13770 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _14873_
timestamp 0
transform -1 0 13370 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _14874_
timestamp 0
transform -1 0 12670 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _14875_
timestamp 0
transform 1 0 11570 0 -1 1690
box -6 -8 246 248
use DFFPOSX1  _14876_
timestamp 0
transform 1 0 14290 0 -1 1690
box -6 -8 246 248
use DFFPOSX1  _14877_
timestamp 0
transform -1 0 15570 0 -1 1690
box -6 -8 246 248
use DFFPOSX1  _14878_
timestamp 0
transform -1 0 14290 0 -1 1690
box -6 -8 246 248
use DFFPOSX1  _14879_
timestamp 0
transform 1 0 13690 0 -1 730
box -6 -8 246 248
use DFFPOSX1  _14880_
timestamp 0
transform -1 0 16630 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _14881_
timestamp 0
transform 1 0 16770 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _14882_
timestamp 0
transform 1 0 16870 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _14883_
timestamp 0
transform -1 0 16630 0 1 730
box -6 -8 246 248
use DFFPOSX1  _14884_
timestamp 0
transform -1 0 15350 0 -1 1210
box -6 -8 246 248
use DFFPOSX1  _14885_
timestamp 0
transform 1 0 14290 0 1 730
box -6 -8 246 248
use DFFPOSX1  _14886_
timestamp 0
transform 1 0 15050 0 1 730
box -6 -8 246 248
use DFFPOSX1  _14887_
timestamp 0
transform -1 0 15830 0 1 730
box -6 -8 246 248
use DFFPOSX1  _14888_
timestamp 0
transform -1 0 12750 0 1 730
box -6 -8 246 248
use DFFPOSX1  _14889_
timestamp 0
transform -1 0 12510 0 1 730
box -6 -8 246 248
use DFFPOSX1  _14890_
timestamp 0
transform -1 0 12750 0 -1 730
box -6 -8 246 248
use DFFPOSX1  _14891_
timestamp 0
transform 1 0 13330 0 1 730
box -6 -8 246 248
use DFFPOSX1  _14892_
timestamp 0
transform -1 0 11990 0 1 730
box -6 -8 246 248
use DFFPOSX1  _14893_
timestamp 0
transform -1 0 11390 0 1 730
box -6 -8 246 248
use DFFPOSX1  _14894_
timestamp 0
transform -1 0 11150 0 1 730
box -6 -8 246 248
use DFFPOSX1  _14895_
timestamp 0
transform -1 0 10910 0 1 730
box -6 -8 246 248
use DFFPOSX1  _14896_
timestamp 0
transform -1 0 12910 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _14897_
timestamp 0
transform 1 0 11390 0 -1 1210
box -6 -8 246 248
use DFFPOSX1  _14898_
timestamp 0
transform -1 0 15770 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _14899_
timestamp 0
transform -1 0 13290 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _14900_
timestamp 0
transform -1 0 15050 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _14901_
timestamp 0
transform -1 0 12810 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _14902_
timestamp 0
transform -1 0 14370 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _14903_
timestamp 0
transform -1 0 13770 0 -1 1690
box -6 -8 246 248
use DFFPOSX1  _14904_
timestamp 0
transform -1 0 12470 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _14905_
timestamp 0
transform 1 0 11390 0 1 730
box -6 -8 246 248
use DFFPOSX1  _14906_
timestamp 0
transform 1 0 11330 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _14907_
timestamp 0
transform -1 0 12330 0 1 1690
box -6 -8 246 248
use BUFX2  _14908_
timestamp 0
transform -1 0 7690 0 -1 6970
box -6 -8 86 248
use BUFX2  _14909_
timestamp 0
transform -1 0 150 0 1 7930
box -6 -8 86 248
use BUFX2  _14910_
timestamp 0
transform -1 0 8590 0 -1 250
box -6 -8 86 248
use BUFX2  _14911_
timestamp 0
transform -1 0 9870 0 1 250
box -6 -8 86 248
use BUFX2  _14912_
timestamp 0
transform -1 0 6870 0 1 6970
box -6 -8 86 248
use BUFX2  _14913_
timestamp 0
transform -1 0 130 0 1 6970
box -6 -8 86 248
use BUFX2  _14914_
timestamp 0
transform 1 0 8270 0 1 6010
box -6 -8 86 248
use BUFX2  _14915_
timestamp 0
transform 1 0 16210 0 -1 250
box -6 -8 86 248
use BUFX2  _14916_
timestamp 0
transform 1 0 8470 0 -1 6010
box -6 -8 86 248
use BUFX2  _14917_
timestamp 0
transform -1 0 8050 0 -1 6010
box -6 -8 86 248
use BUFX2  _14918_
timestamp 0
transform -1 0 8210 0 1 6010
box -6 -8 86 248
use BUFX2  _14919_
timestamp 0
transform -1 0 6390 0 1 7450
box -6 -8 86 248
use BUFX2  _14920_
timestamp 0
transform 1 0 9010 0 -1 250
box -6 -8 86 248
use BUFX2  BUFX2_insert0
timestamp 0
transform 1 0 8230 0 -1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert1
timestamp 0
transform 1 0 9530 0 -1 8410
box -6 -8 86 248
use BUFX2  BUFX2_insert2
timestamp 0
transform -1 0 7930 0 -1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert3
timestamp 0
transform 1 0 9490 0 1 8410
box -6 -8 86 248
use BUFX2  BUFX2_insert4
timestamp 0
transform -1 0 9430 0 1 8410
box -6 -8 86 248
use BUFX2  BUFX2_insert5
timestamp 0
transform 1 0 5450 0 1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert6
timestamp 0
transform 1 0 4650 0 1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert7
timestamp 0
transform -1 0 1410 0 1 10810
box -6 -8 86 248
use BUFX2  BUFX2_insert8
timestamp 0
transform -1 0 1270 0 -1 8410
box -6 -8 86 248
use BUFX2  BUFX2_insert9
timestamp 0
transform 1 0 4550 0 1 6010
box -6 -8 86 248
use BUFX2  BUFX2_insert10
timestamp 0
transform 1 0 4170 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert11
timestamp 0
transform 1 0 3610 0 1 6010
box -6 -8 86 248
use BUFX2  BUFX2_insert12
timestamp 0
transform -1 0 3390 0 -1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert13
timestamp 0
transform -1 0 4530 0 1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert14
timestamp 0
transform -1 0 4190 0 -1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert15
timestamp 0
transform 1 0 6890 0 1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert16
timestamp 0
transform -1 0 4870 0 1 7450
box -6 -8 86 248
use BUFX2  BUFX2_insert17
timestamp 0
transform -1 0 3330 0 1 7450
box -6 -8 86 248
use BUFX2  BUFX2_insert18
timestamp 0
transform -1 0 4610 0 1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert19
timestamp 0
transform -1 0 16230 0 1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert20
timestamp 0
transform -1 0 16370 0 1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert21
timestamp 0
transform -1 0 12970 0 1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert22
timestamp 0
transform -1 0 12210 0 1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert23
timestamp 0
transform -1 0 3110 0 -1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert24
timestamp 0
transform 1 0 4690 0 1 10330
box -6 -8 86 248
use BUFX2  BUFX2_insert25
timestamp 0
transform 1 0 1090 0 -1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert26
timestamp 0
transform -1 0 130 0 1 10810
box -6 -8 86 248
use BUFX2  BUFX2_insert27
timestamp 0
transform -1 0 1290 0 1 10810
box -6 -8 86 248
use BUFX2  BUFX2_insert28
timestamp 0
transform -1 0 130 0 1 10330
box -6 -8 86 248
use BUFX2  BUFX2_insert108
timestamp 0
transform -1 0 7910 0 1 7450
box -6 -8 86 248
use BUFX2  BUFX2_insert109
timestamp 0
transform 1 0 9310 0 1 7450
box -6 -8 86 248
use BUFX2  BUFX2_insert110
timestamp 0
transform -1 0 9130 0 -1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert111
timestamp 0
transform 1 0 8830 0 -1 7450
box -6 -8 86 248
use BUFX2  BUFX2_insert112
timestamp 0
transform 1 0 8330 0 -1 7450
box -6 -8 86 248
use BUFX2  BUFX2_insert113
timestamp 0
transform -1 0 13950 0 -1 14650
box -6 -8 86 248
use BUFX2  BUFX2_insert114
timestamp 0
transform -1 0 13610 0 1 13210
box -6 -8 86 248
use BUFX2  BUFX2_insert115
timestamp 0
transform -1 0 14450 0 -1 12730
box -6 -8 86 248
use BUFX2  BUFX2_insert116
timestamp 0
transform 1 0 15110 0 1 14650
box -6 -8 86 248
use BUFX2  BUFX2_insert117
timestamp 0
transform -1 0 7070 0 -1 6970
box -6 -8 86 248
use BUFX2  BUFX2_insert118
timestamp 0
transform 1 0 8170 0 1 6490
box -6 -8 86 248
use BUFX2  BUFX2_insert119
timestamp 0
transform 1 0 7730 0 -1 6970
box -6 -8 86 248
use BUFX2  BUFX2_insert120
timestamp 0
transform 1 0 7130 0 -1 6970
box -6 -8 86 248
use BUFX2  BUFX2_insert121
timestamp 0
transform -1 0 5890 0 1 6490
box -6 -8 86 248
use BUFX2  BUFX2_insert122
timestamp 0
transform -1 0 7690 0 1 6010
box -6 -8 86 248
use BUFX2  BUFX2_insert123
timestamp 0
transform 1 0 7770 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert124
timestamp 0
transform -1 0 6670 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert125
timestamp 0
transform -1 0 6110 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert126
timestamp 0
transform 1 0 5370 0 1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert127
timestamp 0
transform -1 0 4190 0 -1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert128
timestamp 0
transform 1 0 4630 0 -1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert129
timestamp 0
transform -1 0 4290 0 1 7450
box -6 -8 86 248
use BUFX2  BUFX2_insert130
timestamp 0
transform -1 0 5190 0 -1 8410
box -6 -8 86 248
use BUFX2  BUFX2_insert131
timestamp 0
transform -1 0 2650 0 -1 15130
box -6 -8 86 248
use BUFX2  BUFX2_insert132
timestamp 0
transform 1 0 2710 0 -1 15130
box -6 -8 86 248
use BUFX2  BUFX2_insert133
timestamp 0
transform 1 0 910 0 -1 16570
box -6 -8 86 248
use BUFX2  BUFX2_insert134
timestamp 0
transform -1 0 530 0 -1 16570
box -6 -8 86 248
use BUFX2  BUFX2_insert135
timestamp 0
transform 1 0 630 0 -1 17050
box -6 -8 86 248
use BUFX2  BUFX2_insert136
timestamp 0
transform 1 0 13610 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert137
timestamp 0
transform -1 0 12010 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert138
timestamp 0
transform -1 0 12130 0 1 250
box -6 -8 86 248
use BUFX2  BUFX2_insert139
timestamp 0
transform 1 0 15550 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert140
timestamp 0
transform 1 0 14570 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert141
timestamp 0
transform -1 0 11070 0 1 11290
box -6 -8 86 248
use BUFX2  BUFX2_insert142
timestamp 0
transform 1 0 12150 0 -1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert143
timestamp 0
transform -1 0 11390 0 -1 10330
box -6 -8 86 248
use BUFX2  BUFX2_insert144
timestamp 0
transform 1 0 12230 0 1 11290
box -6 -8 86 248
use BUFX2  BUFX2_insert145
timestamp 0
transform 1 0 12330 0 -1 11290
box -6 -8 86 248
use BUFX2  BUFX2_insert146
timestamp 0
transform -1 0 10630 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert147
timestamp 0
transform 1 0 10670 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert148
timestamp 0
transform 1 0 8530 0 1 250
box -6 -8 86 248
use BUFX2  BUFX2_insert149
timestamp 0
transform 1 0 8110 0 -1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert150
timestamp 0
transform -1 0 8010 0 1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert151
timestamp 0
transform -1 0 16170 0 -1 14170
box -6 -8 86 248
use BUFX2  BUFX2_insert152
timestamp 0
transform 1 0 16070 0 1 13690
box -6 -8 86 248
use BUFX2  BUFX2_insert153
timestamp 0
transform -1 0 16030 0 -1 14170
box -6 -8 86 248
use BUFX2  BUFX2_insert154
timestamp 0
transform -1 0 16010 0 1 12730
box -6 -8 86 248
use BUFX2  BUFX2_insert155
timestamp 0
transform -1 0 16070 0 -1 13210
box -6 -8 86 248
use BUFX2  BUFX2_insert156
timestamp 0
transform -1 0 15830 0 1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert157
timestamp 0
transform -1 0 15110 0 -1 9850
box -6 -8 86 248
use BUFX2  BUFX2_insert158
timestamp 0
transform 1 0 16990 0 -1 9850
box -6 -8 86 248
use BUFX2  BUFX2_insert159
timestamp 0
transform 1 0 15910 0 -1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert160
timestamp 0
transform 1 0 16450 0 -1 9850
box -6 -8 86 248
use BUFX2  BUFX2_insert161
timestamp 0
transform 1 0 11970 0 -1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert162
timestamp 0
transform 1 0 12750 0 -1 9850
box -6 -8 86 248
use BUFX2  BUFX2_insert163
timestamp 0
transform 1 0 12770 0 -1 10330
box -6 -8 86 248
use BUFX2  BUFX2_insert164
timestamp 0
transform -1 0 10610 0 -1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert165
timestamp 0
transform -1 0 11790 0 -1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert166
timestamp 0
transform -1 0 1270 0 1 9850
box -6 -8 86 248
use BUFX2  BUFX2_insert167
timestamp 0
transform -1 0 1250 0 1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert168
timestamp 0
transform 1 0 3670 0 1 9850
box -6 -8 86 248
use BUFX2  BUFX2_insert169
timestamp 0
transform 1 0 3730 0 1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert170
timestamp 0
transform 1 0 1550 0 -1 9850
box -6 -8 86 248
use BUFX2  BUFX2_insert171
timestamp 0
transform -1 0 14510 0 1 12730
box -6 -8 86 248
use BUFX2  BUFX2_insert172
timestamp 0
transform 1 0 12890 0 1 12730
box -6 -8 86 248
use BUFX2  BUFX2_insert173
timestamp 0
transform -1 0 12030 0 1 13690
box -6 -8 86 248
use BUFX2  BUFX2_insert174
timestamp 0
transform -1 0 12190 0 -1 13210
box -6 -8 86 248
use BUFX2  BUFX2_insert175
timestamp 0
transform 1 0 14790 0 1 12250
box -6 -8 86 248
use BUFX2  BUFX2_insert176
timestamp 0
transform -1 0 14110 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert177
timestamp 0
transform 1 0 15890 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert178
timestamp 0
transform -1 0 14130 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert179
timestamp 0
transform 1 0 15870 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert180
timestamp 0
transform 1 0 15270 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert181
timestamp 0
transform 1 0 11510 0 1 6490
box -6 -8 86 248
use BUFX2  BUFX2_insert182
timestamp 0
transform -1 0 10150 0 -1 6010
box -6 -8 86 248
use BUFX2  BUFX2_insert183
timestamp 0
transform 1 0 11750 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert184
timestamp 0
transform 1 0 11850 0 -1 7450
box -6 -8 86 248
use BUFX2  BUFX2_insert185
timestamp 0
transform -1 0 10410 0 -1 7450
box -6 -8 86 248
use BUFX2  BUFX2_insert186
timestamp 0
transform -1 0 6090 0 1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert187
timestamp 0
transform 1 0 8270 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert188
timestamp 0
transform -1 0 6910 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert189
timestamp 0
transform -1 0 6070 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert190
timestamp 0
transform 1 0 9630 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert191
timestamp 0
transform 1 0 12550 0 -1 16570
box -6 -8 86 248
use BUFX2  BUFX2_insert192
timestamp 0
transform 1 0 12410 0 1 14650
box -6 -8 86 248
use BUFX2  BUFX2_insert193
timestamp 0
transform 1 0 12150 0 1 15130
box -6 -8 86 248
use BUFX2  BUFX2_insert194
timestamp 0
transform -1 0 11530 0 -1 15130
box -6 -8 86 248
use BUFX2  BUFX2_insert195
timestamp 0
transform -1 0 11930 0 1 14170
box -6 -8 86 248
use BUFX2  BUFX2_insert196
timestamp 0
transform -1 0 1490 0 1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert197
timestamp 0
transform -1 0 1950 0 1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert198
timestamp 0
transform -1 0 830 0 1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert199
timestamp 0
transform 1 0 1910 0 -1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert200
timestamp 0
transform 1 0 12770 0 1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert201
timestamp 0
transform -1 0 11990 0 1 10810
box -6 -8 86 248
use BUFX2  BUFX2_insert202
timestamp 0
transform 1 0 12850 0 1 10810
box -6 -8 86 248
use BUFX2  BUFX2_insert203
timestamp 0
transform -1 0 12710 0 -1 10330
box -6 -8 86 248
use BUFX2  BUFX2_insert204
timestamp 0
transform -1 0 12590 0 -1 10810
box -6 -8 86 248
use BUFX2  BUFX2_insert205
timestamp 0
transform 1 0 12070 0 1 5530
box -6 -8 86 248
use BUFX2  BUFX2_insert206
timestamp 0
transform 1 0 14070 0 1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert207
timestamp 0
transform -1 0 11910 0 1 5530
box -6 -8 86 248
use BUFX2  BUFX2_insert208
timestamp 0
transform 1 0 15530 0 1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert209
timestamp 0
transform 1 0 170 0 1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert210
timestamp 0
transform 1 0 1170 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert211
timestamp 0
transform 1 0 330 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert212
timestamp 0
transform -1 0 870 0 -1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert213
timestamp 0
transform -1 0 150 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert214
timestamp 0
transform 1 0 6430 0 1 6970
box -6 -8 86 248
use BUFX2  BUFX2_insert215
timestamp 0
transform -1 0 5830 0 -1 6970
box -6 -8 86 248
use BUFX2  BUFX2_insert216
timestamp 0
transform -1 0 4890 0 -1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert217
timestamp 0
transform -1 0 3570 0 1 6970
box -6 -8 86 248
use BUFX2  BUFX2_insert218
timestamp 0
transform 1 0 6730 0 -1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert219
timestamp 0
transform -1 0 11650 0 1 5530
box -6 -8 86 248
use BUFX2  BUFX2_insert220
timestamp 0
transform 1 0 11790 0 -1 6490
box -6 -8 86 248
use BUFX2  BUFX2_insert221
timestamp 0
transform -1 0 12190 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert222
timestamp 0
transform -1 0 10070 0 -1 6490
box -6 -8 86 248
use BUFX2  BUFX2_insert223
timestamp 0
transform 1 0 12310 0 -1 6490
box -6 -8 86 248
use BUFX2  BUFX2_insert224
timestamp 0
transform -1 0 9030 0 1 14170
box -6 -8 86 248
use BUFX2  BUFX2_insert225
timestamp 0
transform 1 0 6990 0 -1 16570
box -6 -8 86 248
use BUFX2  BUFX2_insert226
timestamp 0
transform -1 0 10650 0 1 15610
box -6 -8 86 248
use BUFX2  BUFX2_insert227
timestamp 0
transform -1 0 6950 0 1 15130
box -6 -8 86 248
use BUFX2  BUFX2_insert228
timestamp 0
transform -1 0 7630 0 -1 16090
box -6 -8 86 248
use BUFX2  BUFX2_insert229
timestamp 0
transform 1 0 9010 0 -1 15130
box -6 -8 86 248
use BUFX2  BUFX2_insert230
timestamp 0
transform 1 0 8750 0 -1 15130
box -6 -8 86 248
use BUFX2  BUFX2_insert231
timestamp 0
transform -1 0 7530 0 1 16090
box -6 -8 86 248
use BUFX2  BUFX2_insert232
timestamp 0
transform -1 0 9030 0 1 15130
box -6 -8 86 248
use BUFX2  BUFX2_insert233
timestamp 0
transform -1 0 15230 0 1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert234
timestamp 0
transform 1 0 15410 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert235
timestamp 0
transform -1 0 13010 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert236
timestamp 0
transform -1 0 12210 0 -1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert237
timestamp 0
transform -1 0 13330 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert238
timestamp 0
transform -1 0 2370 0 -1 12250
box -6 -8 86 248
use BUFX2  BUFX2_insert239
timestamp 0
transform -1 0 4770 0 1 13210
box -6 -8 86 248
use BUFX2  BUFX2_insert240
timestamp 0
transform 1 0 5230 0 -1 12250
box -6 -8 86 248
use BUFX2  BUFX2_insert241
timestamp 0
transform 1 0 5670 0 -1 14170
box -6 -8 86 248
use BUFX2  BUFX2_insert242
timestamp 0
transform 1 0 5430 0 -1 12730
box -6 -8 86 248
use BUFX2  BUFX2_insert243
timestamp 0
transform -1 0 1930 0 1 5530
box -6 -8 86 248
use BUFX2  BUFX2_insert244
timestamp 0
transform -1 0 1510 0 1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert245
timestamp 0
transform 1 0 4490 0 1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert246
timestamp 0
transform 1 0 2470 0 1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert247
timestamp 0
transform 1 0 3890 0 1 5530
box -6 -8 86 248
use BUFX2  BUFX2_insert248
timestamp 0
transform 1 0 2290 0 -1 16090
box -6 -8 86 248
use BUFX2  BUFX2_insert249
timestamp 0
transform 1 0 3290 0 -1 14650
box -6 -8 86 248
use BUFX2  BUFX2_insert250
timestamp 0
transform -1 0 530 0 -1 16090
box -6 -8 86 248
use BUFX2  BUFX2_insert251
timestamp 0
transform -1 0 2010 0 -1 15610
box -6 -8 86 248
use BUFX2  BUFX2_insert252
timestamp 0
transform 1 0 3070 0 -1 15130
box -6 -8 86 248
use BUFX2  BUFX2_insert253
timestamp 0
transform 1 0 8670 0 1 6010
box -6 -8 86 248
use BUFX2  BUFX2_insert254
timestamp 0
transform 1 0 11390 0 -1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert255
timestamp 0
transform -1 0 10310 0 1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert256
timestamp 0
transform 1 0 11150 0 1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert257
timestamp 0
transform 1 0 12070 0 1 6010
box -6 -8 86 248
use BUFX2  BUFX2_insert258
timestamp 0
transform -1 0 14090 0 -1 14650
box -6 -8 86 248
use BUFX2  BUFX2_insert259
timestamp 0
transform -1 0 13830 0 -1 13690
box -6 -8 86 248
use BUFX2  BUFX2_insert260
timestamp 0
transform 1 0 16510 0 1 15610
box -6 -8 86 248
use BUFX2  BUFX2_insert261
timestamp 0
transform -1 0 15950 0 -1 16090
box -6 -8 86 248
use BUFX2  BUFX2_insert262
timestamp 0
transform -1 0 13530 0 -1 16090
box -6 -8 86 248
use BUFX2  BUFX2_insert263
timestamp 0
transform -1 0 13450 0 1 13690
box -6 -8 86 248
use BUFX2  BUFX2_insert264
timestamp 0
transform 1 0 4570 0 1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert265
timestamp 0
transform 1 0 5470 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert266
timestamp 0
transform -1 0 4370 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert267
timestamp 0
transform -1 0 4490 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert268
timestamp 0
transform -1 0 4470 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert269
timestamp 0
transform -1 0 7610 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert270
timestamp 0
transform -1 0 7290 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert271
timestamp 0
transform 1 0 9870 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert272
timestamp 0
transform 1 0 8110 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert273
timestamp 0
transform 1 0 9030 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert274
timestamp 0
transform -1 0 8350 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert275
timestamp 0
transform 1 0 9910 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert276
timestamp 0
transform 1 0 9710 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert277
timestamp 0
transform -1 0 7130 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert278
timestamp 0
transform 1 0 7470 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert279
timestamp 0
transform 1 0 9950 0 1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert280
timestamp 0
transform -1 0 16010 0 1 14170
box -6 -8 86 248
use BUFX2  BUFX2_insert281
timestamp 0
transform -1 0 15950 0 -1 13210
box -6 -8 86 248
use BUFX2  BUFX2_insert282
timestamp 0
transform 1 0 15950 0 1 13690
box -6 -8 86 248
use BUFX2  BUFX2_insert283
timestamp 0
transform -1 0 16670 0 1 14170
box -6 -8 86 248
use BUFX2  BUFX2_insert284
timestamp 0
transform 1 0 16130 0 -1 13210
box -6 -8 86 248
use BUFX2  BUFX2_insert285
timestamp 0
transform -1 0 15950 0 1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert286
timestamp 0
transform -1 0 16410 0 1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert287
timestamp 0
transform 1 0 16410 0 1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert288
timestamp 0
transform 1 0 15090 0 1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert289
timestamp 0
transform -1 0 13110 0 1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert290
timestamp 0
transform 1 0 6750 0 1 12730
box -6 -8 86 248
use BUFX2  BUFX2_insert291
timestamp 0
transform 1 0 6630 0 1 12730
box -6 -8 86 248
use BUFX2  BUFX2_insert292
timestamp 0
transform -1 0 6570 0 1 12730
box -6 -8 86 248
use BUFX2  BUFX2_insert293
timestamp 0
transform 1 0 8310 0 1 12730
box -6 -8 86 248
use BUFX2  BUFX2_insert294
timestamp 0
transform -1 0 11970 0 -1 8410
box -6 -8 86 248
use BUFX2  BUFX2_insert295
timestamp 0
transform -1 0 11970 0 1 10330
box -6 -8 86 248
use BUFX2  BUFX2_insert296
timestamp 0
transform 1 0 15270 0 -1 8410
box -6 -8 86 248
use BUFX2  BUFX2_insert297
timestamp 0
transform 1 0 15030 0 -1 10330
box -6 -8 86 248
use BUFX2  BUFX2_insert298
timestamp 0
transform 1 0 17090 0 1 10330
box -6 -8 86 248
use BUFX2  BUFX2_insert299
timestamp 0
transform 1 0 16950 0 -1 8410
box -6 -8 86 248
use BUFX2  BUFX2_insert300
timestamp 0
transform 1 0 9130 0 1 14650
box -6 -8 86 248
use BUFX2  BUFX2_insert301
timestamp 0
transform -1 0 8090 0 -1 12730
box -6 -8 86 248
use BUFX2  BUFX2_insert302
timestamp 0
transform -1 0 8150 0 1 14650
box -6 -8 86 248
use BUFX2  BUFX2_insert303
timestamp 0
transform -1 0 8150 0 1 12730
box -6 -8 86 248
use BUFX2  BUFX2_insert304
timestamp 0
transform -1 0 8650 0 1 6970
box -6 -8 86 248
use BUFX2  BUFX2_insert305
timestamp 0
transform 1 0 8630 0 1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert306
timestamp 0
transform -1 0 9790 0 -1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert307
timestamp 0
transform 1 0 9730 0 1 6970
box -6 -8 86 248
use BUFX2  BUFX2_insert308
timestamp 0
transform 1 0 10250 0 1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert309
timestamp 0
transform -1 0 13730 0 -1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert310
timestamp 0
transform 1 0 13790 0 -1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert311
timestamp 0
transform -1 0 15990 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert312
timestamp 0
transform -1 0 16070 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert313
timestamp 0
transform -1 0 15190 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert314
timestamp 0
transform 1 0 15630 0 -1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert315
timestamp 0
transform 1 0 16430 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert316
timestamp 0
transform 1 0 14270 0 -1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert317
timestamp 0
transform 1 0 16390 0 1 5530
box -6 -8 86 248
use BUFX2  BUFX2_insert318
timestamp 0
transform -1 0 11790 0 1 5530
box -6 -8 86 248
use BUFX2  BUFX2_insert319
timestamp 0
transform 1 0 11950 0 1 5530
box -6 -8 86 248
use BUFX2  BUFX2_insert320
timestamp 0
transform 1 0 8610 0 -1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert321
timestamp 0
transform -1 0 7030 0 -1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert322
timestamp 0
transform 1 0 7070 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert323
timestamp 0
transform 1 0 8670 0 -1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert324
timestamp 0
transform -1 0 730 0 -1 14170
box -6 -8 86 248
use BUFX2  BUFX2_insert325
timestamp 0
transform 1 0 3010 0 -1 12730
box -6 -8 86 248
use BUFX2  BUFX2_insert326
timestamp 0
transform 1 0 2110 0 -1 16570
box -6 -8 86 248
use BUFX2  BUFX2_insert327
timestamp 0
transform -1 0 2990 0 1 15130
box -6 -8 86 248
use BUFX2  BUFX2_insert328
timestamp 0
transform 1 0 1070 0 1 15610
box -6 -8 86 248
use BUFX2  BUFX2_insert329
timestamp 0
transform 1 0 2090 0 1 16570
box -6 -8 86 248
use BUFX2  BUFX2_insert330
timestamp 0
transform -1 0 2950 0 1 15610
box -6 -8 86 248
use BUFX2  BUFX2_insert331
timestamp 0
transform 1 0 3770 0 1 14170
box -6 -8 86 248
use BUFX2  BUFX2_insert332
timestamp 0
transform -1 0 2930 0 1 12730
box -6 -8 86 248
use BUFX2  BUFX2_insert333
timestamp 0
transform -1 0 1890 0 1 15130
box -6 -8 86 248
use BUFX2  BUFX2_insert334
timestamp 0
transform 1 0 2850 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert335
timestamp 0
transform 1 0 2590 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert336
timestamp 0
transform 1 0 330 0 1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert337
timestamp 0
transform -1 0 1270 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert338
timestamp 0
transform -1 0 1610 0 1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert339
timestamp 0
transform -1 0 910 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert340
timestamp 0
transform 1 0 330 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert341
timestamp 0
transform -1 0 650 0 -1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert342
timestamp 0
transform 1 0 1210 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert343
timestamp 0
transform 1 0 210 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert344
timestamp 0
transform -1 0 150 0 -1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert345
timestamp 0
transform 1 0 10890 0 -1 16570
box -6 -8 86 248
use BUFX2  BUFX2_insert346
timestamp 0
transform -1 0 11170 0 -1 13690
box -6 -8 86 248
use BUFX2  BUFX2_insert347
timestamp 0
transform 1 0 11510 0 1 15130
box -6 -8 86 248
use BUFX2  BUFX2_insert348
timestamp 0
transform -1 0 11010 0 1 13690
box -6 -8 86 248
use BUFX2  BUFX2_insert349
timestamp 0
transform 1 0 8130 0 -1 16090
box -6 -8 86 248
use BUFX2  BUFX2_insert350
timestamp 0
transform -1 0 7890 0 -1 16090
box -6 -8 86 248
use BUFX2  BUFX2_insert351
timestamp 0
transform -1 0 7730 0 1 15130
box -6 -8 86 248
use BUFX2  BUFX2_insert352
timestamp 0
transform 1 0 7770 0 1 15130
box -6 -8 86 248
use BUFX2  BUFX2_insert353
timestamp 0
transform 1 0 10770 0 -1 14650
box -6 -8 86 248
use BUFX2  BUFX2_insert354
timestamp 0
transform -1 0 6550 0 1 16090
box -6 -8 86 248
use BUFX2  BUFX2_insert355
timestamp 0
transform -1 0 9530 0 -1 14170
box -6 -8 86 248
use BUFX2  BUFX2_insert356
timestamp 0
transform 1 0 9490 0 1 16090
box -6 -8 86 248
use BUFX2  BUFX2_insert357
timestamp 0
transform -1 0 7130 0 -1 14170
box -6 -8 86 248
use BUFX2  BUFX2_insert358
timestamp 0
transform 1 0 10810 0 1 13690
box -6 -8 86 248
use BUFX2  BUFX2_insert359
timestamp 0
transform -1 0 9550 0 1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert360
timestamp 0
transform -1 0 7590 0 1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert361
timestamp 0
transform -1 0 6410 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert362
timestamp 0
transform -1 0 8250 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert363
timestamp 0
transform 1 0 6710 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert364
timestamp 0
transform 1 0 3490 0 1 11770
box -6 -8 86 248
use BUFX2  BUFX2_insert365
timestamp 0
transform -1 0 4910 0 1 13210
box -6 -8 86 248
use BUFX2  BUFX2_insert366
timestamp 0
transform -1 0 3750 0 1 13210
box -6 -8 86 248
use BUFX2  BUFX2_insert367
timestamp 0
transform -1 0 3050 0 -1 13210
box -6 -8 86 248
use BUFX2  BUFX2_insert368
timestamp 0
transform -1 0 4850 0 -1 12250
box -6 -8 86 248
use BUFX2  BUFX2_insert369
timestamp 0
transform 1 0 13350 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert370
timestamp 0
transform -1 0 13010 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert371
timestamp 0
transform 1 0 12050 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert372
timestamp 0
transform 1 0 13230 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert373
timestamp 0
transform -1 0 11270 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert374
timestamp 0
transform 1 0 2890 0 1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert375
timestamp 0
transform 1 0 3030 0 1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert376
timestamp 0
transform -1 0 1530 0 1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert377
timestamp 0
transform -1 0 2090 0 1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert378
timestamp 0
transform -1 0 1410 0 -1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert379
timestamp 0
transform 1 0 6370 0 1 11770
box -6 -8 86 248
use BUFX2  BUFX2_insert380
timestamp 0
transform 1 0 4970 0 1 13210
box -6 -8 86 248
use BUFX2  BUFX2_insert381
timestamp 0
transform -1 0 2950 0 -1 12730
box -6 -8 86 248
use BUFX2  BUFX2_insert382
timestamp 0
transform 1 0 5790 0 1 11290
box -6 -8 86 248
use BUFX2  BUFX2_insert383
timestamp 0
transform -1 0 4590 0 1 11290
box -6 -8 86 248
use CLKBUF1  CLKBUF1_insert29
timestamp 0
transform -1 0 9630 0 1 4570
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert30
timestamp 0
transform 1 0 10490 0 1 16570
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert31
timestamp 0
transform -1 0 1950 0 1 5050
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert32
timestamp 0
transform -1 0 6430 0 1 12250
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert33
timestamp 0
transform -1 0 5990 0 -1 14170
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert34
timestamp 0
transform -1 0 10270 0 1 7450
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert35
timestamp 0
transform -1 0 13390 0 -1 2170
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert36
timestamp 0
transform 1 0 3550 0 -1 8410
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert37
timestamp 0
transform -1 0 14890 0 -1 12250
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert38
timestamp 0
transform 1 0 5650 0 1 10810
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert39
timestamp 0
transform -1 0 6090 0 -1 6970
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert40
timestamp 0
transform 1 0 15910 0 -1 2170
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert41
timestamp 0
transform -1 0 11530 0 1 3130
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert42
timestamp 0
transform 1 0 9490 0 1 11290
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert43
timestamp 0
transform 1 0 7390 0 -1 9850
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert44
timestamp 0
transform 1 0 2790 0 -1 4570
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert45
timestamp 0
transform 1 0 11070 0 -1 15130
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert46
timestamp 0
transform 1 0 3530 0 1 6490
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert47
timestamp 0
transform 1 0 13010 0 1 7930
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert48
timestamp 0
transform -1 0 2310 0 -1 12730
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert49
timestamp 0
transform 1 0 6130 0 -1 6970
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert50
timestamp 0
transform -1 0 13690 0 -1 12250
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert51
timestamp 0
transform 1 0 14750 0 1 13690
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert52
timestamp 0
transform -1 0 7230 0 -1 7930
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert53
timestamp 0
transform -1 0 4470 0 -1 9850
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert54
timestamp 0
transform 1 0 13130 0 1 6970
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert55
timestamp 0
transform 1 0 14190 0 1 12730
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert56
timestamp 0
transform -1 0 11390 0 1 7930
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert57
timestamp 0
transform -1 0 14890 0 1 1690
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert58
timestamp 0
transform 1 0 7190 0 -1 11770
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert59
timestamp 0
transform -1 0 6050 0 -1 8890
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert60
timestamp 0
transform -1 0 9070 0 -1 11290
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert61
timestamp 0
transform 1 0 6370 0 -1 6970
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert62
timestamp 0
transform 1 0 11210 0 1 7450
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert63
timestamp 0
transform 1 0 10370 0 1 12250
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert64
timestamp 0
transform 1 0 3810 0 -1 5050
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert65
timestamp 0
transform 1 0 6970 0 1 2170
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert66
timestamp 0
transform 1 0 10590 0 1 16090
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert67
timestamp 0
transform -1 0 15430 0 -1 2170
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert68
timestamp 0
transform -1 0 6450 0 1 14170
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert69
timestamp 0
transform 1 0 6950 0 -1 10810
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert70
timestamp 0
transform 1 0 3070 0 -1 5050
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert71
timestamp 0
transform -1 0 2810 0 1 11770
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert72
timestamp 0
transform 1 0 9450 0 -1 4090
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert73
timestamp 0
transform 1 0 12410 0 -1 2650
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert74
timestamp 0
transform 1 0 15310 0 -1 12250
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert75
timestamp 0
transform 1 0 10370 0 -1 11770
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert76
timestamp 0
transform 1 0 8330 0 -1 3610
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert77
timestamp 0
transform 1 0 11450 0 1 7930
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert78
timestamp 0
transform 1 0 10850 0 1 15610
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert79
timestamp 0
transform 1 0 11410 0 1 4570
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert80
timestamp 0
transform 1 0 4530 0 -1 4570
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert81
timestamp 0
transform -1 0 5530 0 1 13210
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert82
timestamp 0
transform 1 0 11990 0 -1 7450
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert83
timestamp 0
transform -1 0 2010 0 1 6490
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert84
timestamp 0
transform 1 0 8490 0 1 11290
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert85
timestamp 0
transform -1 0 5490 0 -1 13690
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert86
timestamp 0
transform 1 0 12630 0 1 3130
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert87
timestamp 0
transform -1 0 12250 0 1 7450
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert88
timestamp 0
transform 1 0 8090 0 -1 11290
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert89
timestamp 0
transform 1 0 6550 0 -1 3610
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert90
timestamp 0
transform -1 0 2990 0 1 13210
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert91
timestamp 0
transform -1 0 2350 0 -1 3610
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert92
timestamp 0
transform 1 0 9390 0 1 3610
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert93
timestamp 0
transform -1 0 2330 0 1 7450
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert94
timestamp 0
transform -1 0 4330 0 1 4090
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert95
timestamp 0
transform -1 0 3290 0 1 11770
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert96
timestamp 0
transform -1 0 9210 0 1 5050
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert97
timestamp 0
transform -1 0 9450 0 -1 12250
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert98
timestamp 0
transform -1 0 8330 0 -1 6490
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert99
timestamp 0
transform -1 0 10110 0 -1 4570
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert100
timestamp 0
transform 1 0 11650 0 1 4570
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert101
timestamp 0
transform -1 0 15150 0 -1 12250
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert102
timestamp 0
transform 1 0 12290 0 1 7450
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert103
timestamp 0
transform -1 0 10350 0 1 6970
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert104
timestamp 0
transform -1 0 6390 0 -1 10810
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert105
timestamp 0
transform -1 0 6790 0 1 2170
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert106
timestamp 0
transform -1 0 2410 0 -1 5050
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert107
timestamp 0
transform 1 0 9730 0 1 11290
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert384
timestamp 0
transform 1 0 8950 0 -1 17050
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert385
timestamp 0
transform -1 0 5770 0 1 6490
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert386
timestamp 0
transform -1 0 4870 0 1 5050
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert387
timestamp 0
transform 1 0 10810 0 1 7450
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert388
timestamp 0
transform -1 0 8050 0 -1 11290
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert389
timestamp 0
transform 1 0 8410 0 1 6010
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert390
timestamp 0
transform -1 0 10550 0 1 4570
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert391
timestamp 0
transform -1 0 7250 0 1 10810
box -6 -8 206 248
use FILL  FILL256050x21750
timestamp 0
transform -1 0 17090 0 -1 1690
box -6 -8 26 248
use FILL  FILL256050x64950
timestamp 0
transform -1 0 17090 0 -1 4570
box -6 -8 26 248
use FILL  FILL256050x144150
timestamp 0
transform -1 0 17090 0 -1 9850
box -6 -8 26 248
use FILL  FILL256050x216150
timestamp 0
transform -1 0 17090 0 -1 14650
box -6 -8 26 248
use FILL  FILL256050x219750
timestamp 0
transform 1 0 17070 0 1 14650
box -6 -8 26 248
use FILL  FILL256050x223350
timestamp 0
transform -1 0 17090 0 -1 15130
box -6 -8 26 248
use FILL  FILL256050x252150
timestamp 0
transform -1 0 17090 0 -1 17050
box -6 -8 26 248
use FILL  FILL256350x21750
timestamp 0
transform -1 0 17110 0 -1 1690
box -6 -8 26 248
use FILL  FILL256350x28950
timestamp 0
transform -1 0 17110 0 -1 2170
box -6 -8 26 248
use FILL  FILL256350x43350
timestamp 0
transform -1 0 17110 0 -1 3130
box -6 -8 26 248
use FILL  FILL256350x57750
timestamp 0
transform -1 0 17110 0 -1 4090
box -6 -8 26 248
use FILL  FILL256350x64950
timestamp 0
transform -1 0 17110 0 -1 4570
box -6 -8 26 248
use FILL  FILL256350x75750
timestamp 0
transform 1 0 17090 0 1 5050
box -6 -8 26 248
use FILL  FILL256350x108150
timestamp 0
transform -1 0 17110 0 -1 7450
box -6 -8 26 248
use FILL  FILL256350x144150
timestamp 0
transform -1 0 17110 0 -1 9850
box -6 -8 26 248
use FILL  FILL256350x201750
timestamp 0
transform -1 0 17110 0 -1 13690
box -6 -8 26 248
use FILL  FILL256350x216150
timestamp 0
transform -1 0 17110 0 -1 14650
box -6 -8 26 248
use FILL  FILL256350x219750
timestamp 0
transform 1 0 17090 0 1 14650
box -6 -8 26 248
use FILL  FILL256350x223350
timestamp 0
transform -1 0 17110 0 -1 15130
box -6 -8 26 248
use FILL  FILL256350x252150
timestamp 0
transform -1 0 17110 0 -1 17050
box -6 -8 26 248
use FILL  FILL256650x150
timestamp 0
transform -1 0 17130 0 -1 250
box -6 -8 26 248
use FILL  FILL256650x3750
timestamp 0
transform 1 0 17110 0 1 250
box -6 -8 26 248
use FILL  FILL256650x7350
timestamp 0
transform -1 0 17130 0 -1 730
box -6 -8 26 248
use FILL  FILL256650x18150
timestamp 0
transform 1 0 17110 0 1 1210
box -6 -8 26 248
use FILL  FILL256650x21750
timestamp 0
transform -1 0 17130 0 -1 1690
box -6 -8 26 248
use FILL  FILL256650x28950
timestamp 0
transform -1 0 17130 0 -1 2170
box -6 -8 26 248
use FILL  FILL256650x43350
timestamp 0
transform -1 0 17130 0 -1 3130
box -6 -8 26 248
use FILL  FILL256650x57750
timestamp 0
transform -1 0 17130 0 -1 4090
box -6 -8 26 248
use FILL  FILL256650x64950
timestamp 0
transform -1 0 17130 0 -1 4570
box -6 -8 26 248
use FILL  FILL256650x72150
timestamp 0
transform -1 0 17130 0 -1 5050
box -6 -8 26 248
use FILL  FILL256650x75750
timestamp 0
transform 1 0 17110 0 1 5050
box -6 -8 26 248
use FILL  FILL256650x86550
timestamp 0
transform -1 0 17130 0 -1 6010
box -6 -8 26 248
use FILL  FILL256650x108150
timestamp 0
transform -1 0 17130 0 -1 7450
box -6 -8 26 248
use FILL  FILL256650x111750
timestamp 0
transform 1 0 17110 0 1 7450
box -6 -8 26 248
use FILL  FILL256650x126150
timestamp 0
transform 1 0 17110 0 1 8410
box -6 -8 26 248
use FILL  FILL256650x136950
timestamp 0
transform -1 0 17130 0 -1 9370
box -6 -8 26 248
use FILL  FILL256650x144150
timestamp 0
transform -1 0 17130 0 -1 9850
box -6 -8 26 248
use FILL  FILL256650x183750
timestamp 0
transform 1 0 17110 0 1 12250
box -6 -8 26 248
use FILL  FILL256650x198150
timestamp 0
transform 1 0 17110 0 1 13210
box -6 -8 26 248
use FILL  FILL256650x201750
timestamp 0
transform -1 0 17130 0 -1 13690
box -6 -8 26 248
use FILL  FILL256650x216150
timestamp 0
transform -1 0 17130 0 -1 14650
box -6 -8 26 248
use FILL  FILL256650x219750
timestamp 0
transform 1 0 17110 0 1 14650
box -6 -8 26 248
use FILL  FILL256650x223350
timestamp 0
transform -1 0 17130 0 -1 15130
box -6 -8 26 248
use FILL  FILL256650x248550
timestamp 0
transform 1 0 17110 0 1 16570
box -6 -8 26 248
use FILL  FILL256650x252150
timestamp 0
transform -1 0 17130 0 -1 17050
box -6 -8 26 248
use FILL  FILL256950x150
timestamp 0
transform -1 0 17150 0 -1 250
box -6 -8 26 248
use FILL  FILL256950x3750
timestamp 0
transform 1 0 17130 0 1 250
box -6 -8 26 248
use FILL  FILL256950x7350
timestamp 0
transform -1 0 17150 0 -1 730
box -6 -8 26 248
use FILL  FILL256950x10950
timestamp 0
transform 1 0 17130 0 1 730
box -6 -8 26 248
use FILL  FILL256950x18150
timestamp 0
transform 1 0 17130 0 1 1210
box -6 -8 26 248
use FILL  FILL256950x21750
timestamp 0
transform -1 0 17150 0 -1 1690
box -6 -8 26 248
use FILL  FILL256950x28950
timestamp 0
transform -1 0 17150 0 -1 2170
box -6 -8 26 248
use FILL  FILL256950x36150
timestamp 0
transform -1 0 17150 0 -1 2650
box -6 -8 26 248
use FILL  FILL256950x43350
timestamp 0
transform -1 0 17150 0 -1 3130
box -6 -8 26 248
use FILL  FILL256950x46950
timestamp 0
transform 1 0 17130 0 1 3130
box -6 -8 26 248
use FILL  FILL256950x57750
timestamp 0
transform -1 0 17150 0 -1 4090
box -6 -8 26 248
use FILL  FILL256950x64950
timestamp 0
transform -1 0 17150 0 -1 4570
box -6 -8 26 248
use FILL  FILL256950x68550
timestamp 0
transform 1 0 17130 0 1 4570
box -6 -8 26 248
use FILL  FILL256950x72150
timestamp 0
transform -1 0 17150 0 -1 5050
box -6 -8 26 248
use FILL  FILL256950x75750
timestamp 0
transform 1 0 17130 0 1 5050
box -6 -8 26 248
use FILL  FILL256950x86550
timestamp 0
transform -1 0 17150 0 -1 6010
box -6 -8 26 248
use FILL  FILL256950x93750
timestamp 0
transform -1 0 17150 0 -1 6490
box -6 -8 26 248
use FILL  FILL256950x104550
timestamp 0
transform 1 0 17130 0 1 6970
box -6 -8 26 248
use FILL  FILL256950x108150
timestamp 0
transform -1 0 17150 0 -1 7450
box -6 -8 26 248
use FILL  FILL256950x111750
timestamp 0
transform 1 0 17130 0 1 7450
box -6 -8 26 248
use FILL  FILL256950x115350
timestamp 0
transform -1 0 17150 0 -1 7930
box -6 -8 26 248
use FILL  FILL256950x122550
timestamp 0
transform -1 0 17150 0 -1 8410
box -6 -8 26 248
use FILL  FILL256950x126150
timestamp 0
transform 1 0 17130 0 1 8410
box -6 -8 26 248
use FILL  FILL256950x136950
timestamp 0
transform -1 0 17150 0 -1 9370
box -6 -8 26 248
use FILL  FILL256950x140550
timestamp 0
transform 1 0 17130 0 1 9370
box -6 -8 26 248
use FILL  FILL256950x144150
timestamp 0
transform -1 0 17150 0 -1 9850
box -6 -8 26 248
use FILL  FILL256950x147750
timestamp 0
transform 1 0 17130 0 1 9850
box -6 -8 26 248
use FILL  FILL256950x165750
timestamp 0
transform -1 0 17150 0 -1 11290
box -6 -8 26 248
use FILL  FILL256950x169350
timestamp 0
transform 1 0 17130 0 1 11290
box -6 -8 26 248
use FILL  FILL256950x176550
timestamp 0
transform 1 0 17130 0 1 11770
box -6 -8 26 248
use FILL  FILL256950x183750
timestamp 0
transform 1 0 17130 0 1 12250
box -6 -8 26 248
use FILL  FILL256950x198150
timestamp 0
transform 1 0 17130 0 1 13210
box -6 -8 26 248
use FILL  FILL256950x201750
timestamp 0
transform -1 0 17150 0 -1 13690
box -6 -8 26 248
use FILL  FILL256950x208950
timestamp 0
transform -1 0 17150 0 -1 14170
box -6 -8 26 248
use FILL  FILL256950x216150
timestamp 0
transform -1 0 17150 0 -1 14650
box -6 -8 26 248
use FILL  FILL256950x219750
timestamp 0
transform 1 0 17130 0 1 14650
box -6 -8 26 248
use FILL  FILL256950x223350
timestamp 0
transform -1 0 17150 0 -1 15130
box -6 -8 26 248
use FILL  FILL256950x230550
timestamp 0
transform -1 0 17150 0 -1 15610
box -6 -8 26 248
use FILL  FILL256950x237750
timestamp 0
transform -1 0 17150 0 -1 16090
box -6 -8 26 248
use FILL  FILL256950x241350
timestamp 0
transform 1 0 17130 0 1 16090
box -6 -8 26 248
use FILL  FILL256950x244950
timestamp 0
transform -1 0 17150 0 -1 16570
box -6 -8 26 248
use FILL  FILL256950x248550
timestamp 0
transform 1 0 17130 0 1 16570
box -6 -8 26 248
use FILL  FILL256950x252150
timestamp 0
transform -1 0 17150 0 -1 17050
box -6 -8 26 248
use FILL  FILL257250x150
timestamp 0
transform -1 0 17170 0 -1 250
box -6 -8 26 248
use FILL  FILL257250x3750
timestamp 0
transform 1 0 17150 0 1 250
box -6 -8 26 248
use FILL  FILL257250x7350
timestamp 0
transform -1 0 17170 0 -1 730
box -6 -8 26 248
use FILL  FILL257250x10950
timestamp 0
transform 1 0 17150 0 1 730
box -6 -8 26 248
use FILL  FILL257250x18150
timestamp 0
transform 1 0 17150 0 1 1210
box -6 -8 26 248
use FILL  FILL257250x21750
timestamp 0
transform -1 0 17170 0 -1 1690
box -6 -8 26 248
use FILL  FILL257250x25350
timestamp 0
transform 1 0 17150 0 1 1690
box -6 -8 26 248
use FILL  FILL257250x28950
timestamp 0
transform -1 0 17170 0 -1 2170
box -6 -8 26 248
use FILL  FILL257250x36150
timestamp 0
transform -1 0 17170 0 -1 2650
box -6 -8 26 248
use FILL  FILL257250x43350
timestamp 0
transform -1 0 17170 0 -1 3130
box -6 -8 26 248
use FILL  FILL257250x46950
timestamp 0
transform 1 0 17150 0 1 3130
box -6 -8 26 248
use FILL  FILL257250x50550
timestamp 0
transform -1 0 17170 0 -1 3610
box -6 -8 26 248
use FILL  FILL257250x54150
timestamp 0
transform 1 0 17150 0 1 3610
box -6 -8 26 248
use FILL  FILL257250x57750
timestamp 0
transform -1 0 17170 0 -1 4090
box -6 -8 26 248
use FILL  FILL257250x61350
timestamp 0
transform 1 0 17150 0 1 4090
box -6 -8 26 248
use FILL  FILL257250x64950
timestamp 0
transform -1 0 17170 0 -1 4570
box -6 -8 26 248
use FILL  FILL257250x68550
timestamp 0
transform 1 0 17150 0 1 4570
box -6 -8 26 248
use FILL  FILL257250x72150
timestamp 0
transform -1 0 17170 0 -1 5050
box -6 -8 26 248
use FILL  FILL257250x75750
timestamp 0
transform 1 0 17150 0 1 5050
box -6 -8 26 248
use FILL  FILL257250x79350
timestamp 0
transform -1 0 17170 0 -1 5530
box -6 -8 26 248
use FILL  FILL257250x86550
timestamp 0
transform -1 0 17170 0 -1 6010
box -6 -8 26 248
use FILL  FILL257250x90150
timestamp 0
transform 1 0 17150 0 1 6010
box -6 -8 26 248
use FILL  FILL257250x93750
timestamp 0
transform -1 0 17170 0 -1 6490
box -6 -8 26 248
use FILL  FILL257250x100950
timestamp 0
transform -1 0 17170 0 -1 6970
box -6 -8 26 248
use FILL  FILL257250x104550
timestamp 0
transform 1 0 17150 0 1 6970
box -6 -8 26 248
use FILL  FILL257250x108150
timestamp 0
transform -1 0 17170 0 -1 7450
box -6 -8 26 248
use FILL  FILL257250x111750
timestamp 0
transform 1 0 17150 0 1 7450
box -6 -8 26 248
use FILL  FILL257250x115350
timestamp 0
transform -1 0 17170 0 -1 7930
box -6 -8 26 248
use FILL  FILL257250x122550
timestamp 0
transform -1 0 17170 0 -1 8410
box -6 -8 26 248
use FILL  FILL257250x126150
timestamp 0
transform 1 0 17150 0 1 8410
box -6 -8 26 248
use FILL  FILL257250x129750
timestamp 0
transform -1 0 17170 0 -1 8890
box -6 -8 26 248
use FILL  FILL257250x133350
timestamp 0
transform 1 0 17150 0 1 8890
box -6 -8 26 248
use FILL  FILL257250x136950
timestamp 0
transform -1 0 17170 0 -1 9370
box -6 -8 26 248
use FILL  FILL257250x140550
timestamp 0
transform 1 0 17150 0 1 9370
box -6 -8 26 248
use FILL  FILL257250x144150
timestamp 0
transform -1 0 17170 0 -1 9850
box -6 -8 26 248
use FILL  FILL257250x147750
timestamp 0
transform 1 0 17150 0 1 9850
box -6 -8 26 248
use FILL  FILL257250x158550
timestamp 0
transform -1 0 17170 0 -1 10810
box -6 -8 26 248
use FILL  FILL257250x165750
timestamp 0
transform -1 0 17170 0 -1 11290
box -6 -8 26 248
use FILL  FILL257250x169350
timestamp 0
transform 1 0 17150 0 1 11290
box -6 -8 26 248
use FILL  FILL257250x176550
timestamp 0
transform 1 0 17150 0 1 11770
box -6 -8 26 248
use FILL  FILL257250x180150
timestamp 0
transform -1 0 17170 0 -1 12250
box -6 -8 26 248
use FILL  FILL257250x183750
timestamp 0
transform 1 0 17150 0 1 12250
box -6 -8 26 248
use FILL  FILL257250x187350
timestamp 0
transform -1 0 17170 0 -1 12730
box -6 -8 26 248
use FILL  FILL257250x190950
timestamp 0
transform 1 0 17150 0 1 12730
box -6 -8 26 248
use FILL  FILL257250x198150
timestamp 0
transform 1 0 17150 0 1 13210
box -6 -8 26 248
use FILL  FILL257250x201750
timestamp 0
transform -1 0 17170 0 -1 13690
box -6 -8 26 248
use FILL  FILL257250x208950
timestamp 0
transform -1 0 17170 0 -1 14170
box -6 -8 26 248
use FILL  FILL257250x212550
timestamp 0
transform 1 0 17150 0 1 14170
box -6 -8 26 248
use FILL  FILL257250x216150
timestamp 0
transform -1 0 17170 0 -1 14650
box -6 -8 26 248
use FILL  FILL257250x219750
timestamp 0
transform 1 0 17150 0 1 14650
box -6 -8 26 248
use FILL  FILL257250x223350
timestamp 0
transform -1 0 17170 0 -1 15130
box -6 -8 26 248
use FILL  FILL257250x226950
timestamp 0
transform 1 0 17150 0 1 15130
box -6 -8 26 248
use FILL  FILL257250x230550
timestamp 0
transform -1 0 17170 0 -1 15610
box -6 -8 26 248
use FILL  FILL257250x234150
timestamp 0
transform 1 0 17150 0 1 15610
box -6 -8 26 248
use FILL  FILL257250x237750
timestamp 0
transform -1 0 17170 0 -1 16090
box -6 -8 26 248
use FILL  FILL257250x241350
timestamp 0
transform 1 0 17150 0 1 16090
box -6 -8 26 248
use FILL  FILL257250x244950
timestamp 0
transform -1 0 17170 0 -1 16570
box -6 -8 26 248
use FILL  FILL257250x248550
timestamp 0
transform 1 0 17150 0 1 16570
box -6 -8 26 248
use FILL  FILL257250x252150
timestamp 0
transform -1 0 17170 0 -1 17050
box -6 -8 26 248
use FILL  FILL257550x150
timestamp 0
transform -1 0 17190 0 -1 250
box -6 -8 26 248
use FILL  FILL257550x3750
timestamp 0
transform 1 0 17170 0 1 250
box -6 -8 26 248
use FILL  FILL257550x7350
timestamp 0
transform -1 0 17190 0 -1 730
box -6 -8 26 248
use FILL  FILL257550x10950
timestamp 0
transform 1 0 17170 0 1 730
box -6 -8 26 248
use FILL  FILL257550x14550
timestamp 0
transform -1 0 17190 0 -1 1210
box -6 -8 26 248
use FILL  FILL257550x18150
timestamp 0
transform 1 0 17170 0 1 1210
box -6 -8 26 248
use FILL  FILL257550x21750
timestamp 0
transform -1 0 17190 0 -1 1690
box -6 -8 26 248
use FILL  FILL257550x25350
timestamp 0
transform 1 0 17170 0 1 1690
box -6 -8 26 248
use FILL  FILL257550x28950
timestamp 0
transform -1 0 17190 0 -1 2170
box -6 -8 26 248
use FILL  FILL257550x32550
timestamp 0
transform 1 0 17170 0 1 2170
box -6 -8 26 248
use FILL  FILL257550x36150
timestamp 0
transform -1 0 17190 0 -1 2650
box -6 -8 26 248
use FILL  FILL257550x39750
timestamp 0
transform 1 0 17170 0 1 2650
box -6 -8 26 248
use FILL  FILL257550x43350
timestamp 0
transform -1 0 17190 0 -1 3130
box -6 -8 26 248
use FILL  FILL257550x46950
timestamp 0
transform 1 0 17170 0 1 3130
box -6 -8 26 248
use FILL  FILL257550x50550
timestamp 0
transform -1 0 17190 0 -1 3610
box -6 -8 26 248
use FILL  FILL257550x54150
timestamp 0
transform 1 0 17170 0 1 3610
box -6 -8 26 248
use FILL  FILL257550x57750
timestamp 0
transform -1 0 17190 0 -1 4090
box -6 -8 26 248
use FILL  FILL257550x61350
timestamp 0
transform 1 0 17170 0 1 4090
box -6 -8 26 248
use FILL  FILL257550x64950
timestamp 0
transform -1 0 17190 0 -1 4570
box -6 -8 26 248
use FILL  FILL257550x68550
timestamp 0
transform 1 0 17170 0 1 4570
box -6 -8 26 248
use FILL  FILL257550x72150
timestamp 0
transform -1 0 17190 0 -1 5050
box -6 -8 26 248
use FILL  FILL257550x75750
timestamp 0
transform 1 0 17170 0 1 5050
box -6 -8 26 248
use FILL  FILL257550x79350
timestamp 0
transform -1 0 17190 0 -1 5530
box -6 -8 26 248
use FILL  FILL257550x82950
timestamp 0
transform 1 0 17170 0 1 5530
box -6 -8 26 248
use FILL  FILL257550x86550
timestamp 0
transform -1 0 17190 0 -1 6010
box -6 -8 26 248
use FILL  FILL257550x90150
timestamp 0
transform 1 0 17170 0 1 6010
box -6 -8 26 248
use FILL  FILL257550x93750
timestamp 0
transform -1 0 17190 0 -1 6490
box -6 -8 26 248
use FILL  FILL257550x97350
timestamp 0
transform 1 0 17170 0 1 6490
box -6 -8 26 248
use FILL  FILL257550x100950
timestamp 0
transform -1 0 17190 0 -1 6970
box -6 -8 26 248
use FILL  FILL257550x104550
timestamp 0
transform 1 0 17170 0 1 6970
box -6 -8 26 248
use FILL  FILL257550x108150
timestamp 0
transform -1 0 17190 0 -1 7450
box -6 -8 26 248
use FILL  FILL257550x111750
timestamp 0
transform 1 0 17170 0 1 7450
box -6 -8 26 248
use FILL  FILL257550x115350
timestamp 0
transform -1 0 17190 0 -1 7930
box -6 -8 26 248
use FILL  FILL257550x118950
timestamp 0
transform 1 0 17170 0 1 7930
box -6 -8 26 248
use FILL  FILL257550x122550
timestamp 0
transform -1 0 17190 0 -1 8410
box -6 -8 26 248
use FILL  FILL257550x126150
timestamp 0
transform 1 0 17170 0 1 8410
box -6 -8 26 248
use FILL  FILL257550x129750
timestamp 0
transform -1 0 17190 0 -1 8890
box -6 -8 26 248
use FILL  FILL257550x133350
timestamp 0
transform 1 0 17170 0 1 8890
box -6 -8 26 248
use FILL  FILL257550x136950
timestamp 0
transform -1 0 17190 0 -1 9370
box -6 -8 26 248
use FILL  FILL257550x140550
timestamp 0
transform 1 0 17170 0 1 9370
box -6 -8 26 248
use FILL  FILL257550x144150
timestamp 0
transform -1 0 17190 0 -1 9850
box -6 -8 26 248
use FILL  FILL257550x147750
timestamp 0
transform 1 0 17170 0 1 9850
box -6 -8 26 248
use FILL  FILL257550x151350
timestamp 0
transform -1 0 17190 0 -1 10330
box -6 -8 26 248
use FILL  FILL257550x154950
timestamp 0
transform 1 0 17170 0 1 10330
box -6 -8 26 248
use FILL  FILL257550x158550
timestamp 0
transform -1 0 17190 0 -1 10810
box -6 -8 26 248
use FILL  FILL257550x165750
timestamp 0
transform -1 0 17190 0 -1 11290
box -6 -8 26 248
use FILL  FILL257550x169350
timestamp 0
transform 1 0 17170 0 1 11290
box -6 -8 26 248
use FILL  FILL257550x172950
timestamp 0
transform -1 0 17190 0 -1 11770
box -6 -8 26 248
use FILL  FILL257550x176550
timestamp 0
transform 1 0 17170 0 1 11770
box -6 -8 26 248
use FILL  FILL257550x180150
timestamp 0
transform -1 0 17190 0 -1 12250
box -6 -8 26 248
use FILL  FILL257550x183750
timestamp 0
transform 1 0 17170 0 1 12250
box -6 -8 26 248
use FILL  FILL257550x187350
timestamp 0
transform -1 0 17190 0 -1 12730
box -6 -8 26 248
use FILL  FILL257550x190950
timestamp 0
transform 1 0 17170 0 1 12730
box -6 -8 26 248
use FILL  FILL257550x194550
timestamp 0
transform -1 0 17190 0 -1 13210
box -6 -8 26 248
use FILL  FILL257550x198150
timestamp 0
transform 1 0 17170 0 1 13210
box -6 -8 26 248
use FILL  FILL257550x201750
timestamp 0
transform -1 0 17190 0 -1 13690
box -6 -8 26 248
use FILL  FILL257550x208950
timestamp 0
transform -1 0 17190 0 -1 14170
box -6 -8 26 248
use FILL  FILL257550x212550
timestamp 0
transform 1 0 17170 0 1 14170
box -6 -8 26 248
use FILL  FILL257550x216150
timestamp 0
transform -1 0 17190 0 -1 14650
box -6 -8 26 248
use FILL  FILL257550x219750
timestamp 0
transform 1 0 17170 0 1 14650
box -6 -8 26 248
use FILL  FILL257550x223350
timestamp 0
transform -1 0 17190 0 -1 15130
box -6 -8 26 248
use FILL  FILL257550x226950
timestamp 0
transform 1 0 17170 0 1 15130
box -6 -8 26 248
use FILL  FILL257550x230550
timestamp 0
transform -1 0 17190 0 -1 15610
box -6 -8 26 248
use FILL  FILL257550x234150
timestamp 0
transform 1 0 17170 0 1 15610
box -6 -8 26 248
use FILL  FILL257550x237750
timestamp 0
transform -1 0 17190 0 -1 16090
box -6 -8 26 248
use FILL  FILL257550x241350
timestamp 0
transform 1 0 17170 0 1 16090
box -6 -8 26 248
use FILL  FILL257550x244950
timestamp 0
transform -1 0 17190 0 -1 16570
box -6 -8 26 248
use FILL  FILL257550x248550
timestamp 0
transform 1 0 17170 0 1 16570
box -6 -8 26 248
use FILL  FILL257550x252150
timestamp 0
transform -1 0 17190 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__7072_
timestamp 0
transform 1 0 6130 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__7073_
timestamp 0
transform 1 0 8790 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7074_
timestamp 0
transform 1 0 6670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7075_
timestamp 0
transform 1 0 7630 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__7076_
timestamp 0
transform -1 0 5810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7077_
timestamp 0
transform -1 0 8590 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7078_
timestamp 0
transform -1 0 5450 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7079_
timestamp 0
transform -1 0 6770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7080_
timestamp 0
transform -1 0 8590 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7081_
timestamp 0
transform -1 0 5390 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7082_
timestamp 0
transform -1 0 6370 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7083_
timestamp 0
transform 1 0 5930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7084_
timestamp 0
transform 1 0 8650 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7085_
timestamp 0
transform 1 0 5810 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7086_
timestamp 0
transform -1 0 5590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7087_
timestamp 0
transform -1 0 5470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7088_
timestamp 0
transform -1 0 5170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7089_
timestamp 0
transform -1 0 5330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7090_
timestamp 0
transform -1 0 7850 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7091_
timestamp 0
transform -1 0 5410 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7092_
timestamp 0
transform -1 0 5550 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7093_
timestamp 0
transform -1 0 5230 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7094_
timestamp 0
transform 1 0 5290 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7095_
timestamp 0
transform -1 0 5190 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7096_
timestamp 0
transform -1 0 5670 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7097_
timestamp 0
transform -1 0 5790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7098_
timestamp 0
transform -1 0 5790 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7099_
timestamp 0
transform 1 0 5610 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7100_
timestamp 0
transform 1 0 5430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7101_
timestamp 0
transform 1 0 5350 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__7102_
timestamp 0
transform -1 0 5230 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__7103_
timestamp 0
transform 1 0 6370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7104_
timestamp 0
transform 1 0 5090 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__7105_
timestamp 0
transform 1 0 5310 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7106_
timestamp 0
transform 1 0 4950 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__7107_
timestamp 0
transform 1 0 4870 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7108_
timestamp 0
transform 1 0 5930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7109_
timestamp 0
transform 1 0 5190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7110_
timestamp 0
transform -1 0 5330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7111_
timestamp 0
transform 1 0 5470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7112_
timestamp 0
transform -1 0 6210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7113_
timestamp 0
transform -1 0 5570 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7114_
timestamp 0
transform -1 0 10350 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7115_
timestamp 0
transform -1 0 8950 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__7116_
timestamp 0
transform -1 0 8810 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__7117_
timestamp 0
transform -1 0 10770 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7118_
timestamp 0
transform -1 0 8990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7119_
timestamp 0
transform 1 0 8630 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__7120_
timestamp 0
transform -1 0 8010 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__7121_
timestamp 0
transform -1 0 8070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7122_
timestamp 0
transform -1 0 7870 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__7123_
timestamp 0
transform -1 0 9430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7124_
timestamp 0
transform 1 0 9090 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__7125_
timestamp 0
transform -1 0 9230 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7126_
timestamp 0
transform 1 0 9230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7127_
timestamp 0
transform 1 0 9070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7128_
timestamp 0
transform 1 0 8750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7129_
timestamp 0
transform -1 0 8930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7130_
timestamp 0
transform 1 0 7430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7131_
timestamp 0
transform 1 0 8450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7132_
timestamp 0
transform 1 0 8430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7133_
timestamp 0
transform 1 0 7370 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7134_
timestamp 0
transform 1 0 13030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7135_
timestamp 0
transform 1 0 13250 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7136_
timestamp 0
transform 1 0 13090 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7137_
timestamp 0
transform 1 0 11990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7138_
timestamp 0
transform -1 0 10450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7139_
timestamp 0
transform -1 0 10830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7140_
timestamp 0
transform 1 0 10750 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7141_
timestamp 0
transform -1 0 9270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7142_
timestamp 0
transform -1 0 8990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7143_
timestamp 0
transform -1 0 9110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7144_
timestamp 0
transform -1 0 9250 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7145_
timestamp 0
transform 1 0 9690 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7146_
timestamp 0
transform 1 0 9530 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7147_
timestamp 0
transform 1 0 9510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7148_
timestamp 0
transform -1 0 9970 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7149_
timestamp 0
transform 1 0 8330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7150_
timestamp 0
transform 1 0 8870 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7151_
timestamp 0
transform -1 0 7850 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7152_
timestamp 0
transform -1 0 9730 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7153_
timestamp 0
transform 1 0 9710 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7154_
timestamp 0
transform 1 0 10990 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7155_
timestamp 0
transform 1 0 7930 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7156_
timestamp 0
transform 1 0 7530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7157_
timestamp 0
transform -1 0 6470 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7158_
timestamp 0
transform -1 0 6450 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7159_
timestamp 0
transform 1 0 9310 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7160_
timestamp 0
transform -1 0 10150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7161_
timestamp 0
transform -1 0 9990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7162_
timestamp 0
transform 1 0 9170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7163_
timestamp 0
transform 1 0 7950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7164_
timestamp 0
transform -1 0 8590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7165_
timestamp 0
transform 1 0 8630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7166_
timestamp 0
transform 1 0 8810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7167_
timestamp 0
transform -1 0 9170 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7168_
timestamp 0
transform -1 0 9030 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7169_
timestamp 0
transform 1 0 8790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7170_
timestamp 0
transform -1 0 7590 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7171_
timestamp 0
transform -1 0 8610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7172_
timestamp 0
transform 1 0 11110 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7173_
timestamp 0
transform -1 0 9730 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7174_
timestamp 0
transform -1 0 9850 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7175_
timestamp 0
transform 1 0 8290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7176_
timestamp 0
transform 1 0 8470 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7177_
timestamp 0
transform 1 0 8310 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7178_
timestamp 0
transform -1 0 8350 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7179_
timestamp 0
transform 1 0 10310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7180_
timestamp 0
transform 1 0 9270 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7181_
timestamp 0
transform 1 0 9110 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7182_
timestamp 0
transform 1 0 9430 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7183_
timestamp 0
transform 1 0 8830 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7184_
timestamp 0
transform -1 0 8970 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7185_
timestamp 0
transform 1 0 8670 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7186_
timestamp 0
transform 1 0 8490 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7187_
timestamp 0
transform -1 0 8370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7188_
timestamp 0
transform -1 0 7970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7189_
timestamp 0
transform -1 0 8150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7190_
timestamp 0
transform 1 0 7790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7191_
timestamp 0
transform 1 0 10310 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7192_
timestamp 0
transform 1 0 9790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7193_
timestamp 0
transform -1 0 10150 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7194_
timestamp 0
transform 1 0 9550 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7195_
timestamp 0
transform 1 0 8490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7196_
timestamp 0
transform -1 0 7930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7197_
timestamp 0
transform 1 0 8070 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7198_
timestamp 0
transform 1 0 8070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7199_
timestamp 0
transform 1 0 8170 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7200_
timestamp 0
transform 1 0 8430 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7201_
timestamp 0
transform 1 0 8730 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7202_
timestamp 0
transform -1 0 8610 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7203_
timestamp 0
transform -1 0 6590 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7204_
timestamp 0
transform 1 0 7730 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__7205_
timestamp 0
transform 1 0 9370 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7206_
timestamp 0
transform 1 0 7930 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__7207_
timestamp 0
transform -1 0 6330 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7208_
timestamp 0
transform -1 0 7770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7209_
timestamp 0
transform -1 0 9830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7210_
timestamp 0
transform -1 0 8870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7211_
timestamp 0
transform -1 0 9670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7212_
timestamp 0
transform -1 0 9370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7213_
timestamp 0
transform 1 0 9490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7214_
timestamp 0
transform 1 0 9030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7215_
timestamp 0
transform 1 0 8870 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7216_
timestamp 0
transform 1 0 9030 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7217_
timestamp 0
transform 1 0 9150 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7218_
timestamp 0
transform 1 0 9410 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7219_
timestamp 0
transform 1 0 9270 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7220_
timestamp 0
transform -1 0 8610 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7221_
timestamp 0
transform 1 0 8730 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7222_
timestamp 0
transform -1 0 8330 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7223_
timestamp 0
transform -1 0 7810 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7224_
timestamp 0
transform -1 0 7670 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7225_
timestamp 0
transform -1 0 7570 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7226_
timestamp 0
transform 1 0 7930 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7227_
timestamp 0
transform -1 0 7410 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7228_
timestamp 0
transform -1 0 7710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7229_
timestamp 0
transform -1 0 6110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7230_
timestamp 0
transform 1 0 6350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7231_
timestamp 0
transform -1 0 5890 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7232_
timestamp 0
transform 1 0 6250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7233_
timestamp 0
transform 1 0 8450 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7234_
timestamp 0
transform 1 0 8330 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7235_
timestamp 0
transform -1 0 6930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7236_
timestamp 0
transform -1 0 8710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7237_
timestamp 0
transform 1 0 11230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7238_
timestamp 0
transform -1 0 9310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7239_
timestamp 0
transform -1 0 9430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7240_
timestamp 0
transform 1 0 7770 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7241_
timestamp 0
transform 1 0 7610 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7242_
timestamp 0
transform 1 0 7950 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7243_
timestamp 0
transform -1 0 8070 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7244_
timestamp 0
transform -1 0 8170 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7245_
timestamp 0
transform 1 0 7290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7246_
timestamp 0
transform -1 0 6450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7247_
timestamp 0
transform 1 0 6350 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7248_
timestamp 0
transform 1 0 6490 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7249_
timestamp 0
transform 1 0 6350 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7250_
timestamp 0
transform -1 0 6150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7251_
timestamp 0
transform -1 0 6310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7252_
timestamp 0
transform 1 0 6390 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7253_
timestamp 0
transform 1 0 6390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7254_
timestamp 0
transform 1 0 8190 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7255_
timestamp 0
transform -1 0 8050 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7256_
timestamp 0
transform 1 0 6250 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7257_
timestamp 0
transform -1 0 6270 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7258_
timestamp 0
transform -1 0 5750 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7259_
timestamp 0
transform -1 0 9810 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7260_
timestamp 0
transform -1 0 7910 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7261_
timestamp 0
transform -1 0 8030 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7262_
timestamp 0
transform -1 0 8210 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7263_
timestamp 0
transform 1 0 7550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7264_
timestamp 0
transform -1 0 7950 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7265_
timestamp 0
transform -1 0 6650 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7266_
timestamp 0
transform -1 0 6470 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7267_
timestamp 0
transform -1 0 5650 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7268_
timestamp 0
transform -1 0 5010 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7269_
timestamp 0
transform 1 0 5790 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7270_
timestamp 0
transform -1 0 5150 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7271_
timestamp 0
transform 1 0 4850 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7272_
timestamp 0
transform -1 0 5450 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7273_
timestamp 0
transform 1 0 5290 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7274_
timestamp 0
transform 1 0 5570 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7275_
timestamp 0
transform -1 0 5610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7276_
timestamp 0
transform -1 0 5970 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7277_
timestamp 0
transform 1 0 5790 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7278_
timestamp 0
transform 1 0 5710 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7279_
timestamp 0
transform 1 0 6090 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7280_
timestamp 0
transform 1 0 6550 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7281_
timestamp 0
transform -1 0 6210 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7282_
timestamp 0
transform -1 0 7390 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7283_
timestamp 0
transform 1 0 7430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7284_
timestamp 0
transform -1 0 7330 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7285_
timestamp 0
transform 1 0 6790 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7286_
timestamp 0
transform 1 0 6750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7287_
timestamp 0
transform -1 0 6070 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7288_
timestamp 0
transform -1 0 6570 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7289_
timestamp 0
transform -1 0 5530 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7290_
timestamp 0
transform -1 0 5630 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7291_
timestamp 0
transform -1 0 5770 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7292_
timestamp 0
transform 1 0 5910 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7293_
timestamp 0
transform 1 0 5930 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7294_
timestamp 0
transform 1 0 6010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7295_
timestamp 0
transform -1 0 7790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7296_
timestamp 0
transform 1 0 7870 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7297_
timestamp 0
transform -1 0 7270 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7298_
timestamp 0
transform 1 0 6030 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7299_
timestamp 0
transform 1 0 5370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7300_
timestamp 0
transform -1 0 4250 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7301_
timestamp 0
transform -1 0 5110 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7302_
timestamp 0
transform -1 0 7490 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7303_
timestamp 0
transform 1 0 7050 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7304_
timestamp 0
transform 1 0 6910 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7305_
timestamp 0
transform -1 0 4790 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7306_
timestamp 0
transform -1 0 4370 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7307_
timestamp 0
transform -1 0 5390 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7308_
timestamp 0
transform -1 0 4110 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7309_
timestamp 0
transform 1 0 3950 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7310_
timestamp 0
transform -1 0 4630 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7311_
timestamp 0
transform -1 0 4470 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7312_
timestamp 0
transform -1 0 4470 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7313_
timestamp 0
transform -1 0 4610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7314_
timestamp 0
transform -1 0 4730 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7315_
timestamp 0
transform 1 0 5470 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7316_
timestamp 0
transform -1 0 5470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7317_
timestamp 0
transform -1 0 5330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7318_
timestamp 0
transform 1 0 5650 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7319_
timestamp 0
transform 1 0 5510 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7320_
timestamp 0
transform 1 0 5470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7321_
timestamp 0
transform 1 0 5190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7322_
timestamp 0
transform -1 0 3810 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7323_
timestamp 0
transform 1 0 5790 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7324_
timestamp 0
transform -1 0 5870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7325_
timestamp 0
transform 1 0 5650 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7326_
timestamp 0
transform -1 0 5730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7327_
timestamp 0
transform -1 0 4730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7328_
timestamp 0
transform -1 0 6630 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7329_
timestamp 0
transform 1 0 5150 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7330_
timestamp 0
transform -1 0 7330 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7331_
timestamp 0
transform -1 0 7250 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7332_
timestamp 0
transform -1 0 7150 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7333_
timestamp 0
transform -1 0 7030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7334_
timestamp 0
transform -1 0 6210 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7335_
timestamp 0
transform -1 0 5070 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7336_
timestamp 0
transform -1 0 4950 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7337_
timestamp 0
transform -1 0 4950 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7338_
timestamp 0
transform -1 0 6070 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7339_
timestamp 0
transform 1 0 5310 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7340_
timestamp 0
transform 1 0 5530 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7341_
timestamp 0
transform 1 0 5370 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7342_
timestamp 0
transform 1 0 5250 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7343_
timestamp 0
transform -1 0 4990 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7344_
timestamp 0
transform -1 0 4870 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7345_
timestamp 0
transform -1 0 5050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7346_
timestamp 0
transform 1 0 5110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7347_
timestamp 0
transform -1 0 5250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7348_
timestamp 0
transform 1 0 5290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7349_
timestamp 0
transform 1 0 5250 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7350_
timestamp 0
transform 1 0 5290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7351_
timestamp 0
transform 1 0 6130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7352_
timestamp 0
transform 1 0 5170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7353_
timestamp 0
transform -1 0 5250 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7354_
timestamp 0
transform 1 0 5370 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7355_
timestamp 0
transform -1 0 5410 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7356_
timestamp 0
transform 1 0 5910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7357_
timestamp 0
transform -1 0 6650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7358_
timestamp 0
transform -1 0 5810 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7359_
timestamp 0
transform -1 0 5530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7360_
timestamp 0
transform -1 0 5690 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7361_
timestamp 0
transform -1 0 5650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7362_
timestamp 0
transform 1 0 5510 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7363_
timestamp 0
transform 1 0 5950 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7364_
timestamp 0
transform 1 0 5770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7365_
timestamp 0
transform 1 0 6090 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7366_
timestamp 0
transform 1 0 6790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7367_
timestamp 0
transform -1 0 6810 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7368_
timestamp 0
transform -1 0 6290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7369_
timestamp 0
transform -1 0 6150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7370_
timestamp 0
transform -1 0 5970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7371_
timestamp 0
transform 1 0 4970 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7372_
timestamp 0
transform -1 0 4890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7373_
timestamp 0
transform 1 0 4790 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7374_
timestamp 0
transform 1 0 5090 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7375_
timestamp 0
transform -1 0 5110 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7376_
timestamp 0
transform 1 0 6930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7377_
timestamp 0
transform -1 0 6650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7378_
timestamp 0
transform 1 0 7910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7379_
timestamp 0
transform 1 0 6050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7380_
timestamp 0
transform -1 0 6310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7381_
timestamp 0
transform 1 0 6490 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7382_
timestamp 0
transform 1 0 6410 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7383_
timestamp 0
transform 1 0 6530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7384_
timestamp 0
transform 1 0 6570 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7385_
timestamp 0
transform -1 0 7490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7386_
timestamp 0
transform 1 0 6250 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7387_
timestamp 0
transform -1 0 6790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7388_
timestamp 0
transform -1 0 7050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7389_
timestamp 0
transform -1 0 7190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7390_
timestamp 0
transform -1 0 6430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7391_
timestamp 0
transform -1 0 6470 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7392_
timestamp 0
transform -1 0 6330 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7393_
timestamp 0
transform -1 0 5050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7394_
timestamp 0
transform 1 0 7270 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7395_
timestamp 0
transform -1 0 7050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7396_
timestamp 0
transform -1 0 7050 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7397_
timestamp 0
transform 1 0 6890 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7398_
timestamp 0
transform 1 0 6730 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7399_
timestamp 0
transform 1 0 8290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7400_
timestamp 0
transform -1 0 7170 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7401_
timestamp 0
transform -1 0 7290 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7402_
timestamp 0
transform 1 0 7190 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7403_
timestamp 0
transform 1 0 7550 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7404_
timestamp 0
transform 1 0 8410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7405_
timestamp 0
transform 1 0 8150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7406_
timestamp 0
transform 1 0 8010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7407_
timestamp 0
transform 1 0 7750 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7408_
timestamp 0
transform 1 0 7610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7409_
timestamp 0
transform 1 0 7330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7410_
timestamp 0
transform 1 0 7170 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7411_
timestamp 0
transform 1 0 7610 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7412_
timestamp 0
transform 1 0 6930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7413_
timestamp 0
transform 1 0 7330 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7414_
timestamp 0
transform 1 0 7470 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7415_
timestamp 0
transform 1 0 7090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7416_
timestamp 0
transform -1 0 7130 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7417_
timestamp 0
transform 1 0 5910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7418_
timestamp 0
transform -1 0 5430 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7419_
timestamp 0
transform -1 0 6850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7420_
timestamp 0
transform 1 0 7410 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7421_
timestamp 0
transform 1 0 7010 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7422_
timestamp 0
transform 1 0 7630 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7423_
timestamp 0
transform 1 0 7550 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7424_
timestamp 0
transform -1 0 7650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7425_
timestamp 0
transform 1 0 7390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7426_
timestamp 0
transform -1 0 7530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7427_
timestamp 0
transform -1 0 7270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7428_
timestamp 0
transform 1 0 7010 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7429_
timestamp 0
transform -1 0 6790 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7430_
timestamp 0
transform -1 0 6710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7431_
timestamp 0
transform -1 0 6570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7432_
timestamp 0
transform -1 0 6630 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7433_
timestamp 0
transform 1 0 5570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7434_
timestamp 0
transform 1 0 8190 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7435_
timestamp 0
transform 1 0 7450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7436_
timestamp 0
transform -1 0 7190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7437_
timestamp 0
transform -1 0 7330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7438_
timestamp 0
transform -1 0 7550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7439_
timestamp 0
transform 1 0 8010 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7440_
timestamp 0
transform 1 0 7150 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7441_
timestamp 0
transform -1 0 7690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7442_
timestamp 0
transform 1 0 7650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7443_
timestamp 0
transform 1 0 5230 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7444_
timestamp 0
transform -1 0 4590 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7445_
timestamp 0
transform 1 0 6510 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7446_
timestamp 0
transform 1 0 6350 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7447_
timestamp 0
transform -1 0 7670 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7448_
timestamp 0
transform 1 0 8210 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7449_
timestamp 0
transform 1 0 8750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7450_
timestamp 0
transform -1 0 8710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7451_
timestamp 0
transform -1 0 8050 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7452_
timestamp 0
transform -1 0 7550 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7453_
timestamp 0
transform 1 0 8170 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7454_
timestamp 0
transform 1 0 8290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7455_
timestamp 0
transform -1 0 10030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7456_
timestamp 0
transform -1 0 8590 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7457_
timestamp 0
transform -1 0 8490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7458_
timestamp 0
transform 1 0 10330 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7459_
timestamp 0
transform -1 0 5930 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7460_
timestamp 0
transform -1 0 6610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7461_
timestamp 0
transform -1 0 7690 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7462_
timestamp 0
transform -1 0 7810 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7463_
timestamp 0
transform 1 0 8030 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7464_
timestamp 0
transform 1 0 8390 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7465_
timestamp 0
transform 1 0 6850 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7466_
timestamp 0
transform 1 0 6710 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7467_
timestamp 0
transform 1 0 8470 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7468_
timestamp 0
transform -1 0 6790 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7469_
timestamp 0
transform -1 0 6910 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7470_
timestamp 0
transform -1 0 8210 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7471_
timestamp 0
transform 1 0 8330 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7472_
timestamp 0
transform -1 0 8690 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7473_
timestamp 0
transform -1 0 9170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7474_
timestamp 0
transform -1 0 8230 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7475_
timestamp 0
transform 1 0 8510 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7476_
timestamp 0
transform -1 0 9030 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7477_
timestamp 0
transform 1 0 9550 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7478_
timestamp 0
transform -1 0 11070 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7479_
timestamp 0
transform 1 0 9390 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7480_
timestamp 0
transform -1 0 10930 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7481_
timestamp 0
transform -1 0 10130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7482_
timestamp 0
transform -1 0 9970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7483_
timestamp 0
transform -1 0 9390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7484_
timestamp 0
transform -1 0 8610 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7485_
timestamp 0
transform -1 0 8730 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7486_
timestamp 0
transform 1 0 11150 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7487_
timestamp 0
transform -1 0 9250 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7488_
timestamp 0
transform -1 0 7630 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7489_
timestamp 0
transform -1 0 7750 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7490_
timestamp 0
transform -1 0 7830 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7491_
timestamp 0
transform 1 0 8310 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7492_
timestamp 0
transform 1 0 7790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7493_
timestamp 0
transform 1 0 7910 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7494_
timestamp 0
transform -1 0 7790 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7495_
timestamp 0
transform 1 0 8610 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7496_
timestamp 0
transform -1 0 9050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7497_
timestamp 0
transform 1 0 9490 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7498_
timestamp 0
transform 1 0 8830 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7499_
timestamp 0
transform -1 0 8910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7500_
timestamp 0
transform 1 0 10130 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7501_
timestamp 0
transform -1 0 11630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7502_
timestamp 0
transform 1 0 9990 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7503_
timestamp 0
transform 1 0 11590 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7504_
timestamp 0
transform -1 0 11330 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7505_
timestamp 0
transform 1 0 11450 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7506_
timestamp 0
transform -1 0 10910 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7507_
timestamp 0
transform -1 0 8850 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7508_
timestamp 0
transform 1 0 11730 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7509_
timestamp 0
transform 1 0 12190 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7510_
timestamp 0
transform -1 0 7690 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7511_
timestamp 0
transform -1 0 7830 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7512_
timestamp 0
transform 1 0 8590 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7513_
timestamp 0
transform 1 0 9010 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7514_
timestamp 0
transform -1 0 8070 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7515_
timestamp 0
transform -1 0 7930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7516_
timestamp 0
transform -1 0 8190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7517_
timestamp 0
transform 1 0 9150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7518_
timestamp 0
transform -1 0 9370 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7519_
timestamp 0
transform 1 0 10130 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7520_
timestamp 0
transform 1 0 9310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7521_
timestamp 0
transform 1 0 11330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7522_
timestamp 0
transform 1 0 12090 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7523_
timestamp 0
transform 1 0 11470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7524_
timestamp 0
transform 1 0 12210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7525_
timestamp 0
transform 1 0 12410 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7526_
timestamp 0
transform -1 0 12310 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7527_
timestamp 0
transform 1 0 12550 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7528_
timestamp 0
transform 1 0 9750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7529_
timestamp 0
transform -1 0 11910 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7530_
timestamp 0
transform -1 0 7390 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7531_
timestamp 0
transform -1 0 7510 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7532_
timestamp 0
transform -1 0 7950 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7533_
timestamp 0
transform -1 0 8090 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7534_
timestamp 0
transform 1 0 8730 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7535_
timestamp 0
transform 1 0 8590 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7536_
timestamp 0
transform -1 0 10770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7537_
timestamp 0
transform 1 0 9090 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7538_
timestamp 0
transform 1 0 10790 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7539_
timestamp 0
transform 1 0 11650 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7540_
timestamp 0
transform -1 0 10690 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7541_
timestamp 0
transform -1 0 11130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7542_
timestamp 0
transform 1 0 11810 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7543_
timestamp 0
transform 1 0 11430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7544_
timestamp 0
transform 1 0 11270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7545_
timestamp 0
transform 1 0 12890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7546_
timestamp 0
transform 1 0 12610 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7547_
timestamp 0
transform -1 0 12490 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7548_
timestamp 0
transform 1 0 12610 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7549_
timestamp 0
transform -1 0 12450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7550_
timestamp 0
transform 1 0 11110 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7551_
timestamp 0
transform -1 0 9670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7552_
timestamp 0
transform -1 0 11850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7553_
timestamp 0
transform 1 0 11070 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7554_
timestamp 0
transform -1 0 8370 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7555_
timestamp 0
transform 1 0 8750 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7556_
timestamp 0
transform -1 0 8770 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7557_
timestamp 0
transform -1 0 8890 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7558_
timestamp 0
transform 1 0 10390 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7559_
timestamp 0
transform 1 0 10930 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7560_
timestamp 0
transform 1 0 9250 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7561_
timestamp 0
transform 1 0 9110 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7562_
timestamp 0
transform 1 0 10110 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7563_
timestamp 0
transform -1 0 10270 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7564_
timestamp 0
transform 1 0 10970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7565_
timestamp 0
transform 1 0 13670 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7566_
timestamp 0
transform 1 0 10830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7567_
timestamp 0
transform 1 0 13530 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7568_
timestamp 0
transform -1 0 11710 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7569_
timestamp 0
transform -1 0 11730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7570_
timestamp 0
transform -1 0 11550 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7571_
timestamp 0
transform 1 0 10010 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7572_
timestamp 0
transform 1 0 9090 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7573_
timestamp 0
transform -1 0 10510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7574_
timestamp 0
transform 1 0 8910 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7575_
timestamp 0
transform 1 0 9450 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7576_
timestamp 0
transform 1 0 9590 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7577_
timestamp 0
transform 1 0 10330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7578_
timestamp 0
transform 1 0 9490 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7579_
timestamp 0
transform -1 0 9610 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7580_
timestamp 0
transform 1 0 9750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7581_
timestamp 0
transform 1 0 12490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7582_
timestamp 0
transform -1 0 12970 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7583_
timestamp 0
transform -1 0 12370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7584_
timestamp 0
transform -1 0 11990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7585_
timestamp 0
transform -1 0 12770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7586_
timestamp 0
transform -1 0 12630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7587_
timestamp 0
transform 1 0 12230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7588_
timestamp 0
transform -1 0 12130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7589_
timestamp 0
transform 1 0 12050 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7590_
timestamp 0
transform -1 0 11710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7591_
timestamp 0
transform 1 0 13930 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7592_
timestamp 0
transform 1 0 13790 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7593_
timestamp 0
transform 1 0 13390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7594_
timestamp 0
transform 1 0 13370 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7595_
timestamp 0
transform -1 0 11590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7596_
timestamp 0
transform -1 0 10730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7597_
timestamp 0
transform 1 0 10210 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7598_
timestamp 0
transform 1 0 9210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7599_
timestamp 0
transform 1 0 10150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7600_
timestamp 0
transform 1 0 11850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7601_
timestamp 0
transform -1 0 9630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7602_
timestamp 0
transform 1 0 9050 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7603_
timestamp 0
transform 1 0 9170 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7604_
timestamp 0
transform 1 0 9290 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7605_
timestamp 0
transform 1 0 10390 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7606_
timestamp 0
transform 1 0 9990 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7607_
timestamp 0
transform 1 0 10190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7608_
timestamp 0
transform 1 0 10050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7609_
timestamp 0
transform 1 0 10450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7610_
timestamp 0
transform 1 0 9890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7611_
timestamp 0
transform -1 0 10290 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7612_
timestamp 0
transform 1 0 10690 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7613_
timestamp 0
transform 1 0 11370 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7614_
timestamp 0
transform -1 0 10990 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7615_
timestamp 0
transform 1 0 11110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7616_
timestamp 0
transform -1 0 10890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7617_
timestamp 0
transform -1 0 10850 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7618_
timestamp 0
transform 1 0 10670 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7619_
timestamp 0
transform -1 0 12070 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7620_
timestamp 0
transform 1 0 12190 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7621_
timestamp 0
transform 1 0 12330 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7622_
timestamp 0
transform 1 0 11870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7623_
timestamp 0
transform -1 0 9730 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7624_
timestamp 0
transform 1 0 8870 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7625_
timestamp 0
transform 1 0 9290 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7626_
timestamp 0
transform -1 0 10610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7627_
timestamp 0
transform 1 0 10290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7628_
timestamp 0
transform 1 0 10530 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7629_
timestamp 0
transform 1 0 11510 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7630_
timestamp 0
transform 1 0 11730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7631_
timestamp 0
transform 1 0 10150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7632_
timestamp 0
transform 1 0 10690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7633_
timestamp 0
transform 1 0 11230 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7634_
timestamp 0
transform 1 0 11890 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7635_
timestamp 0
transform -1 0 10670 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7636_
timestamp 0
transform -1 0 11770 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7637_
timestamp 0
transform -1 0 11310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7638_
timestamp 0
transform 1 0 10550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7639_
timestamp 0
transform -1 0 10250 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7640_
timestamp 0
transform 1 0 11590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7641_
timestamp 0
transform 1 0 11450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7642_
timestamp 0
transform 1 0 9150 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7643_
timestamp 0
transform 1 0 10030 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7644_
timestamp 0
transform -1 0 10010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7645_
timestamp 0
transform -1 0 10850 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7646_
timestamp 0
transform 1 0 10950 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7647_
timestamp 0
transform 1 0 11030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7648_
timestamp 0
transform 1 0 12810 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7649_
timestamp 0
transform -1 0 12710 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__7650_
timestamp 0
transform 1 0 11170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7651_
timestamp 0
transform -1 0 11010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7652_
timestamp 0
transform 1 0 11150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7653_
timestamp 0
transform -1 0 10390 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7654_
timestamp 0
transform 1 0 10110 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7655_
timestamp 0
transform 1 0 11490 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7656_
timestamp 0
transform -1 0 11610 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7657_
timestamp 0
transform 1 0 11450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7658_
timestamp 0
transform 1 0 11290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7659_
timestamp 0
transform 1 0 11350 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7660_
timestamp 0
transform 1 0 9430 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7661_
timestamp 0
transform -1 0 9410 0 1 730
box -6 -8 26 248
use FILL  FILL_0__7662_
timestamp 0
transform -1 0 9490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__7663_
timestamp 0
transform 1 0 9630 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7664_
timestamp 0
transform -1 0 10290 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7665_
timestamp 0
transform 1 0 10390 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7666_
timestamp 0
transform 1 0 10550 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__7667_
timestamp 0
transform -1 0 9590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7668_
timestamp 0
transform 1 0 9870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7669_
timestamp 0
transform -1 0 9750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7670_
timestamp 0
transform 1 0 10750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7671_
timestamp 0
transform -1 0 10730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7672_
timestamp 0
transform 1 0 10850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7673_
timestamp 0
transform -1 0 10550 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7674_
timestamp 0
transform 1 0 10150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7675_
timestamp 0
transform 1 0 9930 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7676_
timestamp 0
transform 1 0 11250 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7677_
timestamp 0
transform 1 0 11090 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7678_
timestamp 0
transform 1 0 10370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7679_
timestamp 0
transform 1 0 10230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7680_
timestamp 0
transform 1 0 10490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7681_
timestamp 0
transform 1 0 10630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__7682_
timestamp 0
transform -1 0 10570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7683_
timestamp 0
transform -1 0 10430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7684_
timestamp 0
transform -1 0 10090 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7685_
timestamp 0
transform 1 0 6810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7686_
timestamp 0
transform 1 0 6190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7687_
timestamp 0
transform -1 0 6250 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7688_
timestamp 0
transform -1 0 6090 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7689_
timestamp 0
transform -1 0 6110 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7690_
timestamp 0
transform 1 0 5910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7691_
timestamp 0
transform -1 0 5690 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7692_
timestamp 0
transform -1 0 5790 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7693_
timestamp 0
transform 1 0 5130 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__7694_
timestamp 0
transform -1 0 5470 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7695_
timestamp 0
transform 1 0 5050 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7696_
timestamp 0
transform -1 0 6050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7697_
timestamp 0
transform -1 0 6350 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7698_
timestamp 0
transform -1 0 6350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7699_
timestamp 0
transform -1 0 6210 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7700_
timestamp 0
transform -1 0 5890 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7701_
timestamp 0
transform -1 0 5790 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__7702_
timestamp 0
transform -1 0 5750 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7703_
timestamp 0
transform -1 0 5650 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__7704_
timestamp 0
transform -1 0 5410 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__7705_
timestamp 0
transform 1 0 5510 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__7706_
timestamp 0
transform -1 0 5270 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__7707_
timestamp 0
transform -1 0 5010 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__7708_
timestamp 0
transform -1 0 6030 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7709_
timestamp 0
transform -1 0 5950 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__7710_
timestamp 0
transform 1 0 7190 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__7711_
timestamp 0
transform 1 0 7410 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__7712_
timestamp 0
transform 1 0 7250 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__7713_
timestamp 0
transform 1 0 7590 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__7714_
timestamp 0
transform -1 0 7470 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__7715_
timestamp 0
transform 1 0 7310 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__7716_
timestamp 0
transform -1 0 6810 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__7717_
timestamp 0
transform -1 0 6450 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__7718_
timestamp 0
transform -1 0 6770 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__7719_
timestamp 0
transform 1 0 6530 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__7720_
timestamp 0
transform 1 0 6250 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__7721_
timestamp 0
transform -1 0 5770 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__7722_
timestamp 0
transform -1 0 6910 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__7723_
timestamp 0
transform -1 0 6670 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__7724_
timestamp 0
transform -1 0 6670 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7725_
timestamp 0
transform -1 0 7670 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7726_
timestamp 0
transform -1 0 7530 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7727_
timestamp 0
transform 1 0 7030 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__7728_
timestamp 0
transform 1 0 7350 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__7729_
timestamp 0
transform -1 0 6510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7730_
timestamp 0
transform 1 0 6630 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7731_
timestamp 0
transform -1 0 6310 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7732_
timestamp 0
transform -1 0 6330 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__7733_
timestamp 0
transform 1 0 6390 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__7734_
timestamp 0
transform -1 0 6250 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__7735_
timestamp 0
transform 1 0 6110 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__7736_
timestamp 0
transform -1 0 6470 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__7737_
timestamp 0
transform -1 0 8070 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7738_
timestamp 0
transform -1 0 7330 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7739_
timestamp 0
transform 1 0 7150 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7740_
timestamp 0
transform 1 0 6750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7741_
timestamp 0
transform 1 0 7670 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7742_
timestamp 0
transform -1 0 7450 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7743_
timestamp 0
transform 1 0 7550 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7744_
timestamp 0
transform -1 0 6530 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7745_
timestamp 0
transform -1 0 6970 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__7746_
timestamp 0
transform 1 0 7090 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__7747_
timestamp 0
transform -1 0 6830 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__7748_
timestamp 0
transform 1 0 7570 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7749_
timestamp 0
transform -1 0 8110 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7750_
timestamp 0
transform 1 0 8150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7751_
timestamp 0
transform 1 0 8810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7752_
timestamp 0
transform -1 0 8690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7753_
timestamp 0
transform 1 0 8250 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__7754_
timestamp 0
transform -1 0 8130 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7755_
timestamp 0
transform 1 0 8250 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7756_
timestamp 0
transform -1 0 7990 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7757_
timestamp 0
transform -1 0 7730 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7758_
timestamp 0
transform 1 0 7430 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7759_
timestamp 0
transform 1 0 7310 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7760_
timestamp 0
transform 1 0 7130 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7761_
timestamp 0
transform 1 0 7270 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7762_
timestamp 0
transform -1 0 6410 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7763_
timestamp 0
transform -1 0 7470 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7764_
timestamp 0
transform -1 0 7590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7765_
timestamp 0
transform 1 0 7810 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7766_
timestamp 0
transform 1 0 7830 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7767_
timestamp 0
transform 1 0 7690 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7768_
timestamp 0
transform 1 0 7850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7769_
timestamp 0
transform 1 0 7930 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7770_
timestamp 0
transform 1 0 7810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7771_
timestamp 0
transform -1 0 7810 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7772_
timestamp 0
transform -1 0 7690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7773_
timestamp 0
transform 1 0 7590 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7774_
timestamp 0
transform -1 0 7470 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7775_
timestamp 0
transform 1 0 6890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7776_
timestamp 0
transform 1 0 7030 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7777_
timestamp 0
transform 1 0 7310 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7778_
timestamp 0
transform -1 0 7210 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7779_
timestamp 0
transform 1 0 7050 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7780_
timestamp 0
transform -1 0 6930 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7781_
timestamp 0
transform 1 0 5510 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7782_
timestamp 0
transform 1 0 6610 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7783_
timestamp 0
transform 1 0 5110 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7784_
timestamp 0
transform -1 0 4870 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7785_
timestamp 0
transform -1 0 4730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7786_
timestamp 0
transform 1 0 4990 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7787_
timestamp 0
transform -1 0 5130 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7788_
timestamp 0
transform 1 0 5170 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7789_
timestamp 0
transform 1 0 5250 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7790_
timestamp 0
transform 1 0 5610 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7791_
timestamp 0
transform -1 0 6050 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7792_
timestamp 0
transform -1 0 5910 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7793_
timestamp 0
transform 1 0 5730 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7794_
timestamp 0
transform -1 0 8450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7795_
timestamp 0
transform -1 0 6970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7796_
timestamp 0
transform 1 0 7070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7797_
timestamp 0
transform 1 0 7350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7798_
timestamp 0
transform -1 0 7310 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7799_
timestamp 0
transform -1 0 7210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7800_
timestamp 0
transform -1 0 7190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7801_
timestamp 0
transform -1 0 6470 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7802_
timestamp 0
transform 1 0 6750 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7803_
timestamp 0
transform -1 0 6890 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7804_
timestamp 0
transform -1 0 7190 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7805_
timestamp 0
transform -1 0 7050 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__7806_
timestamp 0
transform -1 0 7410 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7807_
timestamp 0
transform -1 0 7730 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7808_
timestamp 0
transform 1 0 8170 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7809_
timestamp 0
transform 1 0 8430 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7810_
timestamp 0
transform -1 0 7030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7811_
timestamp 0
transform -1 0 8010 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7812_
timestamp 0
transform 1 0 8130 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7813_
timestamp 0
transform 1 0 7850 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7814_
timestamp 0
transform -1 0 6530 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7815_
timestamp 0
transform -1 0 6370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7816_
timestamp 0
transform 1 0 6190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7817_
timestamp 0
transform 1 0 5910 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7818_
timestamp 0
transform 1 0 7430 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7819_
timestamp 0
transform -1 0 7730 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7820_
timestamp 0
transform 1 0 7590 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7821_
timestamp 0
transform -1 0 7310 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7822_
timestamp 0
transform 1 0 7030 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7823_
timestamp 0
transform 1 0 6910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7824_
timestamp 0
transform -1 0 6450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7825_
timestamp 0
transform -1 0 6310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7826_
timestamp 0
transform -1 0 6010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7827_
timestamp 0
transform 1 0 6130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7828_
timestamp 0
transform -1 0 5870 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7829_
timestamp 0
transform 1 0 6030 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7830_
timestamp 0
transform 1 0 6290 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7831_
timestamp 0
transform -1 0 6170 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7832_
timestamp 0
transform 1 0 6730 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7833_
timestamp 0
transform 1 0 8350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7834_
timestamp 0
transform 1 0 6870 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__7835_
timestamp 0
transform -1 0 8610 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7836_
timestamp 0
transform -1 0 8730 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__7837_
timestamp 0
transform 1 0 6870 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7838_
timestamp 0
transform -1 0 6910 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7839_
timestamp 0
transform -1 0 10490 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7840_
timestamp 0
transform -1 0 7510 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__7841_
timestamp 0
transform 1 0 9570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7842_
timestamp 0
transform -1 0 9890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7843_
timestamp 0
transform -1 0 8790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7844_
timestamp 0
transform 1 0 9250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7845_
timestamp 0
transform 1 0 9110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7846_
timestamp 0
transform -1 0 6630 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7847_
timestamp 0
transform -1 0 10610 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7848_
timestamp 0
transform 1 0 10710 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7849_
timestamp 0
transform 1 0 9730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7850_
timestamp 0
transform 1 0 9550 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7851_
timestamp 0
transform -1 0 6130 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__7852_
timestamp 0
transform 1 0 11110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7853_
timestamp 0
transform 1 0 10950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__7854_
timestamp 0
transform 1 0 8890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7855_
timestamp 0
transform -1 0 8770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__7856_
timestamp 0
transform 1 0 8890 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7857_
timestamp 0
transform -1 0 9070 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7858_
timestamp 0
transform -1 0 8750 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7859_
timestamp 0
transform -1 0 8610 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7860_
timestamp 0
transform -1 0 8970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7861_
timestamp 0
transform -1 0 9090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7862_
timestamp 0
transform 1 0 10210 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7863_
timestamp 0
transform 1 0 10050 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__7864_
timestamp 0
transform -1 0 7210 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7865_
timestamp 0
transform -1 0 7050 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__7866_
timestamp 0
transform 1 0 7250 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7867_
timestamp 0
transform 1 0 7110 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7868_
timestamp 0
transform -1 0 6770 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7869_
timestamp 0
transform -1 0 6890 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7870_
timestamp 0
transform -1 0 7030 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7871_
timestamp 0
transform -1 0 6950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7872_
timestamp 0
transform -1 0 7910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7873_
timestamp 0
transform 1 0 7510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7874_
timestamp 0
transform 1 0 6470 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7875_
timestamp 0
transform -1 0 6610 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7876_
timestamp 0
transform 1 0 6650 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7877_
timestamp 0
transform -1 0 6790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7878_
timestamp 0
transform -1 0 6250 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7879_
timestamp 0
transform 1 0 6090 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__7880_
timestamp 0
transform -1 0 6050 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7881_
timestamp 0
transform -1 0 6190 0 1 250
box -6 -8 26 248
use FILL  FILL_0__7882_
timestamp 0
transform -1 0 7150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7883_
timestamp 0
transform 1 0 6990 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7884_
timestamp 0
transform -1 0 7190 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7885_
timestamp 0
transform -1 0 7350 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7886_
timestamp 0
transform -1 0 8070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7887_
timestamp 0
transform 1 0 8170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__7888_
timestamp 0
transform -1 0 7310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7889_
timestamp 0
transform -1 0 7430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__7890_
timestamp 0
transform 1 0 7310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7891_
timestamp 0
transform 1 0 7150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__7892_
timestamp 0
transform 1 0 8470 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7893_
timestamp 0
transform 1 0 8330 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__7894_
timestamp 0
transform 1 0 8310 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7895_
timestamp 0
transform 1 0 8030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7896_
timestamp 0
transform -1 0 8190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7897_
timestamp 0
transform -1 0 6930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7898_
timestamp 0
transform 1 0 7890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7899_
timestamp 0
transform 1 0 7490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__7900_
timestamp 0
transform -1 0 7930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7901_
timestamp 0
transform -1 0 8050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7902_
timestamp 0
transform 1 0 5030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7903_
timestamp 0
transform -1 0 4890 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7904_
timestamp 0
transform -1 0 7850 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7905_
timestamp 0
transform -1 0 7970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7906_
timestamp 0
transform 1 0 8810 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7907_
timestamp 0
transform 1 0 8450 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__7908_
timestamp 0
transform -1 0 8270 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7909_
timestamp 0
transform -1 0 7790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__7910_
timestamp 0
transform 1 0 6750 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7911_
timestamp 0
transform -1 0 6910 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__7912_
timestamp 0
transform 1 0 7030 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7913_
timestamp 0
transform 1 0 6750 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7914_
timestamp 0
transform 1 0 6910 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__7915_
timestamp 0
transform 1 0 6130 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__7996_
timestamp 0
transform -1 0 6210 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__7997_
timestamp 0
transform -1 0 5170 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__7998_
timestamp 0
transform -1 0 4910 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__7999_
timestamp 0
transform 1 0 4970 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8000_
timestamp 0
transform 1 0 4310 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8001_
timestamp 0
transform 1 0 4190 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8002_
timestamp 0
transform -1 0 4470 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8003_
timestamp 0
transform -1 0 4630 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8004_
timestamp 0
transform -1 0 4490 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8005_
timestamp 0
transform -1 0 4330 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8006_
timestamp 0
transform -1 0 5270 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8007_
timestamp 0
transform 1 0 4450 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8008_
timestamp 0
transform 1 0 5030 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8009_
timestamp 0
transform 1 0 4290 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8010_
timestamp 0
transform -1 0 3750 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8011_
timestamp 0
transform -1 0 5430 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__8012_
timestamp 0
transform -1 0 3990 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__8013_
timestamp 0
transform -1 0 4150 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__8014_
timestamp 0
transform 1 0 6530 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8015_
timestamp 0
transform -1 0 5010 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8016_
timestamp 0
transform 1 0 4850 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8017_
timestamp 0
transform 1 0 4830 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8018_
timestamp 0
transform -1 0 4870 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8019_
timestamp 0
transform -1 0 4470 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8020_
timestamp 0
transform 1 0 3270 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8021_
timestamp 0
transform 1 0 4350 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8022_
timestamp 0
transform -1 0 4210 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8023_
timestamp 0
transform 1 0 3310 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8024_
timestamp 0
transform 1 0 2950 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8025_
timestamp 0
transform -1 0 3390 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8026_
timestamp 0
transform -1 0 3530 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8027_
timestamp 0
transform -1 0 4210 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8028_
timestamp 0
transform -1 0 3690 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8029_
timestamp 0
transform 1 0 3330 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8030_
timestamp 0
transform 1 0 3770 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8031_
timestamp 0
transform -1 0 3630 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8032_
timestamp 0
transform 1 0 2850 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8033_
timestamp 0
transform 1 0 3090 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8034_
timestamp 0
transform -1 0 3250 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8035_
timestamp 0
transform -1 0 3350 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8036_
timestamp 0
transform -1 0 4330 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8037_
timestamp 0
transform -1 0 3490 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8038_
timestamp 0
transform 1 0 3050 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8039_
timestamp 0
transform 1 0 4070 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8040_
timestamp 0
transform 1 0 3830 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8041_
timestamp 0
transform 1 0 4410 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8042_
timestamp 0
transform 1 0 4650 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8043_
timestamp 0
transform 1 0 4490 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8044_
timestamp 0
transform -1 0 3710 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8045_
timestamp 0
transform 1 0 3890 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8046_
timestamp 0
transform -1 0 3590 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8047_
timestamp 0
transform 1 0 2750 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8048_
timestamp 0
transform -1 0 3530 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8049_
timestamp 0
transform 1 0 3910 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8050_
timestamp 0
transform 1 0 4530 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8051_
timestamp 0
transform 1 0 3590 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8052_
timestamp 0
transform 1 0 3030 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8053_
timestamp 0
transform 1 0 2870 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8054_
timestamp 0
transform 1 0 4590 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8055_
timestamp 0
transform -1 0 5370 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8056_
timestamp 0
transform -1 0 1270 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8057_
timestamp 0
transform 1 0 1530 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8058_
timestamp 0
transform 1 0 2350 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8059_
timestamp 0
transform 1 0 2610 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8060_
timestamp 0
transform 1 0 2450 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8061_
timestamp 0
transform 1 0 3470 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8062_
timestamp 0
transform -1 0 3910 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8063_
timestamp 0
transform 1 0 3750 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8064_
timestamp 0
transform 1 0 3570 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8065_
timestamp 0
transform 1 0 4130 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8066_
timestamp 0
transform 1 0 3770 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8067_
timestamp 0
transform -1 0 3990 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8068_
timestamp 0
transform -1 0 2810 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8069_
timestamp 0
transform -1 0 2910 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8070_
timestamp 0
transform -1 0 3050 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8071_
timestamp 0
transform 1 0 3810 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8072_
timestamp 0
transform 1 0 3770 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8073_
timestamp 0
transform -1 0 5110 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8074_
timestamp 0
transform 1 0 5210 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8075_
timestamp 0
transform -1 0 5110 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8076_
timestamp 0
transform 1 0 5530 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8077_
timestamp 0
transform -1 0 4470 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8078_
timestamp 0
transform -1 0 4370 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8079_
timestamp 0
transform -1 0 4950 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8080_
timestamp 0
transform 1 0 4690 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8081_
timestamp 0
transform 1 0 6810 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8082_
timestamp 0
transform 1 0 4850 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8083_
timestamp 0
transform 1 0 5210 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8084_
timestamp 0
transform -1 0 2850 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8085_
timestamp 0
transform -1 0 3030 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8086_
timestamp 0
transform -1 0 2590 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8087_
timestamp 0
transform -1 0 3690 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8088_
timestamp 0
transform 1 0 3630 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8089_
timestamp 0
transform -1 0 3510 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8090_
timestamp 0
transform 1 0 3230 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8091_
timestamp 0
transform 1 0 3110 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8092_
timestamp 0
transform 1 0 3270 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8093_
timestamp 0
transform -1 0 3330 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8094_
timestamp 0
transform -1 0 5730 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8095_
timestamp 0
transform -1 0 30 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8096_
timestamp 0
transform -1 0 2730 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8097_
timestamp 0
transform -1 0 2470 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8098_
timestamp 0
transform -1 0 2690 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8099_
timestamp 0
transform 1 0 3090 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8100_
timestamp 0
transform 1 0 3330 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8101_
timestamp 0
transform 1 0 3190 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8102_
timestamp 0
transform 1 0 2990 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8103_
timestamp 0
transform -1 0 3190 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8104_
timestamp 0
transform 1 0 3310 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8105_
timestamp 0
transform 1 0 3150 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8106_
timestamp 0
transform -1 0 2630 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8107_
timestamp 0
transform -1 0 2210 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8108_
timestamp 0
transform -1 0 2350 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8109_
timestamp 0
transform 1 0 3430 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8110_
timestamp 0
transform -1 0 3610 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8111_
timestamp 0
transform 1 0 4750 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8112_
timestamp 0
transform -1 0 2110 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8113_
timestamp 0
transform -1 0 2310 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8114_
timestamp 0
transform 1 0 2110 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8115_
timestamp 0
transform -1 0 3490 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8116_
timestamp 0
transform 1 0 3150 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8117_
timestamp 0
transform -1 0 3310 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8118_
timestamp 0
transform 1 0 3750 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8119_
timestamp 0
transform 1 0 4790 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8120_
timestamp 0
transform 1 0 5050 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8121_
timestamp 0
transform 1 0 5330 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8122_
timestamp 0
transform -1 0 4910 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8123_
timestamp 0
transform -1 0 4970 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8124_
timestamp 0
transform -1 0 4790 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8125_
timestamp 0
transform -1 0 4650 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8126_
timestamp 0
transform -1 0 4490 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8127_
timestamp 0
transform 1 0 4710 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8128_
timestamp 0
transform 1 0 7010 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__8129_
timestamp 0
transform 1 0 7170 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__8130_
timestamp 0
transform 1 0 7030 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__8131_
timestamp 0
transform 1 0 4470 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8132_
timestamp 0
transform 1 0 5190 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8133_
timestamp 0
transform -1 0 1890 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8134_
timestamp 0
transform -1 0 1950 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8135_
timestamp 0
transform 1 0 4050 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8136_
timestamp 0
transform -1 0 4050 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8137_
timestamp 0
transform 1 0 4170 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8138_
timestamp 0
transform 1 0 4330 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8139_
timestamp 0
transform -1 0 4670 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8140_
timestamp 0
transform 1 0 4630 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8141_
timestamp 0
transform -1 0 4250 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8142_
timestamp 0
transform 1 0 4490 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8143_
timestamp 0
transform 1 0 4350 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8144_
timestamp 0
transform 1 0 4930 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8145_
timestamp 0
transform -1 0 4790 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8146_
timestamp 0
transform -1 0 4770 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8147_
timestamp 0
transform 1 0 5010 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8148_
timestamp 0
transform 1 0 5250 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8149_
timestamp 0
transform -1 0 5170 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8150_
timestamp 0
transform 1 0 4850 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8151_
timestamp 0
transform -1 0 5090 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8152_
timestamp 0
transform -1 0 1070 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8153_
timestamp 0
transform 1 0 3890 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8154_
timestamp 0
transform 1 0 4330 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8155_
timestamp 0
transform 1 0 3530 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8156_
timestamp 0
transform -1 0 4250 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8157_
timestamp 0
transform -1 0 4610 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8158_
timestamp 0
transform 1 0 2930 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8159_
timestamp 0
transform -1 0 2550 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8160_
timestamp 0
transform -1 0 4510 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8161_
timestamp 0
transform -1 0 1870 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8162_
timestamp 0
transform -1 0 1530 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8163_
timestamp 0
transform -1 0 1570 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8164_
timestamp 0
transform 1 0 1830 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8165_
timestamp 0
transform 1 0 1530 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8166_
timestamp 0
transform -1 0 1350 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8167_
timestamp 0
transform 1 0 5930 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8168_
timestamp 0
transform -1 0 2850 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8169_
timestamp 0
transform 1 0 1550 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8170_
timestamp 0
transform 1 0 1390 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8171_
timestamp 0
transform 1 0 730 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8172_
timestamp 0
transform 1 0 970 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8173_
timestamp 0
transform 1 0 830 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8174_
timestamp 0
transform 1 0 1950 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8175_
timestamp 0
transform 1 0 2110 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8176_
timestamp 0
transform 1 0 2330 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__8177_
timestamp 0
transform -1 0 2430 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8178_
timestamp 0
transform 1 0 2630 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8179_
timestamp 0
transform -1 0 2790 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8180_
timestamp 0
transform -1 0 3390 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8181_
timestamp 0
transform -1 0 2270 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8182_
timestamp 0
transform 1 0 1710 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__8183_
timestamp 0
transform -1 0 690 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8184_
timestamp 0
transform -1 0 410 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8185_
timestamp 0
transform -1 0 550 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8186_
timestamp 0
transform -1 0 1710 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8187_
timestamp 0
transform 1 0 670 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8188_
timestamp 0
transform 1 0 1630 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8189_
timestamp 0
transform -1 0 690 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8190_
timestamp 0
transform 1 0 710 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8191_
timestamp 0
transform 1 0 770 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8192_
timestamp 0
transform -1 0 270 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__8193_
timestamp 0
transform -1 0 830 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8194_
timestamp 0
transform -1 0 610 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8195_
timestamp 0
transform 1 0 690 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__8196_
timestamp 0
transform 1 0 530 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__8197_
timestamp 0
transform 1 0 390 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__8198_
timestamp 0
transform 1 0 670 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__8199_
timestamp 0
transform 1 0 970 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__8200_
timestamp 0
transform 1 0 1090 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8201_
timestamp 0
transform 1 0 1250 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8202_
timestamp 0
transform -1 0 2790 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8203_
timestamp 0
transform -1 0 950 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8204_
timestamp 0
transform -1 0 1390 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__8205_
timestamp 0
transform -1 0 450 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8206_
timestamp 0
transform -1 0 770 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8207_
timestamp 0
transform 1 0 990 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8208_
timestamp 0
transform -1 0 750 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8209_
timestamp 0
transform 1 0 1030 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8210_
timestamp 0
transform 1 0 510 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8211_
timestamp 0
transform -1 0 30 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8212_
timestamp 0
transform -1 0 650 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8213_
timestamp 0
transform -1 0 490 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8214_
timestamp 0
transform -1 0 350 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8215_
timestamp 0
transform 1 0 10 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8216_
timestamp 0
transform 1 0 10 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__8217_
timestamp 0
transform 1 0 150 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__8218_
timestamp 0
transform 1 0 150 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8219_
timestamp 0
transform 1 0 1090 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8220_
timestamp 0
transform -1 0 970 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8221_
timestamp 0
transform 1 0 1250 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8222_
timestamp 0
transform -1 0 2470 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8223_
timestamp 0
transform -1 0 2130 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8224_
timestamp 0
transform 1 0 470 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8225_
timestamp 0
transform 1 0 570 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8226_
timestamp 0
transform -1 0 590 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8227_
timestamp 0
transform 1 0 390 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8228_
timestamp 0
transform -1 0 270 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8229_
timestamp 0
transform -1 0 30 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8230_
timestamp 0
transform 1 0 130 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8231_
timestamp 0
transform -1 0 290 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8232_
timestamp 0
transform 1 0 230 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8233_
timestamp 0
transform 1 0 330 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8234_
timestamp 0
transform -1 0 30 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8235_
timestamp 0
transform 1 0 350 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8236_
timestamp 0
transform 1 0 470 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8237_
timestamp 0
transform 1 0 690 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8238_
timestamp 0
transform -1 0 550 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__8239_
timestamp 0
transform -1 0 430 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__8240_
timestamp 0
transform -1 0 650 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8241_
timestamp 0
transform 1 0 490 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8242_
timestamp 0
transform 1 0 1110 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8243_
timestamp 0
transform 1 0 1170 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8244_
timestamp 0
transform -1 0 1970 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8245_
timestamp 0
transform -1 0 2790 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8246_
timestamp 0
transform -1 0 190 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8247_
timestamp 0
transform -1 0 850 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__8248_
timestamp 0
transform 1 0 170 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8249_
timestamp 0
transform -1 0 290 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__8250_
timestamp 0
transform -1 0 350 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8251_
timestamp 0
transform 1 0 410 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8252_
timestamp 0
transform -1 0 170 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8253_
timestamp 0
transform -1 0 190 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8254_
timestamp 0
transform 1 0 650 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8255_
timestamp 0
transform -1 0 770 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8256_
timestamp 0
transform 1 0 870 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8257_
timestamp 0
transform -1 0 830 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8258_
timestamp 0
transform 1 0 350 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8259_
timestamp 0
transform -1 0 30 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8260_
timestamp 0
transform 1 0 130 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8261_
timestamp 0
transform 1 0 110 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8262_
timestamp 0
transform 1 0 490 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8263_
timestamp 0
transform 1 0 10 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8264_
timestamp 0
transform -1 0 250 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8265_
timestamp 0
transform 1 0 150 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8266_
timestamp 0
transform 1 0 770 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8267_
timestamp 0
transform -1 0 790 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8268_
timestamp 0
transform -1 0 670 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8269_
timestamp 0
transform -1 0 830 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8270_
timestamp 0
transform 1 0 890 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8271_
timestamp 0
transform -1 0 2490 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8272_
timestamp 0
transform -1 0 2150 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8273_
timestamp 0
transform 1 0 970 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8274_
timestamp 0
transform -1 0 2630 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8275_
timestamp 0
transform -1 0 2270 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8276_
timestamp 0
transform 1 0 890 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8277_
timestamp 0
transform -1 0 990 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8278_
timestamp 0
transform 1 0 1030 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8279_
timestamp 0
transform -1 0 370 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8280_
timestamp 0
transform -1 0 30 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8281_
timestamp 0
transform -1 0 530 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8282_
timestamp 0
transform 1 0 150 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8283_
timestamp 0
transform -1 0 30 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8284_
timestamp 0
transform -1 0 30 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8285_
timestamp 0
transform -1 0 30 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8286_
timestamp 0
transform -1 0 210 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8287_
timestamp 0
transform 1 0 130 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8288_
timestamp 0
transform 1 0 290 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8289_
timestamp 0
transform 1 0 450 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8290_
timestamp 0
transform 1 0 470 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8291_
timestamp 0
transform 1 0 1010 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8292_
timestamp 0
transform 1 0 1370 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8293_
timestamp 0
transform 1 0 1510 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8294_
timestamp 0
transform -1 0 1990 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8295_
timestamp 0
transform 1 0 290 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8296_
timestamp 0
transform 1 0 310 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8297_
timestamp 0
transform 1 0 550 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8298_
timestamp 0
transform -1 0 630 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8299_
timestamp 0
transform -1 0 490 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8300_
timestamp 0
transform 1 0 590 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8301_
timestamp 0
transform 1 0 610 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8302_
timestamp 0
transform -1 0 990 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8303_
timestamp 0
transform 1 0 130 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8304_
timestamp 0
transform -1 0 170 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8305_
timestamp 0
transform 1 0 710 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8306_
timestamp 0
transform 1 0 10 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8307_
timestamp 0
transform -1 0 30 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8308_
timestamp 0
transform -1 0 270 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8309_
timestamp 0
transform -1 0 430 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8310_
timestamp 0
transform 1 0 110 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8311_
timestamp 0
transform 1 0 270 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8312_
timestamp 0
transform 1 0 410 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8313_
timestamp 0
transform 1 0 570 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8314_
timestamp 0
transform 1 0 1110 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8315_
timestamp 0
transform 1 0 1250 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8316_
timestamp 0
transform 1 0 1410 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8317_
timestamp 0
transform -1 0 3190 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8318_
timestamp 0
transform 1 0 430 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8319_
timestamp 0
transform 1 0 410 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8320_
timestamp 0
transform 1 0 450 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8321_
timestamp 0
transform -1 0 170 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8322_
timestamp 0
transform 1 0 290 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8323_
timestamp 0
transform -1 0 150 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8324_
timestamp 0
transform -1 0 570 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8325_
timestamp 0
transform 1 0 250 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8326_
timestamp 0
transform -1 0 410 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8327_
timestamp 0
transform -1 0 30 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8328_
timestamp 0
transform -1 0 170 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8329_
timestamp 0
transform -1 0 30 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8330_
timestamp 0
transform -1 0 310 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8331_
timestamp 0
transform -1 0 530 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8332_
timestamp 0
transform 1 0 550 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8333_
timestamp 0
transform 1 0 690 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8334_
timestamp 0
transform 1 0 690 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8335_
timestamp 0
transform 1 0 850 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8336_
timestamp 0
transform 1 0 650 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8337_
timestamp 0
transform 1 0 710 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8338_
timestamp 0
transform 1 0 850 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8339_
timestamp 0
transform 1 0 950 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8340_
timestamp 0
transform 1 0 1090 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8341_
timestamp 0
transform -1 0 2870 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8342_
timestamp 0
transform 1 0 3490 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8343_
timestamp 0
transform -1 0 550 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8344_
timestamp 0
transform -1 0 670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8345_
timestamp 0
transform 1 0 770 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8346_
timestamp 0
transform 1 0 510 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8347_
timestamp 0
transform -1 0 410 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8348_
timestamp 0
transform -1 0 150 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8349_
timestamp 0
transform -1 0 170 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8350_
timestamp 0
transform -1 0 30 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8351_
timestamp 0
transform 1 0 270 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8352_
timestamp 0
transform -1 0 670 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8353_
timestamp 0
transform 1 0 750 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8354_
timestamp 0
transform -1 0 830 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8355_
timestamp 0
transform 1 0 1230 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8356_
timestamp 0
transform 1 0 1390 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8357_
timestamp 0
transform -1 0 3150 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8358_
timestamp 0
transform 1 0 3350 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8359_
timestamp 0
transform 1 0 4550 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8360_
timestamp 0
transform -1 0 4290 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8361_
timestamp 0
transform -1 0 4430 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8362_
timestamp 0
transform 1 0 4090 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8363_
timestamp 0
transform 1 0 5810 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8364_
timestamp 0
transform -1 0 5210 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8365_
timestamp 0
transform 1 0 5670 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8366_
timestamp 0
transform -1 0 3970 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8367_
timestamp 0
transform 1 0 730 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8368_
timestamp 0
transform 1 0 590 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8369_
timestamp 0
transform 1 0 1230 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__8370_
timestamp 0
transform -1 0 1110 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__8371_
timestamp 0
transform 1 0 1250 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8372_
timestamp 0
transform -1 0 1710 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8373_
timestamp 0
transform -1 0 2710 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8374_
timestamp 0
transform -1 0 2670 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8375_
timestamp 0
transform 1 0 1130 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8376_
timestamp 0
transform -1 0 890 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8377_
timestamp 0
transform -1 0 1010 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8378_
timestamp 0
transform 1 0 1990 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8379_
timestamp 0
transform 1 0 2830 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8380_
timestamp 0
transform 1 0 2930 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8381_
timestamp 0
transform -1 0 2750 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8382_
timestamp 0
transform -1 0 2730 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8383_
timestamp 0
transform 1 0 1810 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__8384_
timestamp 0
transform -1 0 1810 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8385_
timestamp 0
transform -1 0 5350 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8386_
timestamp 0
transform -1 0 5470 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8387_
timestamp 0
transform 1 0 2930 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8388_
timestamp 0
transform 1 0 1870 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8389_
timestamp 0
transform -1 0 290 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8390_
timestamp 0
transform -1 0 390 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8391_
timestamp 0
transform 1 0 810 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8392_
timestamp 0
transform -1 0 890 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8393_
timestamp 0
transform -1 0 1010 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8394_
timestamp 0
transform -1 0 1090 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8395_
timestamp 0
transform -1 0 950 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8396_
timestamp 0
transform 1 0 1710 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8397_
timestamp 0
transform 1 0 2470 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8398_
timestamp 0
transform 1 0 1190 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8399_
timestamp 0
transform -1 0 1790 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8400_
timestamp 0
transform -1 0 2590 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8401_
timestamp 0
transform 1 0 2510 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8402_
timestamp 0
transform 1 0 2610 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8403_
timestamp 0
transform -1 0 2370 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8404_
timestamp 0
transform -1 0 2490 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8405_
timestamp 0
transform -1 0 2370 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8406_
timestamp 0
transform 1 0 2490 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8407_
timestamp 0
transform 1 0 2630 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8408_
timestamp 0
transform -1 0 2590 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8409_
timestamp 0
transform -1 0 3550 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8410_
timestamp 0
transform -1 0 2330 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8411_
timestamp 0
transform 1 0 2290 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8412_
timestamp 0
transform -1 0 990 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8413_
timestamp 0
transform 1 0 1110 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8414_
timestamp 0
transform -1 0 1270 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8415_
timestamp 0
transform -1 0 1390 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8416_
timestamp 0
transform 1 0 4030 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8417_
timestamp 0
transform 1 0 1410 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8418_
timestamp 0
transform -1 0 1550 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8419_
timestamp 0
transform 1 0 1590 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8420_
timestamp 0
transform 1 0 2010 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8421_
timestamp 0
transform 1 0 2270 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8422_
timestamp 0
transform 1 0 2130 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8423_
timestamp 0
transform -1 0 2570 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8424_
timestamp 0
transform -1 0 2290 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8425_
timestamp 0
transform 1 0 1950 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8426_
timestamp 0
transform 1 0 2430 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8427_
timestamp 0
transform -1 0 2090 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8428_
timestamp 0
transform 1 0 2210 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8429_
timestamp 0
transform -1 0 2050 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8430_
timestamp 0
transform 1 0 2170 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8431_
timestamp 0
transform 1 0 3370 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8432_
timestamp 0
transform -1 0 2070 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8433_
timestamp 0
transform -1 0 1730 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8434_
timestamp 0
transform -1 0 850 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8435_
timestamp 0
transform -1 0 910 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8436_
timestamp 0
transform 1 0 870 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8437_
timestamp 0
transform -1 0 1390 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8438_
timestamp 0
transform -1 0 2830 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8439_
timestamp 0
transform 1 0 1650 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8440_
timestamp 0
transform -1 0 1810 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8441_
timestamp 0
transform -1 0 1930 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8442_
timestamp 0
transform -1 0 2150 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8443_
timestamp 0
transform 1 0 2210 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8444_
timestamp 0
transform 1 0 2070 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8445_
timestamp 0
transform 1 0 2510 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8446_
timestamp 0
transform -1 0 2570 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8447_
timestamp 0
transform -1 0 2390 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8448_
timestamp 0
transform -1 0 2430 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8449_
timestamp 0
transform 1 0 1810 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8450_
timestamp 0
transform 1 0 1810 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8451_
timestamp 0
transform 1 0 1950 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8452_
timestamp 0
transform -1 0 2370 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8453_
timestamp 0
transform 1 0 2650 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8454_
timestamp 0
transform -1 0 1010 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8455_
timestamp 0
transform 1 0 1110 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8456_
timestamp 0
transform -1 0 1430 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8457_
timestamp 0
transform -1 0 1550 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8458_
timestamp 0
transform 1 0 1670 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8459_
timestamp 0
transform 1 0 1550 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8460_
timestamp 0
transform 1 0 2150 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8461_
timestamp 0
transform -1 0 2430 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8462_
timestamp 0
transform -1 0 1850 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8463_
timestamp 0
transform 1 0 2570 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8464_
timestamp 0
transform 1 0 1990 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8465_
timestamp 0
transform 1 0 2410 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8466_
timestamp 0
transform -1 0 3110 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8467_
timestamp 0
transform 1 0 2110 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8468_
timestamp 0
transform -1 0 2290 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8469_
timestamp 0
transform 1 0 2950 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8470_
timestamp 0
transform 1 0 3390 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8471_
timestamp 0
transform 1 0 4210 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8472_
timestamp 0
transform -1 0 4090 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8473_
timestamp 0
transform 1 0 4150 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8474_
timestamp 0
transform -1 0 4250 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8475_
timestamp 0
transform 1 0 4510 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8476_
timestamp 0
transform -1 0 3950 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8477_
timestamp 0
transform -1 0 2290 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8478_
timestamp 0
transform -1 0 1190 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8479_
timestamp 0
transform 1 0 1250 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8480_
timestamp 0
transform -1 0 1290 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8481_
timestamp 0
transform -1 0 1410 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8482_
timestamp 0
transform 1 0 1910 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8483_
timestamp 0
transform 1 0 2410 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8484_
timestamp 0
transform 1 0 1870 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8485_
timestamp 0
transform -1 0 1750 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8486_
timestamp 0
transform -1 0 1550 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8487_
timestamp 0
transform -1 0 1430 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8488_
timestamp 0
transform 1 0 2690 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8489_
timestamp 0
transform 1 0 3410 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8490_
timestamp 0
transform -1 0 2570 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8491_
timestamp 0
transform 1 0 3530 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8492_
timestamp 0
transform -1 0 3970 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8493_
timestamp 0
transform 1 0 4070 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8494_
timestamp 0
transform 1 0 4230 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8495_
timestamp 0
transform -1 0 4390 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8496_
timestamp 0
transform -1 0 4210 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8497_
timestamp 0
transform -1 0 2030 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8498_
timestamp 0
transform 1 0 1290 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8499_
timestamp 0
transform -1 0 1430 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8500_
timestamp 0
transform -1 0 1470 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8501_
timestamp 0
transform 1 0 2190 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8502_
timestamp 0
transform -1 0 1710 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8503_
timestamp 0
transform -1 0 1550 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8504_
timestamp 0
transform 1 0 2050 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8505_
timestamp 0
transform -1 0 2370 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8506_
timestamp 0
transform -1 0 2650 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8507_
timestamp 0
transform 1 0 2490 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8508_
timestamp 0
transform -1 0 3030 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8509_
timestamp 0
transform 1 0 2810 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8510_
timestamp 0
transform -1 0 2850 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8511_
timestamp 0
transform -1 0 3830 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8512_
timestamp 0
transform 1 0 3670 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8513_
timestamp 0
transform 1 0 3410 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8514_
timestamp 0
transform 1 0 3150 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8515_
timestamp 0
transform 1 0 3230 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8516_
timestamp 0
transform -1 0 3290 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8517_
timestamp 0
transform 1 0 2970 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8518_
timestamp 0
transform -1 0 3150 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8519_
timestamp 0
transform 1 0 3290 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8520_
timestamp 0
transform 1 0 3530 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8521_
timestamp 0
transform -1 0 3930 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8522_
timestamp 0
transform -1 0 4050 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8523_
timestamp 0
transform -1 0 4370 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8524_
timestamp 0
transform -1 0 2750 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8525_
timestamp 0
transform 1 0 1790 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8526_
timestamp 0
transform -1 0 1090 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8527_
timestamp 0
transform 1 0 1190 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8528_
timestamp 0
transform 1 0 1150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8529_
timestamp 0
transform 1 0 1190 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8530_
timestamp 0
transform 1 0 1090 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8531_
timestamp 0
transform -1 0 1930 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8532_
timestamp 0
transform -1 0 1490 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8533_
timestamp 0
transform 1 0 1610 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8534_
timestamp 0
transform 1 0 1750 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8535_
timestamp 0
transform 1 0 1350 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8536_
timestamp 0
transform -1 0 1930 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8537_
timestamp 0
transform -1 0 2090 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8538_
timestamp 0
transform -1 0 2870 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8539_
timestamp 0
transform 1 0 2990 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8540_
timestamp 0
transform 1 0 3690 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8541_
timestamp 0
transform 1 0 3790 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8542_
timestamp 0
transform -1 0 3970 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8543_
timestamp 0
transform -1 0 2210 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__8544_
timestamp 0
transform -1 0 2910 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8545_
timestamp 0
transform -1 0 2770 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8546_
timestamp 0
transform -1 0 2130 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8547_
timestamp 0
transform 1 0 1650 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8548_
timestamp 0
transform -1 0 1610 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8549_
timestamp 0
transform -1 0 1470 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8550_
timestamp 0
transform -1 0 1630 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8551_
timestamp 0
transform 1 0 1670 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8552_
timestamp 0
transform 1 0 1390 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__8553_
timestamp 0
transform 1 0 1830 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8554_
timestamp 0
transform 1 0 1970 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8555_
timestamp 0
transform 1 0 1710 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8556_
timestamp 0
transform 1 0 1710 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8557_
timestamp 0
transform 1 0 1830 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8558_
timestamp 0
transform 1 0 1990 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8559_
timestamp 0
transform 1 0 2150 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8560_
timestamp 0
transform 1 0 1830 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8561_
timestamp 0
transform 1 0 2510 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8562_
timestamp 0
transform -1 0 2670 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8563_
timestamp 0
transform 1 0 2990 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8564_
timestamp 0
transform 1 0 2390 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8565_
timestamp 0
transform 1 0 2250 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8566_
timestamp 0
transform -1 0 1490 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8567_
timestamp 0
transform 1 0 1670 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8568_
timestamp 0
transform -1 0 1730 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8569_
timestamp 0
transform -1 0 1810 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8570_
timestamp 0
transform 1 0 1910 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8571_
timestamp 0
transform 1 0 2210 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8572_
timestamp 0
transform 1 0 2070 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8573_
timestamp 0
transform -1 0 1710 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8574_
timestamp 0
transform -1 0 2190 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8575_
timestamp 0
transform 1 0 2310 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8576_
timestamp 0
transform 1 0 2450 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8577_
timestamp 0
transform 1 0 2590 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8578_
timestamp 0
transform -1 0 3990 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8579_
timestamp 0
transform -1 0 2070 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8580_
timestamp 0
transform -1 0 1790 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8581_
timestamp 0
transform -1 0 1830 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8582_
timestamp 0
transform -1 0 1950 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8583_
timestamp 0
transform -1 0 1930 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8584_
timestamp 0
transform -1 0 1330 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8585_
timestamp 0
transform -1 0 1290 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8586_
timestamp 0
transform -1 0 1570 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8587_
timestamp 0
transform -1 0 1550 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8588_
timestamp 0
transform 1 0 1290 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8589_
timestamp 0
transform 1 0 1550 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8590_
timestamp 0
transform 1 0 1410 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8591_
timestamp 0
transform -1 0 1030 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8592_
timestamp 0
transform 1 0 1170 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8593_
timestamp 0
transform 1 0 1170 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8594_
timestamp 0
transform 1 0 1330 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8595_
timestamp 0
transform 1 0 1710 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8596_
timestamp 0
transform 1 0 1850 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8597_
timestamp 0
transform 1 0 1990 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8598_
timestamp 0
transform -1 0 3670 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8599_
timestamp 0
transform 1 0 2790 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8600_
timestamp 0
transform 1 0 1450 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8601_
timestamp 0
transform -1 0 1570 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8602_
timestamp 0
transform 1 0 530 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8603_
timestamp 0
transform 1 0 390 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8604_
timestamp 0
transform -1 0 270 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8605_
timestamp 0
transform 1 0 250 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8606_
timestamp 0
transform 1 0 2110 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8607_
timestamp 0
transform 1 0 2250 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8608_
timestamp 0
transform 1 0 2390 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8609_
timestamp 0
transform 1 0 5950 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8610_
timestamp 0
transform -1 0 6010 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8611_
timestamp 0
transform -1 0 5610 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8612_
timestamp 0
transform 1 0 5830 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8613_
timestamp 0
transform 1 0 5690 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8614_
timestamp 0
transform 1 0 5670 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8615_
timestamp 0
transform -1 0 4590 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8616_
timestamp 0
transform -1 0 4730 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8617_
timestamp 0
transform 1 0 6590 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8618_
timestamp 0
transform 1 0 6430 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8619_
timestamp 0
transform 1 0 6770 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8620_
timestamp 0
transform 1 0 6610 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8621_
timestamp 0
transform 1 0 6310 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8622_
timestamp 0
transform 1 0 6150 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8623_
timestamp 0
transform 1 0 6390 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8624_
timestamp 0
transform -1 0 6110 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8625_
timestamp 0
transform 1 0 6150 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8626_
timestamp 0
transform -1 0 6270 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8627_
timestamp 0
transform 1 0 6290 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8628_
timestamp 0
transform -1 0 6370 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8629_
timestamp 0
transform 1 0 6210 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8630_
timestamp 0
transform 1 0 6950 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8631_
timestamp 0
transform -1 0 6830 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8632_
timestamp 0
transform -1 0 6050 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8633_
timestamp 0
transform 1 0 6070 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8634_
timestamp 0
transform 1 0 5230 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8635_
timestamp 0
transform -1 0 5550 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8636_
timestamp 0
transform 1 0 5350 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8637_
timestamp 0
transform 1 0 5070 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8638_
timestamp 0
transform -1 0 5030 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8639_
timestamp 0
transform -1 0 5170 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8640_
timestamp 0
transform 1 0 6050 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8641_
timestamp 0
transform -1 0 6570 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8642_
timestamp 0
transform 1 0 6690 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8643_
timestamp 0
transform -1 0 6730 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8644_
timestamp 0
transform 1 0 6530 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8645_
timestamp 0
transform 1 0 6070 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8646_
timestamp 0
transform 1 0 6410 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8647_
timestamp 0
transform -1 0 6270 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8648_
timestamp 0
transform 1 0 5770 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8649_
timestamp 0
transform 1 0 5670 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8650_
timestamp 0
transform -1 0 5470 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8651_
timestamp 0
transform 1 0 6030 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8652_
timestamp 0
transform 1 0 5330 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8653_
timestamp 0
transform 1 0 6010 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8654_
timestamp 0
transform -1 0 5910 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8655_
timestamp 0
transform -1 0 6170 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8656_
timestamp 0
transform 1 0 6130 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8657_
timestamp 0
transform 1 0 5990 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8658_
timestamp 0
transform -1 0 5850 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8659_
timestamp 0
transform -1 0 5970 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8660_
timestamp 0
transform -1 0 7230 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8661_
timestamp 0
transform 1 0 7110 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8662_
timestamp 0
transform 1 0 6430 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8663_
timestamp 0
transform 1 0 6570 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8664_
timestamp 0
transform 1 0 6730 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8665_
timestamp 0
transform 1 0 6930 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8666_
timestamp 0
transform 1 0 6810 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8667_
timestamp 0
transform -1 0 6770 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8668_
timestamp 0
transform 1 0 6270 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8669_
timestamp 0
transform 1 0 7310 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8670_
timestamp 0
transform 1 0 7150 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8671_
timestamp 0
transform 1 0 7350 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8672_
timestamp 0
transform 1 0 7330 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8673_
timestamp 0
transform 1 0 7390 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8674_
timestamp 0
transform 1 0 5850 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8675_
timestamp 0
transform -1 0 6230 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8676_
timestamp 0
transform -1 0 6090 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8677_
timestamp 0
transform 1 0 6090 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8678_
timestamp 0
transform 1 0 7430 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8679_
timestamp 0
transform -1 0 7310 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8680_
timestamp 0
transform -1 0 7230 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8681_
timestamp 0
transform 1 0 7250 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8682_
timestamp 0
transform 1 0 6730 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8683_
timestamp 0
transform 1 0 7450 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8684_
timestamp 0
transform -1 0 7550 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8685_
timestamp 0
transform 1 0 6570 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8686_
timestamp 0
transform -1 0 6890 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8687_
timestamp 0
transform -1 0 6650 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8688_
timestamp 0
transform -1 0 6750 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8689_
timestamp 0
transform 1 0 7090 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8690_
timestamp 0
transform 1 0 6790 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8691_
timestamp 0
transform 1 0 6830 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8692_
timestamp 0
transform -1 0 5210 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8693_
timestamp 0
transform 1 0 5590 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8694_
timestamp 0
transform -1 0 5870 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8695_
timestamp 0
transform 1 0 5710 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8696_
timestamp 0
transform 1 0 5990 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8697_
timestamp 0
transform 1 0 6150 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8698_
timestamp 0
transform 1 0 6130 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8699_
timestamp 0
transform -1 0 6310 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8700_
timestamp 0
transform -1 0 6290 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8701_
timestamp 0
transform 1 0 6370 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8702_
timestamp 0
transform 1 0 6510 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8703_
timestamp 0
transform 1 0 7070 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8704_
timestamp 0
transform -1 0 7030 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8705_
timestamp 0
transform 1 0 6170 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8706_
timestamp 0
transform 1 0 7210 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8707_
timestamp 0
transform -1 0 6530 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8708_
timestamp 0
transform 1 0 6610 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8709_
timestamp 0
transform 1 0 6750 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8710_
timestamp 0
transform 1 0 6890 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8711_
timestamp 0
transform 1 0 7030 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8712_
timestamp 0
transform -1 0 6670 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8713_
timestamp 0
transform 1 0 7150 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8714_
timestamp 0
transform -1 0 6550 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8715_
timestamp 0
transform 1 0 7370 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8716_
timestamp 0
transform -1 0 7250 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8717_
timestamp 0
transform 1 0 6390 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8718_
timestamp 0
transform 1 0 6010 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8719_
timestamp 0
transform -1 0 6450 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8720_
timestamp 0
transform 1 0 6550 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8721_
timestamp 0
transform 1 0 5490 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8722_
timestamp 0
transform 1 0 5670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8723_
timestamp 0
transform -1 0 5370 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8724_
timestamp 0
transform 1 0 5390 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8725_
timestamp 0
transform 1 0 6470 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8726_
timestamp 0
transform -1 0 6430 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8727_
timestamp 0
transform -1 0 6650 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8728_
timestamp 0
transform -1 0 6710 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8729_
timestamp 0
transform -1 0 6550 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8730_
timestamp 0
transform 1 0 5930 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8731_
timestamp 0
transform -1 0 6070 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8732_
timestamp 0
transform -1 0 6150 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8733_
timestamp 0
transform -1 0 5890 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8734_
timestamp 0
transform -1 0 5530 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8735_
timestamp 0
transform 1 0 5790 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8736_
timestamp 0
transform 1 0 5990 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8737_
timestamp 0
transform 1 0 5870 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8738_
timestamp 0
transform 1 0 5550 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8739_
timestamp 0
transform -1 0 5410 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8740_
timestamp 0
transform 1 0 5370 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__8741_
timestamp 0
transform -1 0 4810 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__8742_
timestamp 0
transform 1 0 5730 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8743_
timestamp 0
transform 1 0 6130 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8744_
timestamp 0
transform -1 0 6290 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8745_
timestamp 0
transform -1 0 5270 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8746_
timestamp 0
transform 1 0 5230 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8747_
timestamp 0
transform -1 0 4890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8748_
timestamp 0
transform 1 0 5350 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8749_
timestamp 0
transform 1 0 4990 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8750_
timestamp 0
transform -1 0 5090 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__8751_
timestamp 0
transform 1 0 5210 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__8752_
timestamp 0
transform -1 0 4950 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__8753_
timestamp 0
transform 1 0 4270 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__8754_
timestamp 0
transform -1 0 5130 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8755_
timestamp 0
transform -1 0 4670 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__8756_
timestamp 0
transform 1 0 4050 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8757_
timestamp 0
transform 1 0 3890 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8758_
timestamp 0
transform -1 0 4030 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8759_
timestamp 0
transform -1 0 2930 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8760_
timestamp 0
transform 1 0 1010 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8761_
timestamp 0
transform -1 0 1730 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8762_
timestamp 0
transform 1 0 870 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__8763_
timestamp 0
transform 1 0 4250 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8764_
timestamp 0
transform -1 0 5210 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8765_
timestamp 0
transform -1 0 3970 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8766_
timestamp 0
transform -1 0 4130 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8767_
timestamp 0
transform -1 0 4950 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8768_
timestamp 0
transform -1 0 5070 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8769_
timestamp 0
transform 1 0 4910 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8770_
timestamp 0
transform 1 0 5190 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8771_
timestamp 0
transform -1 0 3410 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8772_
timestamp 0
transform -1 0 3530 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8773_
timestamp 0
transform -1 0 4750 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8774_
timestamp 0
transform -1 0 4870 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8775_
timestamp 0
transform 1 0 5330 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8776_
timestamp 0
transform -1 0 3770 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8777_
timestamp 0
transform 1 0 3770 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8778_
timestamp 0
transform -1 0 2750 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8779_
timestamp 0
transform -1 0 2770 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8780_
timestamp 0
transform -1 0 3930 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8781_
timestamp 0
transform 1 0 3770 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8782_
timestamp 0
transform -1 0 5210 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8783_
timestamp 0
transform 1 0 5050 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8784_
timestamp 0
transform 1 0 3250 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8785_
timestamp 0
transform 1 0 3110 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8786_
timestamp 0
transform 1 0 3110 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8787_
timestamp 0
transform 1 0 2950 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8788_
timestamp 0
transform -1 0 1670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8789_
timestamp 0
transform 1 0 1110 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8790_
timestamp 0
transform -1 0 1450 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8791_
timestamp 0
transform 1 0 1270 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__8792_
timestamp 0
transform 1 0 5610 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8793_
timestamp 0
transform -1 0 4390 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8794_
timestamp 0
transform -1 0 4770 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8795_
timestamp 0
transform 1 0 3650 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__8796_
timestamp 0
transform -1 0 3810 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8797_
timestamp 0
transform 1 0 3650 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8798_
timestamp 0
transform 1 0 5230 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8799_
timestamp 0
transform 1 0 5090 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__8800_
timestamp 0
transform 1 0 3410 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8801_
timestamp 0
transform -1 0 3550 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__8802_
timestamp 0
transform -1 0 2470 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__8803_
timestamp 0
transform 1 0 2170 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__8804_
timestamp 0
transform -1 0 1690 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8805_
timestamp 0
transform 1 0 1530 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__8806_
timestamp 0
transform 1 0 4150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8807_
timestamp 0
transform -1 0 4570 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8808_
timestamp 0
transform -1 0 4010 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8809_
timestamp 0
transform 1 0 3850 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8810_
timestamp 0
transform 1 0 5610 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8811_
timestamp 0
transform 1 0 5470 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__8812_
timestamp 0
transform 1 0 5550 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8813_
timestamp 0
transform 1 0 5390 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__8814_
timestamp 0
transform -1 0 4610 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8815_
timestamp 0
transform -1 0 4730 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__8816_
timestamp 0
transform -1 0 5290 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8817_
timestamp 0
transform 1 0 5110 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__8818_
timestamp 0
transform -1 0 5510 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__8819_
timestamp 0
transform 1 0 5490 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8820_
timestamp 0
transform 1 0 5410 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8821_
timestamp 0
transform -1 0 6010 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8822_
timestamp 0
transform 1 0 5630 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__8823_
timestamp 0
transform 1 0 5570 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__8824_
timestamp 0
transform -1 0 5710 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8825_
timestamp 0
transform 1 0 5290 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8826_
timestamp 0
transform -1 0 6410 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8827_
timestamp 0
transform 1 0 6230 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__8828_
timestamp 0
transform 1 0 6530 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8829_
timestamp 0
transform -1 0 6670 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8830_
timestamp 0
transform 1 0 6890 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8831_
timestamp 0
transform -1 0 7030 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__8832_
timestamp 0
transform 1 0 4710 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8833_
timestamp 0
transform -1 0 4890 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__8834_
timestamp 0
transform 1 0 5470 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8835_
timestamp 0
transform 1 0 5630 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__8836_
timestamp 0
transform -1 0 5330 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8837_
timestamp 0
transform -1 0 5450 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__8838_
timestamp 0
transform 1 0 5950 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8839_
timestamp 0
transform -1 0 5810 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__8920_
timestamp 0
transform 1 0 250 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__8921_
timestamp 0
transform -1 0 2790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__8922_
timestamp 0
transform -1 0 2910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__8923_
timestamp 0
transform -1 0 4170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__8924_
timestamp 0
transform -1 0 4030 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__8925_
timestamp 0
transform 1 0 4950 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__8926_
timestamp 0
transform -1 0 4270 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__8927_
timestamp 0
transform 1 0 4150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__8928_
timestamp 0
transform 1 0 4510 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__8929_
timestamp 0
transform -1 0 4590 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__8930_
timestamp 0
transform 1 0 4450 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__8931_
timestamp 0
transform 1 0 4150 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__8932_
timestamp 0
transform 1 0 3970 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__8933_
timestamp 0
transform 1 0 3970 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__8934_
timestamp 0
transform 1 0 3710 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__8935_
timestamp 0
transform 1 0 3610 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__8936_
timestamp 0
transform 1 0 4290 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__8937_
timestamp 0
transform 1 0 4450 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__8938_
timestamp 0
transform 1 0 4870 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__8939_
timestamp 0
transform -1 0 4610 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__8940_
timestamp 0
transform -1 0 4910 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__8941_
timestamp 0
transform -1 0 4770 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__8942_
timestamp 0
transform 1 0 3070 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__8943_
timestamp 0
transform 1 0 4610 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__8944_
timestamp 0
transform 1 0 5150 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__8945_
timestamp 0
transform 1 0 5570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__8946_
timestamp 0
transform 1 0 5430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__8947_
timestamp 0
transform 1 0 6210 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__8948_
timestamp 0
transform -1 0 6010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__8949_
timestamp 0
transform 1 0 5650 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__8950_
timestamp 0
transform -1 0 5350 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__8951_
timestamp 0
transform -1 0 4010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__8952_
timestamp 0
transform 1 0 4730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__8953_
timestamp 0
transform -1 0 5050 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__8954_
timestamp 0
transform -1 0 5870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__8955_
timestamp 0
transform 1 0 5550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__8956_
timestamp 0
transform 1 0 4950 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__8957_
timestamp 0
transform -1 0 4910 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__8958_
timestamp 0
transform -1 0 4950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__8959_
timestamp 0
transform -1 0 5090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__8960_
timestamp 0
transform 1 0 4670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__8961_
timestamp 0
transform 1 0 5050 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__8962_
timestamp 0
transform 1 0 3550 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__8963_
timestamp 0
transform -1 0 4790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__8964_
timestamp 0
transform 1 0 4490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__8965_
timestamp 0
transform -1 0 5810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__8966_
timestamp 0
transform 1 0 5730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__8967_
timestamp 0
transform -1 0 5510 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__8968_
timestamp 0
transform 1 0 5190 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__8969_
timestamp 0
transform -1 0 3970 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__8970_
timestamp 0
transform -1 0 4830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__8971_
timestamp 0
transform 1 0 5930 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__8972_
timestamp 0
transform -1 0 4390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__8973_
timestamp 0
transform 1 0 4590 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__8974_
timestamp 0
transform 1 0 4190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__8975_
timestamp 0
transform -1 0 4470 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__8976_
timestamp 0
transform 1 0 4130 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__8977_
timestamp 0
transform -1 0 4330 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__8978_
timestamp 0
transform -1 0 3910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__8979_
timestamp 0
transform -1 0 2370 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__8980_
timestamp 0
transform -1 0 30 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__8981_
timestamp 0
transform -1 0 270 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__8982_
timestamp 0
transform 1 0 1430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__8983_
timestamp 0
transform -1 0 1210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__8984_
timestamp 0
transform -1 0 1350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__8985_
timestamp 0
transform -1 0 1050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__8986_
timestamp 0
transform -1 0 890 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__8987_
timestamp 0
transform -1 0 1030 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__8988_
timestamp 0
transform -1 0 1170 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__8989_
timestamp 0
transform 1 0 890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__8990_
timestamp 0
transform -1 0 630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__8991_
timestamp 0
transform -1 0 770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__8992_
timestamp 0
transform -1 0 1570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__8993_
timestamp 0
transform 1 0 1410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__8994_
timestamp 0
transform -1 0 1390 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__8995_
timestamp 0
transform 1 0 1030 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__8996_
timestamp 0
transform 1 0 1210 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__8997_
timestamp 0
transform -1 0 2490 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__8998_
timestamp 0
transform -1 0 2230 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__8999_
timestamp 0
transform -1 0 2610 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9000_
timestamp 0
transform -1 0 430 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9001_
timestamp 0
transform 1 0 3530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9002_
timestamp 0
transform 1 0 3410 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9003_
timestamp 0
transform 1 0 2690 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9004_
timestamp 0
transform -1 0 3530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9005_
timestamp 0
transform 1 0 4490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9006_
timestamp 0
transform 1 0 4550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9007_
timestamp 0
transform -1 0 3570 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9008_
timestamp 0
transform -1 0 430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9009_
timestamp 0
transform -1 0 550 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9010_
timestamp 0
transform 1 0 370 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9011_
timestamp 0
transform 1 0 10 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9012_
timestamp 0
transform -1 0 170 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9013_
timestamp 0
transform 1 0 290 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9014_
timestamp 0
transform -1 0 590 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9015_
timestamp 0
transform -1 0 750 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9016_
timestamp 0
transform -1 0 450 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9017_
timestamp 0
transform 1 0 430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9018_
timestamp 0
transform -1 0 1290 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9019_
timestamp 0
transform -1 0 130 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9020_
timestamp 0
transform -1 0 1050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9021_
timestamp 0
transform -1 0 790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9022_
timestamp 0
transform -1 0 930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9023_
timestamp 0
transform -1 0 1650 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9024_
timestamp 0
transform -1 0 1230 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9025_
timestamp 0
transform -1 0 1370 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9026_
timestamp 0
transform 1 0 1030 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9027_
timestamp 0
transform 1 0 890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9028_
timestamp 0
transform 1 0 1490 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9029_
timestamp 0
transform -1 0 1490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9030_
timestamp 0
transform -1 0 1170 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9031_
timestamp 0
transform 1 0 1670 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9032_
timestamp 0
transform 1 0 1630 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9033_
timestamp 0
transform 1 0 1450 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9034_
timestamp 0
transform 1 0 1510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9035_
timestamp 0
transform 1 0 1510 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9036_
timestamp 0
transform 1 0 710 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9037_
timestamp 0
transform 1 0 710 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9038_
timestamp 0
transform -1 0 750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9039_
timestamp 0
transform -1 0 750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9040_
timestamp 0
transform -1 0 1010 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9041_
timestamp 0
transform 1 0 710 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9042_
timestamp 0
transform -1 0 890 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9043_
timestamp 0
transform -1 0 1670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9044_
timestamp 0
transform -1 0 1550 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9045_
timestamp 0
transform 1 0 1810 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9046_
timestamp 0
transform 1 0 1670 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9047_
timestamp 0
transform 1 0 1930 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9048_
timestamp 0
transform 1 0 2630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9049_
timestamp 0
transform 1 0 2790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9050_
timestamp 0
transform 1 0 2930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9051_
timestamp 0
transform 1 0 4170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9052_
timestamp 0
transform 1 0 7490 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9053_
timestamp 0
transform -1 0 6910 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9054_
timestamp 0
transform 1 0 7110 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9055_
timestamp 0
transform -1 0 3950 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9056_
timestamp 0
transform -1 0 2090 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9057_
timestamp 0
transform -1 0 430 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9058_
timestamp 0
transform 1 0 570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9059_
timestamp 0
transform -1 0 590 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9060_
timestamp 0
transform -1 0 290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9061_
timestamp 0
transform 1 0 410 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9062_
timestamp 0
transform 1 0 550 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9063_
timestamp 0
transform 1 0 1950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9064_
timestamp 0
transform 1 0 2090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9065_
timestamp 0
transform 1 0 2070 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9066_
timestamp 0
transform 1 0 1650 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9067_
timestamp 0
transform 1 0 1930 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9068_
timestamp 0
transform 1 0 2390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9069_
timestamp 0
transform 1 0 2230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9070_
timestamp 0
transform 1 0 3250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9071_
timestamp 0
transform 1 0 3510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9072_
timestamp 0
transform 1 0 3670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9073_
timestamp 0
transform 1 0 3790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9074_
timestamp 0
transform -1 0 3370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9075_
timestamp 0
transform 1 0 3890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9076_
timestamp 0
transform 1 0 3990 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9077_
timestamp 0
transform 1 0 4350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9078_
timestamp 0
transform -1 0 4050 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9079_
timestamp 0
transform 1 0 4830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9080_
timestamp 0
transform 1 0 4450 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9081_
timestamp 0
transform 1 0 3090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9082_
timestamp 0
transform 1 0 3950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9083_
timestamp 0
transform -1 0 2910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9084_
timestamp 0
transform 1 0 1810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9085_
timestamp 0
transform 1 0 530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9086_
timestamp 0
transform -1 0 310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9087_
timestamp 0
transform -1 0 650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9088_
timestamp 0
transform -1 0 910 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9089_
timestamp 0
transform 1 0 890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9090_
timestamp 0
transform -1 0 1630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9091_
timestamp 0
transform 1 0 1510 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9092_
timestamp 0
transform 1 0 1610 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9093_
timestamp 0
transform 1 0 1530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9094_
timestamp 0
transform 1 0 2610 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9095_
timestamp 0
transform -1 0 2650 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9096_
timestamp 0
transform -1 0 2770 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9097_
timestamp 0
transform -1 0 2770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9098_
timestamp 0
transform 1 0 3150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9099_
timestamp 0
transform 1 0 3010 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9100_
timestamp 0
transform 1 0 3470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9101_
timestamp 0
transform 1 0 3590 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9102_
timestamp 0
transform 1 0 4050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9103_
timestamp 0
transform 1 0 4210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9104_
timestamp 0
transform -1 0 4570 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9105_
timestamp 0
transform 1 0 3310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9106_
timestamp 0
transform 1 0 3530 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9107_
timestamp 0
transform -1 0 190 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9108_
timestamp 0
transform -1 0 370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9109_
timestamp 0
transform 1 0 470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9110_
timestamp 0
transform 1 0 610 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9111_
timestamp 0
transform -1 0 770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9112_
timestamp 0
transform -1 0 930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9113_
timestamp 0
transform -1 0 1070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9114_
timestamp 0
transform 1 0 3310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9115_
timestamp 0
transform 1 0 3190 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9116_
timestamp 0
transform 1 0 3610 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9117_
timestamp 0
transform -1 0 2930 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9118_
timestamp 0
transform 1 0 3050 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9119_
timestamp 0
transform 1 0 3910 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9120_
timestamp 0
transform -1 0 3590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9121_
timestamp 0
transform -1 0 3450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9122_
timestamp 0
transform 1 0 3690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9123_
timestamp 0
transform 1 0 4330 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9124_
timestamp 0
transform 1 0 4890 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9125_
timestamp 0
transform 1 0 5050 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9126_
timestamp 0
transform -1 0 5810 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9127_
timestamp 0
transform -1 0 4270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9128_
timestamp 0
transform 1 0 2810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9129_
timestamp 0
transform 1 0 2910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9130_
timestamp 0
transform -1 0 430 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9131_
timestamp 0
transform 1 0 530 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9132_
timestamp 0
transform 1 0 970 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9133_
timestamp 0
transform -1 0 1050 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9134_
timestamp 0
transform -1 0 1310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9135_
timestamp 0
transform 1 0 2610 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9136_
timestamp 0
transform -1 0 3090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9137_
timestamp 0
transform -1 0 2690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9138_
timestamp 0
transform -1 0 2790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9139_
timestamp 0
transform 1 0 3350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9140_
timestamp 0
transform 1 0 3210 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9141_
timestamp 0
transform -1 0 3510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9142_
timestamp 0
transform -1 0 3630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9143_
timestamp 0
transform 1 0 4390 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9144_
timestamp 0
transform 1 0 4550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9145_
timestamp 0
transform 1 0 4690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9146_
timestamp 0
transform -1 0 4690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9147_
timestamp 0
transform -1 0 6310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9148_
timestamp 0
transform 1 0 4490 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9149_
timestamp 0
transform 1 0 3070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9150_
timestamp 0
transform 1 0 650 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9151_
timestamp 0
transform -1 0 610 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9152_
timestamp 0
transform -1 0 830 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9153_
timestamp 0
transform 1 0 4070 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9154_
timestamp 0
transform -1 0 3310 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9155_
timestamp 0
transform 1 0 2750 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9156_
timestamp 0
transform -1 0 3530 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9157_
timestamp 0
transform 1 0 4890 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9158_
timestamp 0
transform 1 0 3630 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9159_
timestamp 0
transform -1 0 3410 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9160_
timestamp 0
transform 1 0 3770 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9161_
timestamp 0
transform 1 0 5010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9162_
timestamp 0
transform 1 0 3750 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9163_
timestamp 0
transform 1 0 4070 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9164_
timestamp 0
transform -1 0 4750 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9165_
timestamp 0
transform 1 0 4650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9166_
timestamp 0
transform 1 0 5130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9167_
timestamp 0
transform 1 0 5270 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9168_
timestamp 0
transform -1 0 6150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9169_
timestamp 0
transform 1 0 5010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9170_
timestamp 0
transform -1 0 4770 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9171_
timestamp 0
transform 1 0 4190 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9172_
timestamp 0
transform -1 0 4050 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9173_
timestamp 0
transform -1 0 3750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9174_
timestamp 0
transform -1 0 3890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9175_
timestamp 0
transform -1 0 4630 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9176_
timestamp 0
transform -1 0 4170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9177_
timestamp 0
transform -1 0 2950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9178_
timestamp 0
transform 1 0 250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9179_
timestamp 0
transform -1 0 390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9180_
timestamp 0
transform 1 0 650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9181_
timestamp 0
transform -1 0 1470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9182_
timestamp 0
transform -1 0 3210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9183_
timestamp 0
transform -1 0 3350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9184_
timestamp 0
transform 1 0 3930 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9185_
timestamp 0
transform 1 0 3870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9186_
timestamp 0
transform 1 0 3990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9187_
timestamp 0
transform 1 0 3450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9188_
timestamp 0
transform 1 0 3730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9189_
timestamp 0
transform -1 0 3610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9190_
timestamp 0
transform -1 0 4130 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9191_
timestamp 0
transform 1 0 4230 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9192_
timestamp 0
transform 1 0 4490 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9193_
timestamp 0
transform 1 0 4850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9194_
timestamp 0
transform 1 0 4350 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9195_
timestamp 0
transform 1 0 4290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9196_
timestamp 0
transform 1 0 4750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9197_
timestamp 0
transform 1 0 4610 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9198_
timestamp 0
transform -1 0 4870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9199_
timestamp 0
transform -1 0 5030 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9200_
timestamp 0
transform -1 0 3710 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9201_
timestamp 0
transform -1 0 4010 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9202_
timestamp 0
transform -1 0 3870 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9203_
timestamp 0
transform -1 0 2350 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9204_
timestamp 0
transform -1 0 3190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9205_
timestamp 0
transform 1 0 1130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9206_
timestamp 0
transform -1 0 2770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9207_
timestamp 0
transform 1 0 2850 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9208_
timestamp 0
transform 1 0 2610 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9209_
timestamp 0
transform -1 0 2730 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9210_
timestamp 0
transform 1 0 2450 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9211_
timestamp 0
transform 1 0 2890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9212_
timestamp 0
transform 1 0 2990 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9213_
timestamp 0
transform 1 0 3030 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9214_
timestamp 0
transform 1 0 4170 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9215_
timestamp 0
transform 1 0 4470 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9216_
timestamp 0
transform 1 0 4450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9217_
timestamp 0
transform 1 0 4590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9218_
timestamp 0
transform -1 0 4870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9219_
timestamp 0
transform -1 0 4290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9220_
timestamp 0
transform 1 0 4410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9221_
timestamp 0
transform 1 0 5050 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9222_
timestamp 0
transform 1 0 4690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9223_
timestamp 0
transform -1 0 4570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9224_
timestamp 0
transform -1 0 4070 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9225_
timestamp 0
transform 1 0 4330 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9226_
timestamp 0
transform -1 0 3630 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9227_
timestamp 0
transform 1 0 3310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9228_
timestamp 0
transform 1 0 3510 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9229_
timestamp 0
transform 1 0 1290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9230_
timestamp 0
transform 1 0 3370 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9231_
timestamp 0
transform 1 0 3110 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9232_
timestamp 0
transform 1 0 3290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9233_
timestamp 0
transform 1 0 3430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9234_
timestamp 0
transform 1 0 3730 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9235_
timestamp 0
transform -1 0 3250 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9236_
timestamp 0
transform 1 0 3890 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9237_
timestamp 0
transform 1 0 4010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9238_
timestamp 0
transform 1 0 4430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9239_
timestamp 0
transform 1 0 4570 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9240_
timestamp 0
transform 1 0 4710 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9241_
timestamp 0
transform -1 0 5150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9242_
timestamp 0
transform -1 0 2250 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9243_
timestamp 0
transform 1 0 870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9244_
timestamp 0
transform 1 0 3390 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9245_
timestamp 0
transform 1 0 3630 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9246_
timestamp 0
transform 1 0 3490 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9247_
timestamp 0
transform -1 0 3690 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9248_
timestamp 0
transform -1 0 3270 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9249_
timestamp 0
transform 1 0 3790 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9250_
timestamp 0
transform 1 0 3710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9251_
timestamp 0
transform 1 0 4070 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9252_
timestamp 0
transform 1 0 3790 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9253_
timestamp 0
transform -1 0 3950 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9254_
timestamp 0
transform 1 0 3930 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9255_
timestamp 0
transform -1 0 4090 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9256_
timestamp 0
transform 1 0 3570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9257_
timestamp 0
transform -1 0 3870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9258_
timestamp 0
transform -1 0 4310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9259_
timestamp 0
transform 1 0 4370 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9260_
timestamp 0
transform 1 0 4210 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9261_
timestamp 0
transform 1 0 4150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9262_
timestamp 0
transform 1 0 4510 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9263_
timestamp 0
transform 1 0 4670 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9264_
timestamp 0
transform 1 0 4810 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9265_
timestamp 0
transform -1 0 4770 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9266_
timestamp 0
transform 1 0 6190 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9267_
timestamp 0
transform -1 0 4190 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9268_
timestamp 0
transform 1 0 10 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9269_
timestamp 0
transform 1 0 250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9270_
timestamp 0
transform -1 0 270 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9271_
timestamp 0
transform -1 0 30 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9272_
timestamp 0
transform -1 0 3550 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9273_
timestamp 0
transform 1 0 3790 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9274_
timestamp 0
transform 1 0 3910 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9275_
timestamp 0
transform 1 0 4050 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9276_
timestamp 0
transform -1 0 4190 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9277_
timestamp 0
transform 1 0 4430 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9278_
timestamp 0
transform -1 0 4310 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9279_
timestamp 0
transform 1 0 4290 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9280_
timestamp 0
transform 1 0 4650 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9281_
timestamp 0
transform -1 0 6070 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9282_
timestamp 0
transform 1 0 3550 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9283_
timestamp 0
transform 1 0 2530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9284_
timestamp 0
transform 1 0 2870 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9285_
timestamp 0
transform 1 0 2450 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9286_
timestamp 0
transform 1 0 1950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9287_
timestamp 0
transform 1 0 1670 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9288_
timestamp 0
transform -1 0 530 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9289_
timestamp 0
transform -1 0 1530 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9290_
timestamp 0
transform 1 0 1810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9291_
timestamp 0
transform -1 0 4230 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9292_
timestamp 0
transform -1 0 4370 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9293_
timestamp 0
transform -1 0 2350 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9294_
timestamp 0
transform -1 0 2490 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9295_
timestamp 0
transform -1 0 2350 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9296_
timestamp 0
transform -1 0 1910 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9297_
timestamp 0
transform -1 0 1910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9298_
timestamp 0
transform 1 0 1790 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9299_
timestamp 0
transform 1 0 2510 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9300_
timestamp 0
transform 1 0 2750 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9301_
timestamp 0
transform 1 0 2630 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9302_
timestamp 0
transform 1 0 1970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9303_
timestamp 0
transform 1 0 2290 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9304_
timestamp 0
transform 1 0 3170 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9305_
timestamp 0
transform -1 0 3830 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9306_
timestamp 0
transform -1 0 2190 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9307_
timestamp 0
transform 1 0 3230 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9308_
timestamp 0
transform 1 0 3090 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9309_
timestamp 0
transform 1 0 1410 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9310_
timestamp 0
transform 1 0 1250 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9311_
timestamp 0
transform -1 0 1790 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9312_
timestamp 0
transform 1 0 1830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9313_
timestamp 0
transform -1 0 2950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9314_
timestamp 0
transform -1 0 3070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9315_
timestamp 0
transform 1 0 1250 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9316_
timestamp 0
transform -1 0 2290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9317_
timestamp 0
transform -1 0 2410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9318_
timestamp 0
transform -1 0 1550 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9319_
timestamp 0
transform 1 0 1370 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9320_
timestamp 0
transform 1 0 1690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9321_
timestamp 0
transform 1 0 1930 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9322_
timestamp 0
transform -1 0 2170 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9323_
timestamp 0
transform 1 0 2110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9324_
timestamp 0
transform -1 0 2190 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9325_
timestamp 0
transform 1 0 2190 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9326_
timestamp 0
transform 1 0 2350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9327_
timestamp 0
transform 1 0 2330 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9328_
timestamp 0
transform 1 0 2470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9329_
timestamp 0
transform -1 0 2610 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9330_
timestamp 0
transform 1 0 2730 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9331_
timestamp 0
transform 1 0 3010 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9332_
timestamp 0
transform 1 0 3670 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9333_
timestamp 0
transform 1 0 4030 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9334_
timestamp 0
transform 1 0 2470 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9335_
timestamp 0
transform -1 0 2150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9336_
timestamp 0
transform 1 0 2090 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9337_
timestamp 0
transform -1 0 1970 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9338_
timestamp 0
transform 1 0 2350 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9339_
timestamp 0
transform 1 0 1830 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9340_
timestamp 0
transform 1 0 1770 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9341_
timestamp 0
transform -1 0 1790 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9342_
timestamp 0
transform -1 0 1670 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9343_
timestamp 0
transform 1 0 1670 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9344_
timestamp 0
transform 1 0 1970 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9345_
timestamp 0
transform 1 0 2210 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9346_
timestamp 0
transform 1 0 2010 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9347_
timestamp 0
transform -1 0 2010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9348_
timestamp 0
transform 1 0 2250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9349_
timestamp 0
transform 1 0 2710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9350_
timestamp 0
transform 1 0 2410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9351_
timestamp 0
transform 1 0 2810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9352_
timestamp 0
transform 1 0 3470 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9353_
timestamp 0
transform -1 0 3350 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9354_
timestamp 0
transform 1 0 3850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9355_
timestamp 0
transform 1 0 3870 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9356_
timestamp 0
transform -1 0 2590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9357_
timestamp 0
transform -1 0 2510 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9358_
timestamp 0
transform -1 0 2270 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9359_
timestamp 0
transform 1 0 2110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9360_
timestamp 0
transform -1 0 1070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9361_
timestamp 0
transform -1 0 1250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9362_
timestamp 0
transform 1 0 2030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9363_
timestamp 0
transform -1 0 1930 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9364_
timestamp 0
transform -1 0 2050 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9365_
timestamp 0
transform 1 0 1350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9366_
timestamp 0
transform -1 0 2090 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9367_
timestamp 0
transform 1 0 1910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9368_
timestamp 0
transform 1 0 1770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9369_
timestamp 0
transform 1 0 2210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9370_
timestamp 0
transform 1 0 2510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9371_
timestamp 0
transform 1 0 2070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9372_
timestamp 0
transform 1 0 2610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9373_
timestamp 0
transform 1 0 3290 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9374_
timestamp 0
transform -1 0 3170 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9375_
timestamp 0
transform 1 0 3430 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9376_
timestamp 0
transform -1 0 5450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9377_
timestamp 0
transform -1 0 2390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9378_
timestamp 0
transform -1 0 150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9379_
timestamp 0
transform -1 0 810 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9380_
timestamp 0
transform -1 0 1410 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9381_
timestamp 0
transform -1 0 1530 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9382_
timestamp 0
transform -1 0 1290 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9383_
timestamp 0
transform -1 0 1410 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9384_
timestamp 0
transform 1 0 1830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9385_
timestamp 0
transform -1 0 1750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9386_
timestamp 0
transform -1 0 1690 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9387_
timestamp 0
transform -1 0 1710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9388_
timestamp 0
transform -1 0 1550 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9389_
timestamp 0
transform -1 0 1430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9390_
timestamp 0
transform 1 0 1550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9391_
timestamp 0
transform 1 0 1950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9392_
timestamp 0
transform -1 0 1730 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9393_
timestamp 0
transform 1 0 1990 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9394_
timestamp 0
transform -1 0 2430 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9395_
timestamp 0
transform 1 0 2670 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9396_
timestamp 0
transform 1 0 2530 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9397_
timestamp 0
transform 1 0 2670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9398_
timestamp 0
transform -1 0 5630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9399_
timestamp 0
transform 1 0 4190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9400_
timestamp 0
transform 1 0 2530 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9401_
timestamp 0
transform -1 0 1790 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9402_
timestamp 0
transform -1 0 530 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9403_
timestamp 0
transform -1 0 970 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9404_
timestamp 0
transform 1 0 1270 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9405_
timestamp 0
transform 1 0 1110 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9406_
timestamp 0
transform 1 0 1550 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9407_
timestamp 0
transform 1 0 1890 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9408_
timestamp 0
transform -1 0 1530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9409_
timestamp 0
transform 1 0 1630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9410_
timestamp 0
transform 1 0 1550 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9411_
timestamp 0
transform -1 0 1670 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9412_
timestamp 0
transform -1 0 1830 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9413_
timestamp 0
transform -1 0 2150 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9414_
timestamp 0
transform 1 0 1970 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9415_
timestamp 0
transform -1 0 2250 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9416_
timestamp 0
transform -1 0 3010 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9417_
timestamp 0
transform 1 0 3110 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9418_
timestamp 0
transform 1 0 3270 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9419_
timestamp 0
transform -1 0 3810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9420_
timestamp 0
transform -1 0 5370 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9421_
timestamp 0
transform -1 0 1430 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9422_
timestamp 0
transform -1 0 650 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9423_
timestamp 0
transform -1 0 610 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9424_
timestamp 0
transform -1 0 1010 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9425_
timestamp 0
transform 1 0 990 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9426_
timestamp 0
transform -1 0 1350 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9427_
timestamp 0
transform 1 0 870 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9428_
timestamp 0
transform -1 0 1150 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9429_
timestamp 0
transform -1 0 1290 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9430_
timestamp 0
transform 1 0 1410 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9431_
timestamp 0
transform 1 0 1530 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9432_
timestamp 0
transform 1 0 1690 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9433_
timestamp 0
transform -1 0 1870 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9434_
timestamp 0
transform 1 0 2250 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9435_
timestamp 0
transform -1 0 2410 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9436_
timestamp 0
transform 1 0 2370 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9437_
timestamp 0
transform 1 0 2510 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9438_
timestamp 0
transform 1 0 2690 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9439_
timestamp 0
transform -1 0 2130 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9440_
timestamp 0
transform -1 0 2010 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9441_
timestamp 0
transform -1 0 1850 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9442_
timestamp 0
transform -1 0 1710 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9443_
timestamp 0
transform 1 0 2850 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9444_
timestamp 0
transform 1 0 3650 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9445_
timestamp 0
transform -1 0 3690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9446_
timestamp 0
transform -1 0 5210 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9447_
timestamp 0
transform -1 0 3710 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9448_
timestamp 0
transform 1 0 2630 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9449_
timestamp 0
transform 1 0 750 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9450_
timestamp 0
transform -1 0 390 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9451_
timestamp 0
transform 1 0 430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9452_
timestamp 0
transform -1 0 730 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9453_
timestamp 0
transform -1 0 130 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9454_
timestamp 0
transform -1 0 30 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9455_
timestamp 0
transform -1 0 990 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9456_
timestamp 0
transform -1 0 590 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9457_
timestamp 0
transform 1 0 430 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9458_
timestamp 0
transform 1 0 270 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9459_
timestamp 0
transform -1 0 710 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9460_
timestamp 0
transform 1 0 810 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9461_
timestamp 0
transform -1 0 1150 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9462_
timestamp 0
transform 1 0 2750 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9463_
timestamp 0
transform 1 0 3010 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9464_
timestamp 0
transform 1 0 2910 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9465_
timestamp 0
transform 1 0 3130 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9466_
timestamp 0
transform -1 0 3310 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9467_
timestamp 0
transform -1 0 1270 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9468_
timestamp 0
transform -1 0 1590 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9469_
timestamp 0
transform -1 0 1430 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__9470_
timestamp 0
transform -1 0 690 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9471_
timestamp 0
transform -1 0 630 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9472_
timestamp 0
transform -1 0 1170 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9473_
timestamp 0
transform -1 0 870 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9474_
timestamp 0
transform 1 0 870 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9475_
timestamp 0
transform 1 0 730 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9476_
timestamp 0
transform -1 0 490 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9477_
timestamp 0
transform 1 0 590 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9478_
timestamp 0
transform 1 0 770 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9479_
timestamp 0
transform 1 0 310 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9480_
timestamp 0
transform 1 0 990 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9481_
timestamp 0
transform 1 0 1110 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9482_
timestamp 0
transform 1 0 2210 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9483_
timestamp 0
transform 1 0 2490 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9484_
timestamp 0
transform 1 0 2050 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9485_
timestamp 0
transform 1 0 2350 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9486_
timestamp 0
transform -1 0 3150 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9487_
timestamp 0
transform 1 0 2990 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9488_
timestamp 0
transform -1 0 2170 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9489_
timestamp 0
transform 1 0 2270 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9490_
timestamp 0
transform -1 0 470 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9491_
timestamp 0
transform -1 0 290 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9492_
timestamp 0
transform 1 0 450 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9493_
timestamp 0
transform -1 0 410 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9494_
timestamp 0
transform 1 0 530 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9495_
timestamp 0
transform 1 0 510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9496_
timestamp 0
transform -1 0 390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9497_
timestamp 0
transform -1 0 670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9498_
timestamp 0
transform 1 0 1270 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9499_
timestamp 0
transform 1 0 2370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9500_
timestamp 0
transform 1 0 2510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9501_
timestamp 0
transform 1 0 2610 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9502_
timestamp 0
transform 1 0 5090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9503_
timestamp 0
transform 1 0 910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9504_
timestamp 0
transform 1 0 910 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9505_
timestamp 0
transform 1 0 1270 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9506_
timestamp 0
transform -1 0 1210 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9507_
timestamp 0
transform -1 0 1070 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9508_
timestamp 0
transform -1 0 310 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9509_
timestamp 0
transform 1 0 270 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9510_
timestamp 0
transform -1 0 170 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9511_
timestamp 0
transform -1 0 30 0 1 250
box -6 -8 26 248
use FILL  FILL_0__9512_
timestamp 0
transform 1 0 310 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9513_
timestamp 0
transform -1 0 30 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9514_
timestamp 0
transform -1 0 30 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9515_
timestamp 0
transform 1 0 150 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9516_
timestamp 0
transform 1 0 150 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9517_
timestamp 0
transform 1 0 130 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9518_
timestamp 0
transform -1 0 30 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__9519_
timestamp 0
transform -1 0 30 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9520_
timestamp 0
transform 1 0 170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__9521_
timestamp 0
transform 1 0 130 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__9522_
timestamp 0
transform -1 0 4930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__9523_
timestamp 0
transform -1 0 3190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9524_
timestamp 0
transform 1 0 10 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9525_
timestamp 0
transform 1 0 130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__9526_
timestamp 0
transform 1 0 2590 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9527_
timestamp 0
transform -1 0 2730 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9528_
timestamp 0
transform 1 0 2990 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9529_
timestamp 0
transform -1 0 2870 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__9530_
timestamp 0
transform 1 0 2810 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9531_
timestamp 0
transform 1 0 2950 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9532_
timestamp 0
transform 1 0 3110 0 1 730
box -6 -8 26 248
use FILL  FILL_0__9533_
timestamp 0
transform 1 0 730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9534_
timestamp 0
transform 1 0 1390 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9535_
timestamp 0
transform 1 0 1550 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9536_
timestamp 0
transform 1 0 1250 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9537_
timestamp 0
transform -1 0 1570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9538_
timestamp 0
transform 1 0 1670 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9539_
timestamp 0
transform 1 0 3590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9540_
timestamp 0
transform 1 0 3210 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9541_
timestamp 0
transform 1 0 2050 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9542_
timestamp 0
transform -1 0 1470 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9543_
timestamp 0
transform 1 0 1230 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9544_
timestamp 0
transform -1 0 1150 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9545_
timestamp 0
transform 1 0 950 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9546_
timestamp 0
transform 1 0 790 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9547_
timestamp 0
transform -1 0 830 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9548_
timestamp 0
transform 1 0 830 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9549_
timestamp 0
transform -1 0 370 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9550_
timestamp 0
transform -1 0 690 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9551_
timestamp 0
transform -1 0 510 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9552_
timestamp 0
transform -1 0 1430 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9553_
timestamp 0
transform -1 0 1290 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9554_
timestamp 0
transform -1 0 1550 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9555_
timestamp 0
transform 1 0 1650 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9556_
timestamp 0
transform 1 0 610 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9557_
timestamp 0
transform 1 0 990 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9558_
timestamp 0
transform 1 0 130 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9559_
timestamp 0
transform 1 0 10 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9560_
timestamp 0
transform -1 0 170 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9561_
timestamp 0
transform -1 0 190 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9562_
timestamp 0
transform -1 0 30 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9563_
timestamp 0
transform -1 0 30 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9564_
timestamp 0
transform -1 0 30 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9565_
timestamp 0
transform 1 0 230 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9566_
timestamp 0
transform -1 0 130 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9567_
timestamp 0
transform -1 0 550 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9568_
timestamp 0
transform -1 0 390 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9569_
timestamp 0
transform -1 0 2070 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9570_
timestamp 0
transform -1 0 150 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9571_
timestamp 0
transform 1 0 270 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9572_
timestamp 0
transform -1 0 890 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9573_
timestamp 0
transform -1 0 30 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9574_
timestamp 0
transform 1 0 430 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9575_
timestamp 0
transform -1 0 570 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9576_
timestamp 0
transform -1 0 610 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9577_
timestamp 0
transform 1 0 610 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9578_
timestamp 0
transform 1 0 750 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9579_
timestamp 0
transform -1 0 690 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9580_
timestamp 0
transform -1 0 570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9581_
timestamp 0
transform -1 0 390 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9582_
timestamp 0
transform 1 0 530 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9583_
timestamp 0
transform -1 0 1950 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9584_
timestamp 0
transform 1 0 4310 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9585_
timestamp 0
transform 1 0 3050 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9586_
timestamp 0
transform 1 0 950 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9587_
timestamp 0
transform -1 0 1130 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9588_
timestamp 0
transform 1 0 1070 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9589_
timestamp 0
transform 1 0 3150 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9590_
timestamp 0
transform 1 0 3310 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9591_
timestamp 0
transform 1 0 3430 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9592_
timestamp 0
transform 1 0 670 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9593_
timestamp 0
transform 1 0 3830 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9594_
timestamp 0
transform -1 0 3710 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9595_
timestamp 0
transform 1 0 3730 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9596_
timestamp 0
transform -1 0 3670 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9597_
timestamp 0
transform -1 0 2390 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9598_
timestamp 0
transform -1 0 1470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9599_
timestamp 0
transform -1 0 1130 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9600_
timestamp 0
transform 1 0 1350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9601_
timestamp 0
transform 1 0 1490 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9602_
timestamp 0
transform 1 0 2850 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9603_
timestamp 0
transform -1 0 2730 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9604_
timestamp 0
transform -1 0 3010 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9605_
timestamp 0
transform 1 0 3250 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9606_
timestamp 0
transform 1 0 3850 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9607_
timestamp 0
transform -1 0 3750 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9608_
timestamp 0
transform -1 0 4650 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9609_
timestamp 0
transform -1 0 4790 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9610_
timestamp 0
transform -1 0 4450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9611_
timestamp 0
transform -1 0 3570 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9612_
timestamp 0
transform -1 0 3830 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9613_
timestamp 0
transform -1 0 3130 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9614_
timestamp 0
transform 1 0 3370 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9615_
timestamp 0
transform 1 0 3950 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9616_
timestamp 0
transform 1 0 290 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9617_
timestamp 0
transform 1 0 330 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9618_
timestamp 0
transform 1 0 290 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9619_
timestamp 0
transform 1 0 470 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9620_
timestamp 0
transform -1 0 430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9621_
timestamp 0
transform -1 0 2430 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9622_
timestamp 0
transform 1 0 2430 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9623_
timestamp 0
transform -1 0 2750 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9624_
timestamp 0
transform 1 0 2970 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9625_
timestamp 0
transform 1 0 4230 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9626_
timestamp 0
transform -1 0 4130 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9627_
timestamp 0
transform -1 0 4510 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9628_
timestamp 0
transform 1 0 4350 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9629_
timestamp 0
transform -1 0 4590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9630_
timestamp 0
transform 1 0 3990 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9631_
timestamp 0
transform -1 0 2270 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9632_
timestamp 0
transform 1 0 1370 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9633_
timestamp 0
transform 1 0 1490 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9634_
timestamp 0
transform -1 0 1650 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9635_
timestamp 0
transform -1 0 2030 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9636_
timestamp 0
transform 1 0 2190 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9637_
timestamp 0
transform -1 0 2150 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9638_
timestamp 0
transform 1 0 2310 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9639_
timestamp 0
transform 1 0 4110 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9640_
timestamp 0
transform 1 0 4110 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9641_
timestamp 0
transform -1 0 4270 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9642_
timestamp 0
transform 1 0 3890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9643_
timestamp 0
transform -1 0 1330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9644_
timestamp 0
transform 1 0 1610 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9645_
timestamp 0
transform 1 0 1930 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9646_
timestamp 0
transform 1 0 2790 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9647_
timestamp 0
transform 1 0 1930 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9648_
timestamp 0
transform 1 0 2650 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9649_
timestamp 0
transform -1 0 2610 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9650_
timestamp 0
transform -1 0 2870 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9651_
timestamp 0
transform 1 0 3090 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9652_
timestamp 0
transform -1 0 3430 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9653_
timestamp 0
transform -1 0 3270 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9654_
timestamp 0
transform -1 0 3290 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9655_
timestamp 0
transform -1 0 3250 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9656_
timestamp 0
transform -1 0 3410 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9657_
timestamp 0
transform 1 0 3510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9658_
timestamp 0
transform -1 0 2930 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9659_
timestamp 0
transform 1 0 2090 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9660_
timestamp 0
transform -1 0 1970 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9661_
timestamp 0
transform -1 0 2370 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9662_
timestamp 0
transform -1 0 2830 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9663_
timestamp 0
transform 1 0 2970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9664_
timestamp 0
transform -1 0 3130 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9665_
timestamp 0
transform -1 0 3610 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9666_
timestamp 0
transform -1 0 2550 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9667_
timestamp 0
transform 1 0 2370 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9668_
timestamp 0
transform 1 0 2550 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9669_
timestamp 0
transform -1 0 2690 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9670_
timestamp 0
transform 1 0 2650 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9671_
timestamp 0
transform -1 0 2790 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9672_
timestamp 0
transform 1 0 2630 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9673_
timestamp 0
transform 1 0 2890 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9674_
timestamp 0
transform 1 0 3150 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9675_
timestamp 0
transform 1 0 3310 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9676_
timestamp 0
transform 1 0 3450 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9677_
timestamp 0
transform -1 0 4150 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9678_
timestamp 0
transform -1 0 3030 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9679_
timestamp 0
transform 1 0 3970 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9680_
timestamp 0
transform -1 0 2990 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9681_
timestamp 0
transform -1 0 3590 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9682_
timestamp 0
transform -1 0 2850 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9683_
timestamp 0
transform -1 0 170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9684_
timestamp 0
transform -1 0 270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9685_
timestamp 0
transform -1 0 30 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9686_
timestamp 0
transform -1 0 30 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9687_
timestamp 0
transform -1 0 190 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9688_
timestamp 0
transform -1 0 430 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9689_
timestamp 0
transform 1 0 670 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9690_
timestamp 0
transform -1 0 850 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9691_
timestamp 0
transform -1 0 30 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9692_
timestamp 0
transform -1 0 430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9693_
timestamp 0
transform -1 0 290 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9694_
timestamp 0
transform 1 0 4330 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9695_
timestamp 0
transform -1 0 30 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9696_
timestamp 0
transform -1 0 30 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9697_
timestamp 0
transform -1 0 150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9698_
timestamp 0
transform -1 0 270 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9699_
timestamp 0
transform -1 0 3650 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9700_
timestamp 0
transform 1 0 1390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9701_
timestamp 0
transform 1 0 1230 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9702_
timestamp 0
transform 1 0 1330 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9703_
timestamp 0
transform -1 0 1750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9704_
timestamp 0
transform 1 0 1130 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9705_
timestamp 0
transform 1 0 970 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9706_
timestamp 0
transform -1 0 670 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9707_
timestamp 0
transform 1 0 370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9708_
timestamp 0
transform -1 0 1810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9709_
timestamp 0
transform -1 0 1670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9710_
timestamp 0
transform -1 0 890 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9711_
timestamp 0
transform -1 0 1030 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9712_
timestamp 0
transform -1 0 2870 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9713_
timestamp 0
transform -1 0 2910 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9714_
timestamp 0
transform -1 0 270 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9715_
timestamp 0
transform -1 0 270 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9716_
timestamp 0
transform -1 0 2330 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9717_
timestamp 0
transform 1 0 1990 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9718_
timestamp 0
transform -1 0 1870 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9719_
timestamp 0
transform -1 0 3350 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9720_
timestamp 0
transform 1 0 3570 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9721_
timestamp 0
transform 1 0 3430 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9722_
timestamp 0
transform 1 0 2310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9723_
timestamp 0
transform 1 0 2170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9724_
timestamp 0
transform -1 0 3010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9725_
timestamp 0
transform -1 0 3150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9726_
timestamp 0
transform 1 0 2970 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9727_
timestamp 0
transform -1 0 3390 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9728_
timestamp 0
transform -1 0 2090 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9729_
timestamp 0
transform -1 0 2430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9730_
timestamp 0
transform 1 0 2170 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9731_
timestamp 0
transform 1 0 2030 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9732_
timestamp 0
transform -1 0 2810 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9733_
timestamp 0
transform -1 0 3210 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9734_
timestamp 0
transform -1 0 2470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9735_
timestamp 0
transform 1 0 2590 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9736_
timestamp 0
transform -1 0 810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9737_
timestamp 0
transform -1 0 950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9738_
timestamp 0
transform -1 0 2250 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9739_
timestamp 0
transform -1 0 2490 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9740_
timestamp 0
transform 1 0 1230 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9741_
timestamp 0
transform 1 0 1070 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9742_
timestamp 0
transform -1 0 1810 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9743_
timestamp 0
transform 1 0 1630 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9744_
timestamp 0
transform -1 0 1810 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9745_
timestamp 0
transform 1 0 1250 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9746_
timestamp 0
transform 1 0 2070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9747_
timestamp 0
transform -1 0 2250 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9748_
timestamp 0
transform -1 0 2290 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9749_
timestamp 0
transform 1 0 2130 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9750_
timestamp 0
transform 1 0 2570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9751_
timestamp 0
transform 1 0 2410 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9752_
timestamp 0
transform -1 0 2550 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9753_
timestamp 0
transform -1 0 2670 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9754_
timestamp 0
transform 1 0 3090 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9755_
timestamp 0
transform 1 0 2930 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9756_
timestamp 0
transform 1 0 1290 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9757_
timestamp 0
transform -1 0 1690 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9758_
timestamp 0
transform -1 0 1010 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9759_
timestamp 0
transform -1 0 1170 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9760_
timestamp 0
transform 1 0 1790 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9761_
timestamp 0
transform 1 0 1650 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9762_
timestamp 0
transform 1 0 1110 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9763_
timestamp 0
transform -1 0 970 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9844_
timestamp 0
transform 1 0 9450 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9845_
timestamp 0
transform 1 0 9790 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9846_
timestamp 0
transform 1 0 11230 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9847_
timestamp 0
transform 1 0 9910 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9848_
timestamp 0
transform 1 0 11650 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__9849_
timestamp 0
transform 1 0 11830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9850_
timestamp 0
transform -1 0 10770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9851_
timestamp 0
transform -1 0 10970 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9852_
timestamp 0
transform 1 0 10490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9853_
timestamp 0
transform 1 0 10610 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9854_
timestamp 0
transform -1 0 10650 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9855_
timestamp 0
transform -1 0 10830 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9856_
timestamp 0
transform -1 0 9770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9857_
timestamp 0
transform 1 0 9830 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9858_
timestamp 0
transform -1 0 9030 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9859_
timestamp 0
transform 1 0 11650 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__9860_
timestamp 0
transform -1 0 11790 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__9861_
timestamp 0
transform -1 0 11530 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__9862_
timestamp 0
transform -1 0 10430 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__9863_
timestamp 0
transform 1 0 9830 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9864_
timestamp 0
transform -1 0 10370 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__9865_
timestamp 0
transform -1 0 10210 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__9866_
timestamp 0
transform 1 0 9390 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9867_
timestamp 0
transform -1 0 9250 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__9868_
timestamp 0
transform -1 0 14130 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9869_
timestamp 0
transform -1 0 12570 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9870_
timestamp 0
transform -1 0 12570 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9871_
timestamp 0
transform -1 0 13610 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9872_
timestamp 0
transform -1 0 12850 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9873_
timestamp 0
transform 1 0 12690 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9874_
timestamp 0
transform -1 0 12410 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9875_
timestamp 0
transform -1 0 12170 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9876_
timestamp 0
transform -1 0 12150 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9877_
timestamp 0
transform -1 0 13190 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__9878_
timestamp 0
transform -1 0 12890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__9879_
timestamp 0
transform -1 0 13050 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__9880_
timestamp 0
transform -1 0 12970 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__9881_
timestamp 0
transform -1 0 12870 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9882_
timestamp 0
transform 1 0 12710 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__9883_
timestamp 0
transform -1 0 12730 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__9884_
timestamp 0
transform 1 0 12310 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9885_
timestamp 0
transform 1 0 12570 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__9886_
timestamp 0
transform 1 0 13550 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__9887_
timestamp 0
transform -1 0 12210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9888_
timestamp 0
transform -1 0 12150 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9889_
timestamp 0
transform 1 0 12290 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__9890_
timestamp 0
transform -1 0 11210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9891_
timestamp 0
transform -1 0 11350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9892_
timestamp 0
transform -1 0 11070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9893_
timestamp 0
transform -1 0 10870 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9894_
timestamp 0
transform -1 0 10750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9895_
timestamp 0
transform 1 0 11850 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9896_
timestamp 0
transform -1 0 11570 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9897_
timestamp 0
transform -1 0 11690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9898_
timestamp 0
transform 1 0 11250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9899_
timestamp 0
transform -1 0 11430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9900_
timestamp 0
transform 1 0 10410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9901_
timestamp 0
transform -1 0 10290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9902_
timestamp 0
transform -1 0 12490 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9903_
timestamp 0
transform 1 0 12910 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9904_
timestamp 0
transform 1 0 14990 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9905_
timestamp 0
transform 1 0 15490 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9906_
timestamp 0
transform 1 0 14990 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9907_
timestamp 0
transform -1 0 14730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9908_
timestamp 0
transform -1 0 14870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__9909_
timestamp 0
transform -1 0 13330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9910_
timestamp 0
transform -1 0 14130 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9911_
timestamp 0
transform 1 0 13970 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9912_
timestamp 0
transform -1 0 13950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9913_
timestamp 0
transform -1 0 13370 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9914_
timestamp 0
transform -1 0 13090 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9915_
timestamp 0
transform -1 0 13230 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9916_
timestamp 0
transform -1 0 12550 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9917_
timestamp 0
transform 1 0 13770 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9918_
timestamp 0
transform 1 0 13630 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9919_
timestamp 0
transform 1 0 13450 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9920_
timestamp 0
transform -1 0 13470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9921_
timestamp 0
transform 1 0 12530 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9922_
timestamp 0
transform 1 0 13010 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9923_
timestamp 0
transform -1 0 12830 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9924_
timestamp 0
transform 1 0 12610 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9925_
timestamp 0
transform -1 0 12310 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__9926_
timestamp 0
transform -1 0 12350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9927_
timestamp 0
transform 1 0 12670 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9928_
timestamp 0
transform 1 0 12670 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9929_
timestamp 0
transform -1 0 10910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9930_
timestamp 0
transform -1 0 12190 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9931_
timestamp 0
transform -1 0 13890 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9932_
timestamp 0
transform 1 0 14290 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9933_
timestamp 0
transform 1 0 13670 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9934_
timestamp 0
transform -1 0 14390 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9935_
timestamp 0
transform -1 0 11570 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9936_
timestamp 0
transform -1 0 12770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9937_
timestamp 0
transform 1 0 13030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9938_
timestamp 0
transform 1 0 12590 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9939_
timestamp 0
transform -1 0 13910 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9940_
timestamp 0
transform -1 0 12890 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9941_
timestamp 0
transform 1 0 13170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9942_
timestamp 0
transform 1 0 13770 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__9943_
timestamp 0
transform 1 0 14810 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9944_
timestamp 0
transform 1 0 15770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__9945_
timestamp 0
transform -1 0 15910 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9946_
timestamp 0
transform 1 0 15750 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__9947_
timestamp 0
transform -1 0 13730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__9948_
timestamp 0
transform 1 0 14430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9949_
timestamp 0
transform 1 0 14290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9950_
timestamp 0
transform -1 0 14130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9951_
timestamp 0
transform -1 0 13570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9952_
timestamp 0
transform 1 0 13790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9953_
timestamp 0
transform 1 0 13650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__9954_
timestamp 0
transform -1 0 13670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9955_
timestamp 0
transform -1 0 13070 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9956_
timestamp 0
transform -1 0 13210 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9957_
timestamp 0
transform -1 0 13510 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9958_
timestamp 0
transform -1 0 13350 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9959_
timestamp 0
transform 1 0 13190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9960_
timestamp 0
transform 1 0 14450 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9961_
timestamp 0
transform 1 0 13850 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9962_
timestamp 0
transform -1 0 14630 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9963_
timestamp 0
transform 1 0 14290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9964_
timestamp 0
transform 1 0 14110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9965_
timestamp 0
transform 1 0 14450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9966_
timestamp 0
transform 1 0 14610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__9967_
timestamp 0
transform 1 0 13790 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9968_
timestamp 0
transform 1 0 13650 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9969_
timestamp 0
transform -1 0 13590 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9970_
timestamp 0
transform 1 0 13510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9971_
timestamp 0
transform -1 0 13430 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9972_
timestamp 0
transform 1 0 13130 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9973_
timestamp 0
transform -1 0 13290 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9974_
timestamp 0
transform 1 0 13270 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9975_
timestamp 0
transform 1 0 12290 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9976_
timestamp 0
transform 1 0 7690 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__9977_
timestamp 0
transform -1 0 8190 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__9978_
timestamp 0
transform 1 0 7650 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__9979_
timestamp 0
transform 1 0 12830 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__9980_
timestamp 0
transform 1 0 13690 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9981_
timestamp 0
transform -1 0 15330 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__9982_
timestamp 0
transform 1 0 15150 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9983_
timestamp 0
transform 1 0 14190 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9984_
timestamp 0
transform -1 0 13890 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__9985_
timestamp 0
transform 1 0 14030 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9986_
timestamp 0
transform -1 0 14550 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__9987_
timestamp 0
transform -1 0 14170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9988_
timestamp 0
transform 1 0 14130 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9989_
timestamp 0
transform -1 0 14070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9990_
timestamp 0
transform 1 0 13350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9991_
timestamp 0
transform -1 0 13950 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__9992_
timestamp 0
transform -1 0 13850 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9993_
timestamp 0
transform 1 0 13970 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__9994_
timestamp 0
transform 1 0 14570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9995_
timestamp 0
transform -1 0 14130 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9996_
timestamp 0
transform 1 0 13990 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9997_
timestamp 0
transform -1 0 13890 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9998_
timestamp 0
transform -1 0 14290 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__9999_
timestamp 0
transform -1 0 13750 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10000_
timestamp 0
transform 1 0 13270 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10001_
timestamp 0
transform -1 0 13590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10002_
timestamp 0
transform -1 0 13450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10003_
timestamp 0
transform -1 0 13210 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10004_
timestamp 0
transform 1 0 13710 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10005_
timestamp 0
transform 1 0 14410 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10006_
timestamp 0
transform -1 0 14130 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10007_
timestamp 0
transform -1 0 14590 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10008_
timestamp 0
transform 1 0 14290 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10009_
timestamp 0
transform 1 0 16170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10010_
timestamp 0
transform 1 0 16410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10011_
timestamp 0
transform 1 0 16270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10012_
timestamp 0
transform -1 0 15210 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10013_
timestamp 0
transform -1 0 15690 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10014_
timestamp 0
transform -1 0 14710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10015_
timestamp 0
transform 1 0 14430 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10016_
timestamp 0
transform 1 0 14130 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10017_
timestamp 0
transform -1 0 15490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10018_
timestamp 0
transform 1 0 14790 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10019_
timestamp 0
transform -1 0 14290 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10020_
timestamp 0
transform -1 0 14690 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10021_
timestamp 0
transform 1 0 14370 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10022_
timestamp 0
transform -1 0 14690 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10023_
timestamp 0
transform 1 0 14830 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10024_
timestamp 0
transform -1 0 14370 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10025_
timestamp 0
transform -1 0 14230 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10026_
timestamp 0
transform -1 0 13990 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10027_
timestamp 0
transform -1 0 13830 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10028_
timestamp 0
transform 1 0 13550 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10029_
timestamp 0
transform 1 0 14450 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10030_
timestamp 0
transform 1 0 14930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10031_
timestamp 0
transform 1 0 16770 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10032_
timestamp 0
transform -1 0 15150 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__10033_
timestamp 0
transform 1 0 16850 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10034_
timestamp 0
transform -1 0 16010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10035_
timestamp 0
transform -1 0 16150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10036_
timestamp 0
transform -1 0 14670 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10037_
timestamp 0
transform -1 0 14810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10038_
timestamp 0
transform 1 0 15190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10039_
timestamp 0
transform -1 0 14910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10040_
timestamp 0
transform 1 0 15050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10041_
timestamp 0
transform 1 0 15070 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10042_
timestamp 0
transform 1 0 14930 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10043_
timestamp 0
transform -1 0 14990 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10044_
timestamp 0
transform -1 0 14610 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10045_
timestamp 0
transform -1 0 14470 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10046_
timestamp 0
transform 1 0 14730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10047_
timestamp 0
transform -1 0 14630 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10048_
timestamp 0
transform -1 0 14790 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10049_
timestamp 0
transform -1 0 14650 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10050_
timestamp 0
transform 1 0 13950 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10051_
timestamp 0
transform 1 0 14930 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10052_
timestamp 0
transform 1 0 15530 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10053_
timestamp 0
transform 1 0 14510 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10054_
timestamp 0
transform 1 0 16350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10055_
timestamp 0
transform -1 0 16290 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10056_
timestamp 0
transform 1 0 15970 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10057_
timestamp 0
transform -1 0 15770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10058_
timestamp 0
transform -1 0 15770 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10059_
timestamp 0
transform -1 0 15370 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10060_
timestamp 0
transform 1 0 15290 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10061_
timestamp 0
transform 1 0 15670 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10062_
timestamp 0
transform -1 0 15550 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10063_
timestamp 0
transform -1 0 15410 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10064_
timestamp 0
transform -1 0 15270 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10065_
timestamp 0
transform 1 0 15290 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10066_
timestamp 0
transform 1 0 15230 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10067_
timestamp 0
transform -1 0 14850 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__10068_
timestamp 0
transform 1 0 14950 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10069_
timestamp 0
transform -1 0 14830 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10070_
timestamp 0
transform 1 0 12990 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10071_
timestamp 0
transform 1 0 14410 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10072_
timestamp 0
transform -1 0 15570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10073_
timestamp 0
transform 1 0 15210 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10074_
timestamp 0
transform -1 0 16150 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10075_
timestamp 0
transform -1 0 15930 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10076_
timestamp 0
transform -1 0 16070 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10077_
timestamp 0
transform 1 0 15650 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10078_
timestamp 0
transform 1 0 15930 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10079_
timestamp 0
transform 1 0 15490 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10080_
timestamp 0
transform 1 0 15810 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10081_
timestamp 0
transform -1 0 15690 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10082_
timestamp 0
transform 1 0 16030 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10083_
timestamp 0
transform -1 0 15990 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10084_
timestamp 0
transform 1 0 16090 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10085_
timestamp 0
transform -1 0 15610 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10086_
timestamp 0
transform 1 0 15110 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10087_
timestamp 0
transform -1 0 15030 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10088_
timestamp 0
transform 1 0 14870 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10089_
timestamp 0
transform -1 0 15110 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10090_
timestamp 0
transform -1 0 15270 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10091_
timestamp 0
transform -1 0 15110 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10092_
timestamp 0
transform 1 0 14510 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10093_
timestamp 0
transform -1 0 13170 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10094_
timestamp 0
transform 1 0 15810 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10095_
timestamp 0
transform 1 0 14730 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10096_
timestamp 0
transform 1 0 15410 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10097_
timestamp 0
transform 1 0 15150 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10098_
timestamp 0
transform 1 0 15570 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10099_
timestamp 0
transform -1 0 15750 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10100_
timestamp 0
transform 1 0 15870 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10101_
timestamp 0
transform 1 0 15770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10102_
timestamp 0
transform 1 0 16470 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10103_
timestamp 0
transform 1 0 16470 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10104_
timestamp 0
transform 1 0 16610 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10105_
timestamp 0
transform 1 0 16190 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10106_
timestamp 0
transform -1 0 16270 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10107_
timestamp 0
transform -1 0 16070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10108_
timestamp 0
transform 1 0 16190 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10109_
timestamp 0
transform 1 0 16130 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10110_
timestamp 0
transform -1 0 15990 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10111_
timestamp 0
transform -1 0 16110 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10112_
timestamp 0
transform 1 0 16230 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10113_
timestamp 0
transform 1 0 15930 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10114_
timestamp 0
transform 1 0 15850 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10115_
timestamp 0
transform -1 0 15490 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10116_
timestamp 0
transform 1 0 15350 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10117_
timestamp 0
transform 1 0 15530 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10118_
timestamp 0
transform -1 0 15410 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10119_
timestamp 0
transform 1 0 13450 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10120_
timestamp 0
transform 1 0 13650 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10121_
timestamp 0
transform -1 0 14690 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10122_
timestamp 0
transform 1 0 13490 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10123_
timestamp 0
transform 1 0 13870 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__10124_
timestamp 0
transform 1 0 15970 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10125_
timestamp 0
transform 1 0 15690 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10126_
timestamp 0
transform 1 0 15830 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10127_
timestamp 0
transform 1 0 16470 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10128_
timestamp 0
transform 1 0 16350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10129_
timestamp 0
transform 1 0 16430 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10130_
timestamp 0
transform -1 0 16770 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10131_
timestamp 0
transform -1 0 16510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10132_
timestamp 0
transform -1 0 16910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10133_
timestamp 0
transform 1 0 16750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10134_
timestamp 0
transform 1 0 16590 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10135_
timestamp 0
transform 1 0 16890 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10136_
timestamp 0
transform -1 0 16630 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10137_
timestamp 0
transform -1 0 16830 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10138_
timestamp 0
transform 1 0 16590 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10139_
timestamp 0
transform -1 0 16430 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10140_
timestamp 0
transform -1 0 16130 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10141_
timestamp 0
transform -1 0 16270 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10142_
timestamp 0
transform 1 0 14010 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10143_
timestamp 0
transform -1 0 15890 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10144_
timestamp 0
transform -1 0 16010 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10145_
timestamp 0
transform 1 0 15710 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10146_
timestamp 0
transform 1 0 15970 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10147_
timestamp 0
transform 1 0 16130 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10148_
timestamp 0
transform 1 0 16550 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10149_
timestamp 0
transform -1 0 16430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10150_
timestamp 0
transform -1 0 16450 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__10151_
timestamp 0
transform 1 0 16410 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10152_
timestamp 0
transform 1 0 17010 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10153_
timestamp 0
transform 1 0 16590 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10154_
timestamp 0
transform 1 0 16950 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10155_
timestamp 0
transform 1 0 16910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10156_
timestamp 0
transform 1 0 16750 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10157_
timestamp 0
transform 1 0 17030 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10158_
timestamp 0
transform 1 0 16210 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__10159_
timestamp 0
transform 1 0 16650 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10160_
timestamp 0
transform 1 0 16790 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10161_
timestamp 0
transform -1 0 16690 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10162_
timestamp 0
transform -1 0 16310 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10163_
timestamp 0
transform -1 0 16270 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10164_
timestamp 0
transform -1 0 16170 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10165_
timestamp 0
transform 1 0 13290 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10166_
timestamp 0
transform 1 0 16790 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10167_
timestamp 0
transform 1 0 16330 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10168_
timestamp 0
transform -1 0 17030 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10169_
timestamp 0
transform 1 0 15690 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__10170_
timestamp 0
transform -1 0 16870 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10171_
timestamp 0
transform -1 0 16910 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10172_
timestamp 0
transform 1 0 16710 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10173_
timestamp 0
transform -1 0 16090 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__10174_
timestamp 0
transform 1 0 16990 0 1 250
box -6 -8 26 248
use FILL  FILL_0__10175_
timestamp 0
transform -1 0 17070 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__10176_
timestamp 0
transform -1 0 17030 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10177_
timestamp 0
transform 1 0 16930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10178_
timestamp 0
transform -1 0 16810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10179_
timestamp 0
transform 1 0 17010 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10180_
timestamp 0
transform -1 0 17030 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10181_
timestamp 0
transform 1 0 16970 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10182_
timestamp 0
transform 1 0 16430 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10183_
timestamp 0
transform -1 0 16890 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10184_
timestamp 0
transform -1 0 16990 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10185_
timestamp 0
transform -1 0 16750 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10186_
timestamp 0
transform 1 0 16570 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10187_
timestamp 0
transform -1 0 16430 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10188_
timestamp 0
transform -1 0 16290 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10189_
timestamp 0
transform 1 0 14450 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10190_
timestamp 0
transform -1 0 12090 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10191_
timestamp 0
transform -1 0 16870 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10192_
timestamp 0
transform 1 0 17030 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10193_
timestamp 0
transform 1 0 16790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10194_
timestamp 0
transform -1 0 16910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10195_
timestamp 0
transform 1 0 17030 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10196_
timestamp 0
transform 1 0 16710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10197_
timestamp 0
transform 1 0 15270 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__10198_
timestamp 0
transform -1 0 16850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10199_
timestamp 0
transform 1 0 16950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10200_
timestamp 0
transform 1 0 17070 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10201_
timestamp 0
transform -1 0 16850 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10202_
timestamp 0
transform 1 0 16710 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10203_
timestamp 0
transform -1 0 16690 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10204_
timestamp 0
transform -1 0 16550 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10205_
timestamp 0
transform 1 0 12430 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10206_
timestamp 0
transform -1 0 11550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10207_
timestamp 0
transform 1 0 14270 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10208_
timestamp 0
transform 1 0 14510 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10209_
timestamp 0
transform 1 0 14370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10210_
timestamp 0
transform 1 0 14130 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10211_
timestamp 0
transform -1 0 12770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10212_
timestamp 0
transform -1 0 12510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10213_
timestamp 0
transform -1 0 13030 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10214_
timestamp 0
transform -1 0 14010 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10215_
timestamp 0
transform 1 0 15730 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10216_
timestamp 0
transform 1 0 15630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10217_
timestamp 0
transform 1 0 15470 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10218_
timestamp 0
transform 1 0 15310 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10219_
timestamp 0
transform 1 0 15350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10220_
timestamp 0
transform 1 0 15350 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10221_
timestamp 0
transform 1 0 14910 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10222_
timestamp 0
transform 1 0 12950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10223_
timestamp 0
transform -1 0 15230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10224_
timestamp 0
transform 1 0 15630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10225_
timestamp 0
transform 1 0 15330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10226_
timestamp 0
transform -1 0 15090 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10227_
timestamp 0
transform 1 0 13210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10228_
timestamp 0
transform -1 0 11930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10229_
timestamp 0
transform 1 0 10790 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10230_
timestamp 0
transform 1 0 13090 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10231_
timestamp 0
transform -1 0 14850 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10232_
timestamp 0
transform 1 0 14670 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10233_
timestamp 0
transform -1 0 14170 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10234_
timestamp 0
transform -1 0 14290 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10235_
timestamp 0
transform 1 0 14910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10236_
timestamp 0
transform -1 0 15510 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10237_
timestamp 0
transform -1 0 15790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10238_
timestamp 0
transform -1 0 15930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10239_
timestamp 0
transform 1 0 15910 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10240_
timestamp 0
transform -1 0 15630 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10241_
timestamp 0
transform 1 0 15590 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10242_
timestamp 0
transform -1 0 15710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10243_
timestamp 0
transform -1 0 15790 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10244_
timestamp 0
transform -1 0 15630 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10245_
timestamp 0
transform -1 0 14250 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10246_
timestamp 0
transform -1 0 15530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10247_
timestamp 0
transform 1 0 15070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10248_
timestamp 0
transform 1 0 14550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10249_
timestamp 0
transform -1 0 12750 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10250_
timestamp 0
transform -1 0 12350 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10251_
timestamp 0
transform -1 0 12910 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10252_
timestamp 0
transform 1 0 12430 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10253_
timestamp 0
transform 1 0 12650 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10254_
timestamp 0
transform 1 0 12790 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10255_
timestamp 0
transform 1 0 12930 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10256_
timestamp 0
transform -1 0 10950 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10257_
timestamp 0
transform -1 0 11050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10258_
timestamp 0
transform 1 0 12570 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10259_
timestamp 0
transform 1 0 14510 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10260_
timestamp 0
transform 1 0 16290 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10261_
timestamp 0
transform 1 0 16150 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10262_
timestamp 0
transform -1 0 16090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10263_
timestamp 0
transform 1 0 16190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10264_
timestamp 0
transform -1 0 14710 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10265_
timestamp 0
transform -1 0 14930 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10266_
timestamp 0
transform 1 0 14790 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10267_
timestamp 0
transform -1 0 15230 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10268_
timestamp 0
transform -1 0 14510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10269_
timestamp 0
transform 1 0 14370 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10270_
timestamp 0
transform 1 0 15050 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10271_
timestamp 0
transform -1 0 14650 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10272_
timestamp 0
transform -1 0 13410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10273_
timestamp 0
transform 1 0 13150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10274_
timestamp 0
transform -1 0 13270 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10275_
timestamp 0
transform 1 0 13010 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10276_
timestamp 0
transform -1 0 12210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10277_
timestamp 0
transform 1 0 12190 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10278_
timestamp 0
transform -1 0 12070 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10279_
timestamp 0
transform -1 0 11410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10280_
timestamp 0
transform 1 0 12850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10281_
timestamp 0
transform -1 0 12850 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10282_
timestamp 0
transform 1 0 16650 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10283_
timestamp 0
transform 1 0 16510 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10284_
timestamp 0
transform 1 0 16030 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10285_
timestamp 0
transform 1 0 15710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10286_
timestamp 0
transform 1 0 14790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10287_
timestamp 0
transform -1 0 14950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10288_
timestamp 0
transform 1 0 14810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10289_
timestamp 0
transform 1 0 14750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10290_
timestamp 0
transform -1 0 14370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10291_
timestamp 0
transform -1 0 14090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10292_
timestamp 0
transform -1 0 14630 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10293_
timestamp 0
transform -1 0 13450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10294_
timestamp 0
transform -1 0 12770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10295_
timestamp 0
transform 1 0 13570 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10296_
timestamp 0
transform -1 0 12630 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10297_
timestamp 0
transform -1 0 12590 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10298_
timestamp 0
transform -1 0 12730 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10299_
timestamp 0
transform -1 0 12450 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10300_
timestamp 0
transform 1 0 11970 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10301_
timestamp 0
transform 1 0 12870 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10302_
timestamp 0
transform -1 0 16930 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10303_
timestamp 0
transform 1 0 16750 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10304_
timestamp 0
transform 1 0 16350 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10305_
timestamp 0
transform 1 0 16210 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10306_
timestamp 0
transform 1 0 15450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10307_
timestamp 0
transform 1 0 15310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10308_
timestamp 0
transform -1 0 15330 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10309_
timestamp 0
transform 1 0 14770 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10310_
timestamp 0
transform -1 0 14810 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10311_
timestamp 0
transform -1 0 14490 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10312_
timestamp 0
transform 1 0 14930 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10313_
timestamp 0
transform 1 0 15370 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10314_
timestamp 0
transform -1 0 14350 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10315_
timestamp 0
transform -1 0 14650 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10316_
timestamp 0
transform 1 0 15050 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10317_
timestamp 0
transform -1 0 13790 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10318_
timestamp 0
transform -1 0 13490 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10319_
timestamp 0
transform -1 0 13210 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10320_
timestamp 0
transform -1 0 13350 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10321_
timestamp 0
transform -1 0 13090 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10322_
timestamp 0
transform 1 0 12390 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10323_
timestamp 0
transform 1 0 12190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10324_
timestamp 0
transform 1 0 13750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10325_
timestamp 0
transform 1 0 15790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10326_
timestamp 0
transform -1 0 16010 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10327_
timestamp 0
transform 1 0 16110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10328_
timestamp 0
transform 1 0 15810 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10329_
timestamp 0
transform -1 0 15950 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10330_
timestamp 0
transform -1 0 16090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10331_
timestamp 0
transform -1 0 15950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10332_
timestamp 0
transform 1 0 14910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10333_
timestamp 0
transform 1 0 15050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10334_
timestamp 0
transform 1 0 15650 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10335_
timestamp 0
transform 1 0 15530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10336_
timestamp 0
transform -1 0 15110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10337_
timestamp 0
transform -1 0 14610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10338_
timestamp 0
transform 1 0 15230 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10339_
timestamp 0
transform -1 0 13910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10340_
timestamp 0
transform 1 0 13630 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10341_
timestamp 0
transform -1 0 13490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10342_
timestamp 0
transform -1 0 13350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10343_
timestamp 0
transform 1 0 12290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10344_
timestamp 0
transform 1 0 11330 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10345_
timestamp 0
transform -1 0 15670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10346_
timestamp 0
transform 1 0 16270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10347_
timestamp 0
transform 1 0 16470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10348_
timestamp 0
transform 1 0 16330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10349_
timestamp 0
transform 1 0 15130 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10350_
timestamp 0
transform -1 0 15450 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10351_
timestamp 0
transform 1 0 15570 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10352_
timestamp 0
transform 1 0 15290 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10353_
timestamp 0
transform 1 0 14990 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10354_
timestamp 0
transform 1 0 14730 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10355_
timestamp 0
transform -1 0 14870 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10356_
timestamp 0
transform -1 0 14470 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10357_
timestamp 0
transform 1 0 13910 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10358_
timestamp 0
transform 1 0 14190 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10359_
timestamp 0
transform 1 0 14050 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10360_
timestamp 0
transform -1 0 14190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10361_
timestamp 0
transform -1 0 14210 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10362_
timestamp 0
transform -1 0 14610 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10363_
timestamp 0
transform -1 0 13630 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10364_
timestamp 0
transform 1 0 14030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10365_
timestamp 0
transform 1 0 14430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10366_
timestamp 0
transform 1 0 14290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10367_
timestamp 0
transform -1 0 14350 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10368_
timestamp 0
transform -1 0 13830 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10369_
timestamp 0
transform 1 0 12890 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10370_
timestamp 0
transform 1 0 11450 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10371_
timestamp 0
transform 1 0 12790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10372_
timestamp 0
transform -1 0 13990 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10373_
timestamp 0
transform 1 0 15210 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10374_
timestamp 0
transform 1 0 16310 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10375_
timestamp 0
transform 1 0 16430 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10376_
timestamp 0
transform 1 0 16190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10377_
timestamp 0
transform -1 0 14830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10378_
timestamp 0
transform -1 0 15130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10379_
timestamp 0
transform 1 0 15430 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10380_
timestamp 0
transform -1 0 14990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10381_
timestamp 0
transform -1 0 14690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10382_
timestamp 0
transform 1 0 15470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10383_
timestamp 0
transform 1 0 15470 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__10384_
timestamp 0
transform -1 0 15610 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__10385_
timestamp 0
transform 1 0 15190 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__10386_
timestamp 0
transform 1 0 13410 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10387_
timestamp 0
transform -1 0 13290 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10388_
timestamp 0
transform -1 0 13190 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10389_
timestamp 0
transform -1 0 13030 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10390_
timestamp 0
transform 1 0 12890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10391_
timestamp 0
transform 1 0 14530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10392_
timestamp 0
transform -1 0 14270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10393_
timestamp 0
transform 1 0 14390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10394_
timestamp 0
transform 1 0 16110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__10395_
timestamp 0
transform -1 0 15350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10396_
timestamp 0
transform -1 0 16210 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10397_
timestamp 0
transform 1 0 16250 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10398_
timestamp 0
transform 1 0 16570 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__10399_
timestamp 0
transform -1 0 16530 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__10400_
timestamp 0
transform 1 0 15630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10401_
timestamp 0
transform -1 0 16250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__10402_
timestamp 0
transform 1 0 16370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__10403_
timestamp 0
transform -1 0 16690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__10404_
timestamp 0
transform 1 0 16170 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__10405_
timestamp 0
transform -1 0 16050 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__10406_
timestamp 0
transform -1 0 14110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10407_
timestamp 0
transform -1 0 14110 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10408_
timestamp 0
transform -1 0 15330 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__10409_
timestamp 0
transform -1 0 13710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10410_
timestamp 0
transform 1 0 13650 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10411_
timestamp 0
transform 1 0 12750 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10412_
timestamp 0
transform -1 0 13850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10413_
timestamp 0
transform -1 0 13970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10414_
timestamp 0
transform 1 0 16950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10415_
timestamp 0
transform 1 0 16890 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__10416_
timestamp 0
transform -1 0 16850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__10417_
timestamp 0
transform 1 0 16970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__10418_
timestamp 0
transform 1 0 15390 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__10419_
timestamp 0
transform 1 0 16910 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__10420_
timestamp 0
transform 1 0 16910 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__10421_
timestamp 0
transform 1 0 16670 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__10422_
timestamp 0
transform -1 0 16070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10423_
timestamp 0
transform -1 0 13310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10424_
timestamp 0
transform -1 0 13170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10425_
timestamp 0
transform -1 0 13010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10426_
timestamp 0
transform 1 0 13050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10427_
timestamp 0
transform 1 0 16790 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__10428_
timestamp 0
transform -1 0 15930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10429_
timestamp 0
transform -1 0 16310 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__10430_
timestamp 0
transform -1 0 16430 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__10431_
timestamp 0
transform 1 0 15770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10432_
timestamp 0
transform -1 0 16310 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__10433_
timestamp 0
transform 1 0 16370 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__10434_
timestamp 0
transform 1 0 16550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10435_
timestamp 0
transform -1 0 16890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10436_
timestamp 0
transform 1 0 16830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10437_
timestamp 0
transform -1 0 16730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10438_
timestamp 0
transform -1 0 16650 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10439_
timestamp 0
transform 1 0 17010 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10440_
timestamp 0
transform -1 0 17030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__10441_
timestamp 0
transform -1 0 16890 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10442_
timestamp 0
transform 1 0 16490 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10443_
timestamp 0
transform 1 0 15950 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10444_
timestamp 0
transform -1 0 15830 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10445_
timestamp 0
transform -1 0 15710 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10446_
timestamp 0
transform 1 0 13150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__10447_
timestamp 0
transform 1 0 12070 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10448_
timestamp 0
transform 1 0 16390 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10449_
timestamp 0
transform 1 0 16090 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__10450_
timestamp 0
transform 1 0 16670 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10451_
timestamp 0
transform 1 0 16610 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10452_
timestamp 0
transform 1 0 16570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10453_
timestamp 0
transform 1 0 16470 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10454_
timestamp 0
transform -1 0 13190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10455_
timestamp 0
transform -1 0 13050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10456_
timestamp 0
transform -1 0 12470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10457_
timestamp 0
transform 1 0 11150 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10458_
timestamp 0
transform -1 0 9390 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10459_
timestamp 0
transform -1 0 9290 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10460_
timestamp 0
transform 1 0 9670 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10461_
timestamp 0
transform 1 0 9530 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10462_
timestamp 0
transform 1 0 9710 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10463_
timestamp 0
transform 1 0 9950 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10464_
timestamp 0
transform 1 0 9810 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10465_
timestamp 0
transform 1 0 9250 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10466_
timestamp 0
transform -1 0 9110 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10467_
timestamp 0
transform 1 0 10570 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10468_
timestamp 0
transform -1 0 9950 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10469_
timestamp 0
transform -1 0 9830 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10470_
timestamp 0
transform 1 0 9930 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10471_
timestamp 0
transform -1 0 9810 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10472_
timestamp 0
transform -1 0 8890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10473_
timestamp 0
transform -1 0 8630 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10474_
timestamp 0
transform -1 0 8750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10475_
timestamp 0
transform -1 0 8610 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10476_
timestamp 0
transform -1 0 8770 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10477_
timestamp 0
transform -1 0 8850 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10478_
timestamp 0
transform -1 0 8990 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10479_
timestamp 0
transform 1 0 8870 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10480_
timestamp 0
transform 1 0 8770 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10481_
timestamp 0
transform 1 0 8890 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10482_
timestamp 0
transform -1 0 11090 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10483_
timestamp 0
transform -1 0 10230 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10484_
timestamp 0
transform -1 0 10370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10485_
timestamp 0
transform 1 0 9330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10486_
timestamp 0
transform -1 0 9210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10487_
timestamp 0
transform 1 0 9050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10488_
timestamp 0
transform -1 0 8970 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10489_
timestamp 0
transform -1 0 8710 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10490_
timestamp 0
transform -1 0 8850 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10491_
timestamp 0
transform 1 0 9730 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10492_
timestamp 0
transform 1 0 9550 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10493_
timestamp 0
transform -1 0 9490 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10494_
timestamp 0
transform 1 0 9850 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10495_
timestamp 0
transform 1 0 9990 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10496_
timestamp 0
transform 1 0 10230 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10497_
timestamp 0
transform 1 0 11290 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10498_
timestamp 0
transform -1 0 11170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10499_
timestamp 0
transform 1 0 10990 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10500_
timestamp 0
transform -1 0 11030 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10501_
timestamp 0
transform 1 0 10470 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10502_
timestamp 0
transform 1 0 10350 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10503_
timestamp 0
transform -1 0 9610 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10504_
timestamp 0
transform -1 0 9470 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10505_
timestamp 0
transform -1 0 9170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10506_
timestamp 0
transform 1 0 9290 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10507_
timestamp 0
transform 1 0 9590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10508_
timestamp 0
transform 1 0 10970 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__10509_
timestamp 0
transform -1 0 10570 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10510_
timestamp 0
transform -1 0 10870 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10511_
timestamp 0
transform 1 0 10690 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10512_
timestamp 0
transform 1 0 10090 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10513_
timestamp 0
transform 1 0 10470 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10514_
timestamp 0
transform -1 0 10370 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10515_
timestamp 0
transform 1 0 10430 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__10516_
timestamp 0
transform 1 0 10090 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10517_
timestamp 0
transform 1 0 10690 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__10518_
timestamp 0
transform 1 0 10950 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__10519_
timestamp 0
transform -1 0 10850 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__10520_
timestamp 0
transform -1 0 10810 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__10521_
timestamp 0
transform -1 0 11170 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10522_
timestamp 0
transform -1 0 12890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10523_
timestamp 0
transform 1 0 13110 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10524_
timestamp 0
transform -1 0 12990 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10525_
timestamp 0
transform -1 0 12850 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10526_
timestamp 0
transform -1 0 10930 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10527_
timestamp 0
transform -1 0 11070 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10528_
timestamp 0
transform -1 0 10810 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10529_
timestamp 0
transform -1 0 10550 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10530_
timestamp 0
transform 1 0 10950 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__10531_
timestamp 0
transform 1 0 10830 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__10532_
timestamp 0
transform 1 0 10690 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__10533_
timestamp 0
transform 1 0 10530 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__10534_
timestamp 0
transform -1 0 9450 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10535_
timestamp 0
transform 1 0 10570 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__10536_
timestamp 0
transform -1 0 10690 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__10537_
timestamp 0
transform 1 0 10630 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10538_
timestamp 0
transform 1 0 10330 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__10539_
timestamp 0
transform -1 0 10530 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__10540_
timestamp 0
transform -1 0 11430 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10541_
timestamp 0
transform 1 0 10890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10542_
timestamp 0
transform -1 0 10490 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10543_
timestamp 0
transform -1 0 10770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10544_
timestamp 0
transform -1 0 10630 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10545_
timestamp 0
transform 1 0 10830 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10546_
timestamp 0
transform 1 0 10950 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10547_
timestamp 0
transform 1 0 10430 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10548_
timestamp 0
transform -1 0 10110 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__10549_
timestamp 0
transform -1 0 9850 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__10550_
timestamp 0
transform -1 0 9990 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__10551_
timestamp 0
transform 1 0 9690 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10552_
timestamp 0
transform -1 0 9570 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10553_
timestamp 0
transform -1 0 9250 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10554_
timestamp 0
transform -1 0 9810 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10555_
timestamp 0
transform 1 0 10230 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10556_
timestamp 0
transform 1 0 10690 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10557_
timestamp 0
transform -1 0 10570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10558_
timestamp 0
transform -1 0 10430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10559_
timestamp 0
transform -1 0 10170 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10560_
timestamp 0
transform -1 0 10110 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10561_
timestamp 0
transform 1 0 10270 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10562_
timestamp 0
transform -1 0 10250 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10563_
timestamp 0
transform -1 0 9510 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10564_
timestamp 0
transform -1 0 9670 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10565_
timestamp 0
transform 1 0 9330 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10566_
timestamp 0
transform 1 0 11110 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__10567_
timestamp 0
transform -1 0 11310 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10568_
timestamp 0
transform 1 0 11410 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10569_
timestamp 0
transform -1 0 11410 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10570_
timestamp 0
transform -1 0 11110 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10571_
timestamp 0
transform 1 0 11530 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10572_
timestamp 0
transform -1 0 11210 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10573_
timestamp 0
transform 1 0 10070 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10574_
timestamp 0
transform 1 0 9950 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10575_
timestamp 0
transform 1 0 10070 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10576_
timestamp 0
transform -1 0 10410 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10577_
timestamp 0
transform -1 0 10250 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10578_
timestamp 0
transform 1 0 11390 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__10579_
timestamp 0
transform 1 0 11510 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__10580_
timestamp 0
transform 1 0 11630 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__10581_
timestamp 0
transform -1 0 11270 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__10582_
timestamp 0
transform 1 0 11350 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__10583_
timestamp 0
transform 1 0 11490 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10584_
timestamp 0
transform 1 0 11630 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10585_
timestamp 0
transform -1 0 11610 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10586_
timestamp 0
transform -1 0 11350 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__10587_
timestamp 0
transform 1 0 11630 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__10588_
timestamp 0
transform -1 0 11490 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__10589_
timestamp 0
transform -1 0 11790 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__10590_
timestamp 0
transform -1 0 11330 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10591_
timestamp 0
transform -1 0 11470 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10592_
timestamp 0
transform -1 0 11230 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10593_
timestamp 0
transform 1 0 11330 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10594_
timestamp 0
transform -1 0 11850 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10595_
timestamp 0
transform -1 0 12030 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10596_
timestamp 0
transform 1 0 11870 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__10597_
timestamp 0
transform -1 0 11970 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__10598_
timestamp 0
transform 1 0 12450 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__10599_
timestamp 0
transform -1 0 12310 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__10600_
timestamp 0
transform -1 0 12170 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__10601_
timestamp 0
transform -1 0 11930 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__10602_
timestamp 0
transform -1 0 12210 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__10603_
timestamp 0
transform -1 0 12070 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__10604_
timestamp 0
transform 1 0 10430 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10605_
timestamp 0
transform -1 0 11250 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10606_
timestamp 0
transform 1 0 10570 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10607_
timestamp 0
transform 1 0 15190 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10608_
timestamp 0
transform -1 0 16570 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10609_
timestamp 0
transform -1 0 16090 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10610_
timestamp 0
transform 1 0 16710 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__10611_
timestamp 0
transform 1 0 11550 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10612_
timestamp 0
transform 1 0 10710 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10613_
timestamp 0
transform 1 0 11250 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10614_
timestamp 0
transform -1 0 11430 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10615_
timestamp 0
transform -1 0 11170 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10616_
timestamp 0
transform 1 0 10850 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10617_
timestamp 0
transform -1 0 11030 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10618_
timestamp 0
transform -1 0 10610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10619_
timestamp 0
transform -1 0 12750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10620_
timestamp 0
transform 1 0 12570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10621_
timestamp 0
transform 1 0 11950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__10622_
timestamp 0
transform 1 0 11910 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__10623_
timestamp 0
transform 1 0 10110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10624_
timestamp 0
transform 1 0 13570 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10625_
timestamp 0
transform 1 0 13410 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10626_
timestamp 0
transform -1 0 13710 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10627_
timestamp 0
transform -1 0 13830 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__10628_
timestamp 0
transform 1 0 12390 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10629_
timestamp 0
transform 1 0 12050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10630_
timestamp 0
transform -1 0 12250 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10631_
timestamp 0
transform 1 0 11850 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10632_
timestamp 0
transform 1 0 12430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10633_
timestamp 0
transform -1 0 12590 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10634_
timestamp 0
transform -1 0 13390 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10635_
timestamp 0
transform 1 0 13490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10636_
timestamp 0
transform 1 0 16270 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10637_
timestamp 0
transform -1 0 16410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__10638_
timestamp 0
transform 1 0 15190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10639_
timestamp 0
transform -1 0 15850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__10640_
timestamp 0
transform -1 0 11830 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10641_
timestamp 0
transform -1 0 12090 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10642_
timestamp 0
transform 1 0 11910 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10643_
timestamp 0
transform -1 0 11970 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10644_
timestamp 0
transform 1 0 12350 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10645_
timestamp 0
transform 1 0 12210 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10646_
timestamp 0
transform -1 0 12390 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10647_
timestamp 0
transform 1 0 11970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10648_
timestamp 0
transform -1 0 12930 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10649_
timestamp 0
transform 1 0 12750 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10650_
timestamp 0
transform 1 0 15350 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10651_
timestamp 0
transform 1 0 15190 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10652_
timestamp 0
transform -1 0 15050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10653_
timestamp 0
transform -1 0 15170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10654_
timestamp 0
transform -1 0 11690 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10655_
timestamp 0
transform -1 0 11690 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10656_
timestamp 0
transform 1 0 12190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10657_
timestamp 0
transform 1 0 12050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10658_
timestamp 0
transform -1 0 11850 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10659_
timestamp 0
transform -1 0 12170 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__10660_
timestamp 0
transform -1 0 13350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10661_
timestamp 0
transform -1 0 13390 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10662_
timestamp 0
transform 1 0 11750 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10663_
timestamp 0
transform -1 0 11890 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10664_
timestamp 0
transform 1 0 11670 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10665_
timestamp 0
transform -1 0 11810 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10666_
timestamp 0
transform -1 0 9710 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10667_
timestamp 0
transform -1 0 11550 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10668_
timestamp 0
transform 1 0 11130 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10669_
timestamp 0
transform -1 0 10110 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10670_
timestamp 0
transform -1 0 10930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10671_
timestamp 0
transform 1 0 10770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10672_
timestamp 0
transform -1 0 10630 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10673_
timestamp 0
transform -1 0 10750 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__10674_
timestamp 0
transform -1 0 10210 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10675_
timestamp 0
transform -1 0 10330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__10676_
timestamp 0
transform 1 0 11030 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10677_
timestamp 0
transform 1 0 10890 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__10678_
timestamp 0
transform 1 0 11110 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10679_
timestamp 0
transform 1 0 11250 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10680_
timestamp 0
transform -1 0 9650 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10681_
timestamp 0
transform -1 0 9710 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10682_
timestamp 0
transform -1 0 10050 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__10683_
timestamp 0
transform -1 0 10090 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__10684_
timestamp 0
transform 1 0 9350 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10685_
timestamp 0
transform 1 0 9190 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10686_
timestamp 0
transform -1 0 8570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10687_
timestamp 0
transform -1 0 8690 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__10768_
timestamp 0
transform -1 0 5650 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__10769_
timestamp 0
transform -1 0 4830 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__10770_
timestamp 0
transform -1 0 4730 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__10771_
timestamp 0
transform -1 0 5510 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__10772_
timestamp 0
transform 1 0 5610 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__10773_
timestamp 0
transform -1 0 4350 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__10774_
timestamp 0
transform 1 0 5530 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__10775_
timestamp 0
transform 1 0 5550 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__10776_
timestamp 0
transform -1 0 2670 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__10777_
timestamp 0
transform 1 0 5410 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__10778_
timestamp 0
transform 1 0 5910 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__10779_
timestamp 0
transform 1 0 5750 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__10780_
timestamp 0
transform -1 0 4530 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__10781_
timestamp 0
transform -1 0 5790 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__10782_
timestamp 0
transform 1 0 5430 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__10783_
timestamp 0
transform 1 0 5090 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__10784_
timestamp 0
transform 1 0 5310 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__10785_
timestamp 0
transform 1 0 5470 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__10786_
timestamp 0
transform -1 0 6730 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__10787_
timestamp 0
transform -1 0 5590 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__10788_
timestamp 0
transform -1 0 6090 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__10789_
timestamp 0
transform 1 0 6230 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__10790_
timestamp 0
transform 1 0 6450 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__10791_
timestamp 0
transform 1 0 6610 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__10792_
timestamp 0
transform -1 0 5890 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10793_
timestamp 0
transform -1 0 5290 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__10794_
timestamp 0
transform 1 0 5430 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__10795_
timestamp 0
transform 1 0 5810 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10796_
timestamp 0
transform 1 0 6130 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__10797_
timestamp 0
transform 1 0 5990 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__10798_
timestamp 0
transform 1 0 5570 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__10799_
timestamp 0
transform 1 0 5110 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__10800_
timestamp 0
transform 1 0 6290 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__10801_
timestamp 0
transform -1 0 5610 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__10802_
timestamp 0
transform -1 0 5610 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__10803_
timestamp 0
transform 1 0 5730 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__10804_
timestamp 0
transform -1 0 5330 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__10805_
timestamp 0
transform 1 0 5730 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__10806_
timestamp 0
transform 1 0 5870 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__10807_
timestamp 0
transform 1 0 5890 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__10808_
timestamp 0
transform 1 0 5070 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__10809_
timestamp 0
transform 1 0 6170 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__10810_
timestamp 0
transform 1 0 1070 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__10811_
timestamp 0
transform 1 0 1910 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__10812_
timestamp 0
transform 1 0 1210 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__10813_
timestamp 0
transform 1 0 1530 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__10814_
timestamp 0
transform 1 0 1530 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__10815_
timestamp 0
transform -1 0 1390 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__10816_
timestamp 0
transform 1 0 1650 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__10817_
timestamp 0
transform 1 0 2750 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__10818_
timestamp 0
transform -1 0 2270 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__10819_
timestamp 0
transform 1 0 2710 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__10820_
timestamp 0
transform -1 0 2010 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__10821_
timestamp 0
transform -1 0 2130 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__10822_
timestamp 0
transform -1 0 1830 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__10823_
timestamp 0
transform 1 0 2110 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__10824_
timestamp 0
transform -1 0 2770 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__10825_
timestamp 0
transform -1 0 2950 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__10826_
timestamp 0
transform -1 0 5030 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__10827_
timestamp 0
transform -1 0 4970 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10828_
timestamp 0
transform -1 0 630 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__10829_
timestamp 0
transform -1 0 430 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__10830_
timestamp 0
transform -1 0 1250 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__10831_
timestamp 0
transform 1 0 1470 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__10832_
timestamp 0
transform 1 0 1330 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__10833_
timestamp 0
transform -1 0 30 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__10834_
timestamp 0
transform 1 0 2230 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10835_
timestamp 0
transform 1 0 2090 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10836_
timestamp 0
transform 1 0 1850 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__10837_
timestamp 0
transform 1 0 2930 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__10838_
timestamp 0
transform 1 0 3350 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__10839_
timestamp 0
transform 1 0 3030 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__10840_
timestamp 0
transform -1 0 1870 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__10841_
timestamp 0
transform 1 0 2990 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10842_
timestamp 0
transform 1 0 2610 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__10843_
timestamp 0
transform -1 0 2770 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__10844_
timestamp 0
transform -1 0 3210 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__10845_
timestamp 0
transform -1 0 4710 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__10846_
timestamp 0
transform 1 0 4810 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__10847_
timestamp 0
transform -1 0 4550 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__10848_
timestamp 0
transform -1 0 3150 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10849_
timestamp 0
transform -1 0 1430 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__10850_
timestamp 0
transform -1 0 1310 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__10851_
timestamp 0
transform -1 0 4410 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__10852_
timestamp 0
transform -1 0 4890 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__10853_
timestamp 0
transform 1 0 1790 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__10854_
timestamp 0
transform -1 0 4470 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__10855_
timestamp 0
transform 1 0 3850 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10856_
timestamp 0
transform 1 0 2630 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10857_
timestamp 0
transform 1 0 3070 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10858_
timestamp 0
transform 1 0 3370 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10859_
timestamp 0
transform -1 0 2950 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__10860_
timestamp 0
transform 1 0 3550 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__10861_
timestamp 0
transform 1 0 3470 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__10862_
timestamp 0
transform 1 0 2850 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__10863_
timestamp 0
transform 1 0 3270 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10864_
timestamp 0
transform 1 0 3410 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10865_
timestamp 0
transform 1 0 3550 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10866_
timestamp 0
transform 1 0 4390 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10867_
timestamp 0
transform 1 0 710 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__10868_
timestamp 0
transform 1 0 1710 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10869_
timestamp 0
transform 1 0 1970 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10870_
timestamp 0
transform 1 0 1810 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10871_
timestamp 0
transform -1 0 2390 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10872_
timestamp 0
transform -1 0 2030 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10873_
timestamp 0
transform -1 0 2170 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10874_
timestamp 0
transform -1 0 2250 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10875_
timestamp 0
transform -1 0 2630 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__10876_
timestamp 0
transform 1 0 2410 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__10877_
timestamp 0
transform 1 0 2170 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__10878_
timestamp 0
transform -1 0 3010 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10879_
timestamp 0
transform -1 0 1910 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__10880_
timestamp 0
transform -1 0 2050 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__10881_
timestamp 0
transform -1 0 2090 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__10882_
timestamp 0
transform -1 0 2270 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__10883_
timestamp 0
transform 1 0 3850 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10884_
timestamp 0
transform -1 0 2310 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10885_
timestamp 0
transform -1 0 2490 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10886_
timestamp 0
transform 1 0 2410 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10887_
timestamp 0
transform -1 0 3110 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10888_
timestamp 0
transform 1 0 3590 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10889_
timestamp 0
transform 1 0 3250 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10890_
timestamp 0
transform 1 0 3430 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10891_
timestamp 0
transform -1 0 4470 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10892_
timestamp 0
transform 1 0 4270 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10893_
timestamp 0
transform -1 0 4430 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10894_
timestamp 0
transform 1 0 4130 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10895_
timestamp 0
transform 1 0 4530 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10896_
timestamp 0
transform 1 0 4490 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10897_
timestamp 0
transform 1 0 4810 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10898_
timestamp 0
transform -1 0 4670 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10899_
timestamp 0
transform -1 0 4590 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__10900_
timestamp 0
transform -1 0 8330 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__10901_
timestamp 0
transform -1 0 7830 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__10902_
timestamp 0
transform -1 0 7950 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__10903_
timestamp 0
transform 1 0 5470 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__10904_
timestamp 0
transform 1 0 4670 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10905_
timestamp 0
transform -1 0 2450 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__10906_
timestamp 0
transform -1 0 2610 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10907_
timestamp 0
transform -1 0 3770 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10908_
timestamp 0
transform -1 0 3570 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10909_
timestamp 0
transform 1 0 3690 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10910_
timestamp 0
transform 1 0 3910 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10911_
timestamp 0
transform 1 0 4610 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10912_
timestamp 0
transform 1 0 4750 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10913_
timestamp 0
transform -1 0 4230 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10914_
timestamp 0
transform 1 0 3990 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10915_
timestamp 0
transform -1 0 4090 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10916_
timestamp 0
transform 1 0 4890 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10917_
timestamp 0
transform 1 0 5030 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10918_
timestamp 0
transform 1 0 5510 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10919_
timestamp 0
transform -1 0 5070 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10920_
timestamp 0
transform 1 0 4810 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10921_
timestamp 0
transform 1 0 4950 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10922_
timestamp 0
transform -1 0 5210 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10923_
timestamp 0
transform 1 0 5190 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__10924_
timestamp 0
transform -1 0 1010 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__10925_
timestamp 0
transform 1 0 5310 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10926_
timestamp 0
transform 1 0 5450 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10927_
timestamp 0
transform 1 0 5610 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10928_
timestamp 0
transform 1 0 5590 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__10929_
timestamp 0
transform 1 0 5350 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10930_
timestamp 0
transform 1 0 5330 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__10931_
timestamp 0
transform 1 0 3630 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__10932_
timestamp 0
transform -1 0 4330 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10933_
timestamp 0
transform 1 0 1230 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__10934_
timestamp 0
transform 1 0 1590 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__10935_
timestamp 0
transform 1 0 1450 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__10936_
timestamp 0
transform 1 0 1730 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__10937_
timestamp 0
transform 1 0 1450 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__10938_
timestamp 0
transform 1 0 1190 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__10939_
timestamp 0
transform -1 0 3810 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__10940_
timestamp 0
transform -1 0 2030 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__10941_
timestamp 0
transform 1 0 1810 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__10942_
timestamp 0
transform 1 0 3350 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__10943_
timestamp 0
transform 1 0 3630 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__10944_
timestamp 0
transform 1 0 3490 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__10945_
timestamp 0
transform -1 0 3770 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__10946_
timestamp 0
transform 1 0 4030 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__10947_
timestamp 0
transform 1 0 3890 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__10948_
timestamp 0
transform -1 0 4510 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__10949_
timestamp 0
transform -1 0 4630 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__10950_
timestamp 0
transform -1 0 5050 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__10951_
timestamp 0
transform -1 0 5190 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__10952_
timestamp 0
transform -1 0 5370 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__10953_
timestamp 0
transform -1 0 4750 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__10954_
timestamp 0
transform -1 0 4510 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__10955_
timestamp 0
transform -1 0 1750 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__10956_
timestamp 0
transform -1 0 1430 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__10957_
timestamp 0
transform -1 0 1550 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__10958_
timestamp 0
transform 1 0 1670 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__10959_
timestamp 0
transform 1 0 1590 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__10960_
timestamp 0
transform 1 0 3270 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__10961_
timestamp 0
transform 1 0 2370 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__10962_
timestamp 0
transform 1 0 2730 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__10963_
timestamp 0
transform 1 0 3630 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__10964_
timestamp 0
transform 1 0 3930 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__10965_
timestamp 0
transform -1 0 3370 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__10966_
timestamp 0
transform 1 0 3490 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__10967_
timestamp 0
transform 1 0 4390 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__10968_
timestamp 0
transform 1 0 3730 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__10969_
timestamp 0
transform -1 0 3610 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__10970_
timestamp 0
transform 1 0 3850 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__10971_
timestamp 0
transform -1 0 4730 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__10972_
timestamp 0
transform 1 0 4870 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__10973_
timestamp 0
transform 1 0 5030 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__10974_
timestamp 0
transform -1 0 5750 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__10975_
timestamp 0
transform -1 0 4990 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__10976_
timestamp 0
transform -1 0 4110 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__10977_
timestamp 0
transform 1 0 3770 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__10978_
timestamp 0
transform 1 0 1110 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__10979_
timestamp 0
transform 1 0 1250 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__10980_
timestamp 0
transform -1 0 1330 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__10981_
timestamp 0
transform 1 0 2510 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__10982_
timestamp 0
transform 1 0 2430 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__10983_
timestamp 0
transform 1 0 3790 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__10984_
timestamp 0
transform 1 0 2850 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__10985_
timestamp 0
transform -1 0 3110 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__10986_
timestamp 0
transform 1 0 3190 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__10987_
timestamp 0
transform 1 0 4070 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__10988_
timestamp 0
transform 1 0 4210 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__10989_
timestamp 0
transform 1 0 4830 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__10990_
timestamp 0
transform 1 0 5050 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__10991_
timestamp 0
transform 1 0 5110 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__10992_
timestamp 0
transform 1 0 5270 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__10993_
timestamp 0
transform 1 0 5410 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__10994_
timestamp 0
transform 1 0 5410 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__10995_
timestamp 0
transform -1 0 5930 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__10996_
timestamp 0
transform 1 0 1930 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__10997_
timestamp 0
transform -1 0 3170 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__10998_
timestamp 0
transform -1 0 1250 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__10999_
timestamp 0
transform -1 0 2930 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11000_
timestamp 0
transform -1 0 2210 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11001_
timestamp 0
transform 1 0 2470 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11002_
timestamp 0
transform 1 0 2630 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11003_
timestamp 0
transform -1 0 3650 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11004_
timestamp 0
transform 1 0 3170 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11005_
timestamp 0
transform 1 0 2870 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11006_
timestamp 0
transform 1 0 2730 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11007_
timestamp 0
transform 1 0 3290 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11008_
timestamp 0
transform 1 0 3410 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11009_
timestamp 0
transform 1 0 3870 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11010_
timestamp 0
transform 1 0 4230 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11011_
timestamp 0
transform -1 0 4370 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11012_
timestamp 0
transform -1 0 4570 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11013_
timestamp 0
transform -1 0 4630 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11014_
timestamp 0
transform 1 0 5170 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11015_
timestamp 0
transform 1 0 5310 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11016_
timestamp 0
transform -1 0 5770 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11017_
timestamp 0
transform 1 0 5710 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11018_
timestamp 0
transform 1 0 3030 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11019_
timestamp 0
transform 1 0 4830 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11020_
timestamp 0
transform -1 0 4910 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11021_
timestamp 0
transform 1 0 4470 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11022_
timestamp 0
transform -1 0 4750 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11023_
timestamp 0
transform -1 0 3750 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11024_
timestamp 0
transform -1 0 1270 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11025_
timestamp 0
transform -1 0 3030 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11026_
timestamp 0
transform -1 0 2090 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11027_
timestamp 0
transform -1 0 2130 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11028_
timestamp 0
transform -1 0 2030 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11029_
timestamp 0
transform -1 0 1410 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11030_
timestamp 0
transform -1 0 1550 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11031_
timestamp 0
transform 1 0 1670 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11032_
timestamp 0
transform -1 0 2330 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11033_
timestamp 0
transform 1 0 1770 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11034_
timestamp 0
transform 1 0 1370 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11035_
timestamp 0
transform 1 0 1890 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11036_
timestamp 0
transform 1 0 2170 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11037_
timestamp 0
transform 1 0 2030 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11038_
timestamp 0
transform 1 0 3990 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11039_
timestamp 0
transform 1 0 4230 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11040_
timestamp 0
transform -1 0 4130 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11041_
timestamp 0
transform -1 0 4550 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11042_
timestamp 0
transform 1 0 4690 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11043_
timestamp 0
transform 1 0 5210 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11044_
timestamp 0
transform 1 0 5370 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11045_
timestamp 0
transform 1 0 5170 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11046_
timestamp 0
transform -1 0 5330 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11047_
timestamp 0
transform -1 0 5650 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11048_
timestamp 0
transform -1 0 4130 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11049_
timestamp 0
transform 1 0 4410 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11050_
timestamp 0
transform -1 0 4290 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11051_
timestamp 0
transform -1 0 2770 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11052_
timestamp 0
transform 1 0 2170 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11053_
timestamp 0
transform -1 0 1570 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11054_
timestamp 0
transform 1 0 2310 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11055_
timestamp 0
transform -1 0 1950 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11056_
timestamp 0
transform 1 0 2330 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11057_
timestamp 0
transform 1 0 2590 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11058_
timestamp 0
transform -1 0 2610 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11059_
timestamp 0
transform 1 0 2450 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11060_
timestamp 0
transform -1 0 2450 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11061_
timestamp 0
transform 1 0 2870 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11062_
timestamp 0
transform -1 0 3870 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11063_
timestamp 0
transform 1 0 4890 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11064_
timestamp 0
transform 1 0 5010 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11065_
timestamp 0
transform 1 0 5150 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11066_
timestamp 0
transform -1 0 5490 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11067_
timestamp 0
transform -1 0 3310 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11068_
timestamp 0
transform 1 0 3570 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11069_
timestamp 0
transform -1 0 3450 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11070_
timestamp 0
transform 1 0 3570 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11071_
timestamp 0
transform -1 0 3730 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11072_
timestamp 0
transform -1 0 4010 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11073_
timestamp 0
transform 1 0 3930 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11074_
timestamp 0
transform 1 0 3230 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11075_
timestamp 0
transform 1 0 1710 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11076_
timestamp 0
transform 1 0 2930 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11077_
timestamp 0
transform -1 0 2290 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11078_
timestamp 0
transform 1 0 3090 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11079_
timestamp 0
transform 1 0 2590 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11080_
timestamp 0
transform 1 0 2810 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11081_
timestamp 0
transform 1 0 3490 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11082_
timestamp 0
transform 1 0 3030 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11083_
timestamp 0
transform 1 0 2950 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11084_
timestamp 0
transform 1 0 3190 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11085_
timestamp 0
transform 1 0 4010 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11086_
timestamp 0
transform 1 0 4430 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11087_
timestamp 0
transform 1 0 4590 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11088_
timestamp 0
transform 1 0 4730 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11089_
timestamp 0
transform -1 0 5450 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11090_
timestamp 0
transform -1 0 3770 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11091_
timestamp 0
transform 1 0 2110 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11092_
timestamp 0
transform 1 0 2710 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11093_
timestamp 0
transform 1 0 2630 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11094_
timestamp 0
transform 1 0 2770 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11095_
timestamp 0
transform -1 0 2970 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11096_
timestamp 0
transform -1 0 3510 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11097_
timestamp 0
transform 1 0 3630 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11098_
timestamp 0
transform -1 0 3930 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11099_
timestamp 0
transform 1 0 3530 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11100_
timestamp 0
transform 1 0 3070 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11101_
timestamp 0
transform -1 0 3410 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11102_
timestamp 0
transform 1 0 3770 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11103_
timestamp 0
transform -1 0 4350 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11104_
timestamp 0
transform 1 0 3350 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11105_
timestamp 0
transform 1 0 4070 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11106_
timestamp 0
transform 1 0 4290 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11107_
timestamp 0
transform 1 0 4350 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11108_
timestamp 0
transform 1 0 4470 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11109_
timestamp 0
transform 1 0 4150 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11110_
timestamp 0
transform 1 0 4190 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11111_
timestamp 0
transform 1 0 4890 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11112_
timestamp 0
transform 1 0 5070 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11113_
timestamp 0
transform -1 0 5710 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__11114_
timestamp 0
transform -1 0 6070 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11115_
timestamp 0
transform 1 0 4630 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11116_
timestamp 0
transform -1 0 2590 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11117_
timestamp 0
transform -1 0 2430 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11118_
timestamp 0
transform -1 0 1970 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11119_
timestamp 0
transform -1 0 2470 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11120_
timestamp 0
transform -1 0 3010 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11121_
timestamp 0
transform 1 0 3110 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11122_
timestamp 0
transform 1 0 3250 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11123_
timestamp 0
transform 1 0 3230 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11124_
timestamp 0
transform 1 0 4430 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11125_
timestamp 0
transform 1 0 4530 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11126_
timestamp 0
transform -1 0 4770 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11127_
timestamp 0
transform 1 0 4770 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11128_
timestamp 0
transform 1 0 4930 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11129_
timestamp 0
transform -1 0 5930 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11130_
timestamp 0
transform 1 0 1970 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11131_
timestamp 0
transform -1 0 3430 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11132_
timestamp 0
transform 1 0 3490 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11133_
timestamp 0
transform -1 0 3370 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11134_
timestamp 0
transform 1 0 2310 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11135_
timestamp 0
transform -1 0 4070 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11136_
timestamp 0
transform 1 0 3690 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11137_
timestamp 0
transform -1 0 4250 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__11138_
timestamp 0
transform -1 0 2190 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11139_
timestamp 0
transform 1 0 1110 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11140_
timestamp 0
transform 1 0 970 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11141_
timestamp 0
transform -1 0 4070 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11142_
timestamp 0
transform -1 0 4210 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11143_
timestamp 0
transform 1 0 710 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11144_
timestamp 0
transform 1 0 130 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11145_
timestamp 0
transform -1 0 1450 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11146_
timestamp 0
transform -1 0 1350 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11147_
timestamp 0
transform 1 0 870 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11148_
timestamp 0
transform -1 0 1130 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11149_
timestamp 0
transform 1 0 990 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11150_
timestamp 0
transform 1 0 1730 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11151_
timestamp 0
transform -1 0 1630 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11152_
timestamp 0
transform 1 0 1590 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11153_
timestamp 0
transform -1 0 2530 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11154_
timestamp 0
transform -1 0 1910 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__11155_
timestamp 0
transform 1 0 3350 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11156_
timestamp 0
transform 1 0 3210 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11157_
timestamp 0
transform 1 0 3510 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11158_
timestamp 0
transform -1 0 3650 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11159_
timestamp 0
transform 1 0 1670 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11160_
timestamp 0
transform 1 0 430 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11161_
timestamp 0
transform 1 0 850 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11162_
timestamp 0
transform -1 0 730 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11163_
timestamp 0
transform -1 0 30 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11164_
timestamp 0
transform 1 0 1810 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11165_
timestamp 0
transform 1 0 1650 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11166_
timestamp 0
transform 1 0 290 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11167_
timestamp 0
transform 1 0 130 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__11168_
timestamp 0
transform 1 0 290 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11169_
timestamp 0
transform 1 0 1210 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11170_
timestamp 0
transform 1 0 530 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11171_
timestamp 0
transform -1 0 730 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11172_
timestamp 0
transform -1 0 1590 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11173_
timestamp 0
transform 1 0 1630 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11174_
timestamp 0
transform 1 0 1830 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11175_
timestamp 0
transform -1 0 1490 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11176_
timestamp 0
transform 1 0 1930 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11177_
timestamp 0
transform 1 0 1930 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11178_
timestamp 0
transform -1 0 1810 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11179_
timestamp 0
transform 1 0 2070 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11180_
timestamp 0
transform 1 0 2370 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11181_
timestamp 0
transform -1 0 2130 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11182_
timestamp 0
transform -1 0 1690 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11183_
timestamp 0
transform 1 0 1150 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11184_
timestamp 0
transform 1 0 1510 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11185_
timestamp 0
transform 1 0 1370 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11186_
timestamp 0
transform 1 0 570 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11187_
timestamp 0
transform -1 0 450 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11188_
timestamp 0
transform 1 0 1830 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11189_
timestamp 0
transform 1 0 1270 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11190_
timestamp 0
transform -1 0 1170 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11191_
timestamp 0
transform 1 0 870 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11192_
timestamp 0
transform 1 0 770 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11193_
timestamp 0
transform 1 0 870 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11194_
timestamp 0
transform -1 0 1290 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11195_
timestamp 0
transform -1 0 1030 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11196_
timestamp 0
transform -1 0 910 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11197_
timestamp 0
transform 1 0 1030 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11198_
timestamp 0
transform 1 0 1050 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11199_
timestamp 0
transform 1 0 1130 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11200_
timestamp 0
transform 1 0 1390 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11201_
timestamp 0
transform -1 0 1270 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11202_
timestamp 0
transform 1 0 1530 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11203_
timestamp 0
transform 1 0 1950 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11204_
timestamp 0
transform -1 0 910 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11205_
timestamp 0
transform -1 0 310 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11206_
timestamp 0
transform 1 0 1970 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11207_
timestamp 0
transform 1 0 1870 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11208_
timestamp 0
transform -1 0 590 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11209_
timestamp 0
transform 1 0 150 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11210_
timestamp 0
transform -1 0 1550 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11211_
timestamp 0
transform -1 0 1310 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11212_
timestamp 0
transform 1 0 1410 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11213_
timestamp 0
transform -1 0 30 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11214_
timestamp 0
transform -1 0 750 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11215_
timestamp 0
transform 1 0 290 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11216_
timestamp 0
transform 1 0 310 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11217_
timestamp 0
transform 1 0 550 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11218_
timestamp 0
transform -1 0 170 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11219_
timestamp 0
transform -1 0 430 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11220_
timestamp 0
transform -1 0 30 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11221_
timestamp 0
transform 1 0 150 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11222_
timestamp 0
transform -1 0 30 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11223_
timestamp 0
transform 1 0 390 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11224_
timestamp 0
transform -1 0 2330 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11225_
timestamp 0
transform -1 0 270 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11226_
timestamp 0
transform -1 0 2550 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11227_
timestamp 0
transform -1 0 2670 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11228_
timestamp 0
transform -1 0 290 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11229_
timestamp 0
transform -1 0 290 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11230_
timestamp 0
transform 1 0 10 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11231_
timestamp 0
transform -1 0 150 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__11232_
timestamp 0
transform 1 0 310 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11233_
timestamp 0
transform -1 0 470 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11234_
timestamp 0
transform 1 0 130 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11235_
timestamp 0
transform -1 0 170 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__11236_
timestamp 0
transform -1 0 30 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11237_
timestamp 0
transform -1 0 30 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11238_
timestamp 0
transform -1 0 30 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__11239_
timestamp 0
transform 1 0 290 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__11240_
timestamp 0
transform 1 0 170 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11241_
timestamp 0
transform -1 0 30 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11242_
timestamp 0
transform -1 0 30 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11243_
timestamp 0
transform 1 0 310 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11244_
timestamp 0
transform -1 0 190 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11245_
timestamp 0
transform -1 0 470 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11246_
timestamp 0
transform -1 0 1130 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11247_
timestamp 0
transform -1 0 190 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11248_
timestamp 0
transform -1 0 30 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11249_
timestamp 0
transform -1 0 30 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__11250_
timestamp 0
transform 1 0 1070 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11251_
timestamp 0
transform -1 0 770 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11252_
timestamp 0
transform -1 0 30 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11253_
timestamp 0
transform -1 0 150 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11254_
timestamp 0
transform 1 0 450 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__11255_
timestamp 0
transform -1 0 290 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__11256_
timestamp 0
transform -1 0 190 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11257_
timestamp 0
transform 1 0 590 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11258_
timestamp 0
transform -1 0 530 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11259_
timestamp 0
transform 1 0 430 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11260_
timestamp 0
transform -1 0 330 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11261_
timestamp 0
transform -1 0 190 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11262_
timestamp 0
transform 1 0 470 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11263_
timestamp 0
transform -1 0 150 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11264_
timestamp 0
transform -1 0 30 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11265_
timestamp 0
transform 1 0 130 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11266_
timestamp 0
transform 1 0 290 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11267_
timestamp 0
transform -1 0 30 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11268_
timestamp 0
transform -1 0 1490 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11269_
timestamp 0
transform 1 0 130 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__11270_
timestamp 0
transform -1 0 930 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__11271_
timestamp 0
transform 1 0 530 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11272_
timestamp 0
transform 1 0 450 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__11273_
timestamp 0
transform 1 0 410 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__11274_
timestamp 0
transform 1 0 670 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11275_
timestamp 0
transform -1 0 570 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11276_
timestamp 0
transform -1 0 690 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11277_
timestamp 0
transform -1 0 430 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11278_
timestamp 0
transform -1 0 570 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11279_
timestamp 0
transform 1 0 550 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11280_
timestamp 0
transform -1 0 690 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11281_
timestamp 0
transform 1 0 170 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11282_
timestamp 0
transform -1 0 130 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11283_
timestamp 0
transform -1 0 290 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11284_
timestamp 0
transform 1 0 410 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11285_
timestamp 0
transform -1 0 570 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11286_
timestamp 0
transform 1 0 690 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11287_
timestamp 0
transform 1 0 10 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11288_
timestamp 0
transform 1 0 270 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11289_
timestamp 0
transform 1 0 250 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11290_
timestamp 0
transform 1 0 410 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11291_
timestamp 0
transform 1 0 830 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11292_
timestamp 0
transform 1 0 970 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11293_
timestamp 0
transform -1 0 1210 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11294_
timestamp 0
transform -1 0 1330 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11295_
timestamp 0
transform -1 0 1210 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11296_
timestamp 0
transform -1 0 590 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11297_
timestamp 0
transform 1 0 810 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11298_
timestamp 0
transform -1 0 1170 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11299_
timestamp 0
transform -1 0 970 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11300_
timestamp 0
transform 1 0 270 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11301_
timestamp 0
transform 1 0 870 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11302_
timestamp 0
transform 1 0 710 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__11303_
timestamp 0
transform 1 0 550 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__11304_
timestamp 0
transform -1 0 690 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__11305_
timestamp 0
transform -1 0 750 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11306_
timestamp 0
transform 1 0 790 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__11307_
timestamp 0
transform -1 0 570 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__11308_
timestamp 0
transform -1 0 970 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__11309_
timestamp 0
transform 1 0 710 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11310_
timestamp 0
transform 1 0 130 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11311_
timestamp 0
transform -1 0 30 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11312_
timestamp 0
transform 1 0 430 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11313_
timestamp 0
transform 1 0 530 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11314_
timestamp 0
transform -1 0 810 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11315_
timestamp 0
transform 1 0 670 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11316_
timestamp 0
transform 1 0 790 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11317_
timestamp 0
transform 1 0 910 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11318_
timestamp 0
transform -1 0 850 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11319_
timestamp 0
transform 1 0 810 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__11320_
timestamp 0
transform -1 0 30 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__11321_
timestamp 0
transform -1 0 30 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11322_
timestamp 0
transform -1 0 1090 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11323_
timestamp 0
transform 1 0 1210 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__11324_
timestamp 0
transform 1 0 930 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11325_
timestamp 0
transform -1 0 970 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__11326_
timestamp 0
transform 1 0 1030 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11327_
timestamp 0
transform -1 0 1290 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__11328_
timestamp 0
transform -1 0 1110 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__11329_
timestamp 0
transform 1 0 1110 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__11330_
timestamp 0
transform -1 0 710 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11331_
timestamp 0
transform -1 0 710 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11332_
timestamp 0
transform 1 0 1250 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11333_
timestamp 0
transform -1 0 310 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11334_
timestamp 0
transform -1 0 530 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11335_
timestamp 0
transform 1 0 850 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11336_
timestamp 0
transform -1 0 450 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11337_
timestamp 0
transform -1 0 570 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11338_
timestamp 0
transform 1 0 650 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11339_
timestamp 0
transform 1 0 1350 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__11340_
timestamp 0
transform 1 0 1430 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__11341_
timestamp 0
transform 1 0 1310 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11342_
timestamp 0
transform -1 0 1190 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11343_
timestamp 0
transform -1 0 1110 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11344_
timestamp 0
transform -1 0 970 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11345_
timestamp 0
transform -1 0 990 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11346_
timestamp 0
transform 1 0 1110 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11347_
timestamp 0
transform -1 0 850 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11348_
timestamp 0
transform 1 0 970 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11349_
timestamp 0
transform -1 0 710 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11350_
timestamp 0
transform -1 0 1830 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11351_
timestamp 0
transform -1 0 1070 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11352_
timestamp 0
transform 1 0 1170 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11353_
timestamp 0
transform -1 0 850 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11354_
timestamp 0
transform 1 0 1090 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11355_
timestamp 0
transform 1 0 1310 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11356_
timestamp 0
transform 1 0 790 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11357_
timestamp 0
transform 1 0 1050 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__11358_
timestamp 0
transform 1 0 1190 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11359_
timestamp 0
transform 1 0 1350 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11360_
timestamp 0
transform -1 0 1510 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11361_
timestamp 0
transform 1 0 1470 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__11362_
timestamp 0
transform -1 0 1590 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__11363_
timestamp 0
transform 1 0 1630 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__11364_
timestamp 0
transform -1 0 1630 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__11365_
timestamp 0
transform 1 0 1730 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__11366_
timestamp 0
transform -1 0 1490 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11367_
timestamp 0
transform 1 0 1590 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11368_
timestamp 0
transform -1 0 1470 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11369_
timestamp 0
transform 1 0 1730 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11370_
timestamp 0
transform -1 0 1650 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11371_
timestamp 0
transform -1 0 1570 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11372_
timestamp 0
transform -1 0 1430 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11373_
timestamp 0
transform 1 0 1530 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11374_
timestamp 0
transform 1 0 1350 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11375_
timestamp 0
transform -1 0 2350 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11376_
timestamp 0
transform -1 0 2730 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11377_
timestamp 0
transform -1 0 2490 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__11378_
timestamp 0
transform 1 0 1830 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11379_
timestamp 0
transform -1 0 1690 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11380_
timestamp 0
transform -1 0 1690 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11381_
timestamp 0
transform -1 0 2390 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11382_
timestamp 0
transform 1 0 4210 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11383_
timestamp 0
transform 1 0 4370 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11384_
timestamp 0
transform -1 0 3950 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11385_
timestamp 0
transform 1 0 4470 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11386_
timestamp 0
transform 1 0 4730 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11387_
timestamp 0
transform 1 0 5950 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11388_
timestamp 0
transform 1 0 5390 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11389_
timestamp 0
transform -1 0 6090 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11390_
timestamp 0
transform 1 0 4690 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11391_
timestamp 0
transform -1 0 3570 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11392_
timestamp 0
transform -1 0 3670 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11393_
timestamp 0
transform 1 0 4590 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11394_
timestamp 0
transform 1 0 3770 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11395_
timestamp 0
transform 1 0 4710 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11396_
timestamp 0
transform -1 0 4870 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11397_
timestamp 0
transform 1 0 5150 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11398_
timestamp 0
transform 1 0 5010 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11399_
timestamp 0
transform 1 0 5290 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11400_
timestamp 0
transform 1 0 5430 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11401_
timestamp 0
transform 1 0 4930 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11402_
timestamp 0
transform 1 0 5790 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11403_
timestamp 0
transform 1 0 5910 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11404_
timestamp 0
transform -1 0 4610 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11405_
timestamp 0
transform 1 0 4790 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11406_
timestamp 0
transform -1 0 2770 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11407_
timestamp 0
transform 1 0 3250 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11408_
timestamp 0
transform 1 0 3070 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11409_
timestamp 0
transform -1 0 4090 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11410_
timestamp 0
transform 1 0 4190 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11411_
timestamp 0
transform -1 0 4370 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11412_
timestamp 0
transform 1 0 4370 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11413_
timestamp 0
transform 1 0 5190 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11414_
timestamp 0
transform -1 0 5090 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11415_
timestamp 0
transform -1 0 5350 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11416_
timestamp 0
transform -1 0 5490 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11417_
timestamp 0
transform -1 0 6670 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11418_
timestamp 0
transform 1 0 5290 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11419_
timestamp 0
transform -1 0 6270 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11420_
timestamp 0
transform 1 0 5170 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11421_
timestamp 0
transform -1 0 3590 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11422_
timestamp 0
transform -1 0 3710 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11423_
timestamp 0
transform 1 0 3390 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11424_
timestamp 0
transform 1 0 3590 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11425_
timestamp 0
transform 1 0 6630 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11426_
timestamp 0
transform -1 0 6530 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11427_
timestamp 0
transform 1 0 7150 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11428_
timestamp 0
transform 1 0 7030 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11429_
timestamp 0
transform -1 0 6370 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11430_
timestamp 0
transform 1 0 6490 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11431_
timestamp 0
transform 1 0 6770 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11432_
timestamp 0
transform 1 0 6090 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11433_
timestamp 0
transform 1 0 6490 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__11434_
timestamp 0
transform 1 0 3790 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11435_
timestamp 0
transform 1 0 3950 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11436_
timestamp 0
transform -1 0 4470 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11437_
timestamp 0
transform 1 0 6670 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11438_
timestamp 0
transform -1 0 6470 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11439_
timestamp 0
transform 1 0 6830 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11440_
timestamp 0
transform 1 0 6890 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11441_
timestamp 0
transform -1 0 6110 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11442_
timestamp 0
transform -1 0 5970 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11443_
timestamp 0
transform -1 0 5830 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11444_
timestamp 0
transform 1 0 6970 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11445_
timestamp 0
transform 1 0 6110 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__11446_
timestamp 0
transform -1 0 3910 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11447_
timestamp 0
transform -1 0 3910 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11448_
timestamp 0
transform 1 0 3990 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11449_
timestamp 0
transform 1 0 4130 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11450_
timestamp 0
transform 1 0 6350 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__11451_
timestamp 0
transform -1 0 6230 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__11452_
timestamp 0
transform 1 0 6590 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__11453_
timestamp 0
transform 1 0 6870 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__11454_
timestamp 0
transform 1 0 7290 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11455_
timestamp 0
transform 1 0 7250 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__11456_
timestamp 0
transform -1 0 7390 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__11457_
timestamp 0
transform 1 0 7130 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11458_
timestamp 0
transform -1 0 6390 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11459_
timestamp 0
transform -1 0 6350 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11460_
timestamp 0
transform -1 0 6450 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11461_
timestamp 0
transform -1 0 6730 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__11462_
timestamp 0
transform -1 0 6590 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11463_
timestamp 0
transform 1 0 6550 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11464_
timestamp 0
transform 1 0 3850 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11465_
timestamp 0
transform -1 0 4290 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11466_
timestamp 0
transform -1 0 4570 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11467_
timestamp 0
transform 1 0 4410 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11468_
timestamp 0
transform 1 0 4670 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11469_
timestamp 0
transform -1 0 5190 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11470_
timestamp 0
transform 1 0 5290 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11471_
timestamp 0
transform -1 0 5470 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11472_
timestamp 0
transform 1 0 6050 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11473_
timestamp 0
transform 1 0 7030 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11474_
timestamp 0
transform 1 0 6910 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11475_
timestamp 0
transform 1 0 6750 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11476_
timestamp 0
transform -1 0 6790 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11477_
timestamp 0
transform 1 0 5670 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11478_
timestamp 0
transform 1 0 6050 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11479_
timestamp 0
transform 1 0 5290 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11480_
timestamp 0
transform -1 0 3390 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11481_
timestamp 0
transform 1 0 3510 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11482_
timestamp 0
transform 1 0 3650 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11483_
timestamp 0
transform 1 0 5630 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11484_
timestamp 0
transform 1 0 5750 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11485_
timestamp 0
transform -1 0 5530 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11486_
timestamp 0
transform 1 0 5870 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11487_
timestamp 0
transform 1 0 6110 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11488_
timestamp 0
transform -1 0 5990 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11489_
timestamp 0
transform 1 0 5790 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11490_
timestamp 0
transform -1 0 5450 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11491_
timestamp 0
transform -1 0 2530 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11492_
timestamp 0
transform 1 0 2630 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11493_
timestamp 0
transform 1 0 3050 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11494_
timestamp 0
transform -1 0 3490 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11495_
timestamp 0
transform 1 0 3190 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11496_
timestamp 0
transform 1 0 3330 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11497_
timestamp 0
transform -1 0 6010 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11498_
timestamp 0
transform -1 0 5950 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11499_
timestamp 0
transform -1 0 6050 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11500_
timestamp 0
transform -1 0 6210 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11501_
timestamp 0
transform -1 0 5890 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11502_
timestamp 0
transform 1 0 5050 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11503_
timestamp 0
transform -1 0 4930 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11504_
timestamp 0
transform -1 0 5190 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11505_
timestamp 0
transform 1 0 5290 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11506_
timestamp 0
transform -1 0 4310 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11507_
timestamp 0
transform -1 0 3750 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11508_
timestamp 0
transform -1 0 3810 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11509_
timestamp 0
transform -1 0 3890 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11510_
timestamp 0
transform 1 0 4450 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11511_
timestamp 0
transform 1 0 4590 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11512_
timestamp 0
transform -1 0 4770 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11513_
timestamp 0
transform 1 0 5150 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11514_
timestamp 0
transform 1 0 3990 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11515_
timestamp 0
transform 1 0 4130 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11516_
timestamp 0
transform 1 0 4470 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11517_
timestamp 0
transform 1 0 4570 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11518_
timestamp 0
transform 1 0 3270 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11519_
timestamp 0
transform -1 0 3410 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11520_
timestamp 0
transform -1 0 3530 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11521_
timestamp 0
transform 1 0 3650 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11522_
timestamp 0
transform -1 0 4490 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11523_
timestamp 0
transform 1 0 4630 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11524_
timestamp 0
transform 1 0 4770 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11525_
timestamp 0
transform 1 0 5250 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11526_
timestamp 0
transform -1 0 4610 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11527_
timestamp 0
transform 1 0 5090 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11528_
timestamp 0
transform -1 0 4050 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11529_
timestamp 0
transform 1 0 2670 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11530_
timestamp 0
transform -1 0 3770 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11531_
timestamp 0
transform 1 0 2090 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11532_
timestamp 0
transform 1 0 2030 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11533_
timestamp 0
transform 1 0 2790 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11534_
timestamp 0
transform 1 0 2690 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11535_
timestamp 0
transform -1 0 2070 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11536_
timestamp 0
transform -1 0 3430 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11537_
timestamp 0
transform -1 0 2470 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11538_
timestamp 0
transform -1 0 2630 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11539_
timestamp 0
transform -1 0 2750 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11540_
timestamp 0
transform -1 0 2470 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11541_
timestamp 0
transform -1 0 2610 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11542_
timestamp 0
transform -1 0 3290 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11543_
timestamp 0
transform -1 0 2170 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11544_
timestamp 0
transform -1 0 2290 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11545_
timestamp 0
transform -1 0 2310 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11546_
timestamp 0
transform -1 0 2430 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11547_
timestamp 0
transform 1 0 1970 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11548_
timestamp 0
transform 1 0 2170 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11549_
timestamp 0
transform 1 0 2010 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11550_
timestamp 0
transform 1 0 2870 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__11551_
timestamp 0
transform 1 0 2710 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__11552_
timestamp 0
transform -1 0 3410 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11553_
timestamp 0
transform 1 0 3230 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11554_
timestamp 0
transform -1 0 3210 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11555_
timestamp 0
transform 1 0 3050 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11556_
timestamp 0
transform 1 0 2610 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11557_
timestamp 0
transform -1 0 2490 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11558_
timestamp 0
transform 1 0 2930 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__11559_
timestamp 0
transform 1 0 2790 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__11560_
timestamp 0
transform -1 0 4110 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11561_
timestamp 0
transform 1 0 3930 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11562_
timestamp 0
transform -1 0 3170 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11563_
timestamp 0
transform 1 0 3090 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__11564_
timestamp 0
transform -1 0 4250 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11565_
timestamp 0
transform 1 0 3690 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11566_
timestamp 0
transform -1 0 4110 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11567_
timestamp 0
transform 1 0 3530 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__11568_
timestamp 0
transform -1 0 3270 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11569_
timestamp 0
transform -1 0 3430 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__11570_
timestamp 0
transform 1 0 4170 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11571_
timestamp 0
transform 1 0 4310 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11572_
timestamp 0
transform 1 0 3290 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11573_
timestamp 0
transform -1 0 3430 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__11574_
timestamp 0
transform 1 0 4990 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11575_
timestamp 0
transform 1 0 4830 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11576_
timestamp 0
transform 1 0 4370 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11577_
timestamp 0
transform 1 0 4210 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__11578_
timestamp 0
transform -1 0 4270 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11579_
timestamp 0
transform -1 0 4130 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11580_
timestamp 0
transform 1 0 3330 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11581_
timestamp 0
transform -1 0 3510 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__11582_
timestamp 0
transform 1 0 5090 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11583_
timestamp 0
transform 1 0 4950 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11584_
timestamp 0
transform -1 0 3630 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11585_
timestamp 0
transform 1 0 3750 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__11586_
timestamp 0
transform -1 0 3590 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11587_
timestamp 0
transform 1 0 3290 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11588_
timestamp 0
transform -1 0 3270 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11589_
timestamp 0
transform -1 0 3110 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11590_
timestamp 0
transform 1 0 6230 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11591_
timestamp 0
transform 1 0 2910 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__11592_
timestamp 0
transform -1 0 3790 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11593_
timestamp 0
transform 1 0 4170 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11594_
timestamp 0
transform 1 0 3830 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11595_
timestamp 0
transform -1 0 4010 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11596_
timestamp 0
transform -1 0 4810 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11597_
timestamp 0
transform 1 0 4650 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11598_
timestamp 0
transform 1 0 4530 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11599_
timestamp 0
transform 1 0 4370 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__11600_
timestamp 0
transform -1 0 6810 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__11601_
timestamp 0
transform 1 0 6630 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__11602_
timestamp 0
transform -1 0 5870 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__11603_
timestamp 0
transform -1 0 5990 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__11604_
timestamp 0
transform 1 0 3930 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11605_
timestamp 0
transform -1 0 4110 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11606_
timestamp 0
transform 1 0 4770 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11607_
timestamp 0
transform 1 0 4630 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__11608_
timestamp 0
transform -1 0 3710 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11609_
timestamp 0
transform -1 0 3850 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11610_
timestamp 0
transform -1 0 4110 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11611_
timestamp 0
transform -1 0 4230 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11692_
timestamp 0
transform 1 0 9870 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__11693_
timestamp 0
transform 1 0 11310 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11694_
timestamp 0
transform -1 0 12610 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__11695_
timestamp 0
transform 1 0 13250 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__11696_
timestamp 0
transform 1 0 11490 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__11697_
timestamp 0
transform -1 0 11410 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11698_
timestamp 0
transform -1 0 11750 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11699_
timestamp 0
transform -1 0 11070 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__11700_
timestamp 0
transform -1 0 11830 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__11701_
timestamp 0
transform -1 0 11570 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11702_
timestamp 0
transform -1 0 10790 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11703_
timestamp 0
transform -1 0 10910 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__11704_
timestamp 0
transform -1 0 11210 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11705_
timestamp 0
transform -1 0 11870 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__11706_
timestamp 0
transform 1 0 12030 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__11707_
timestamp 0
transform 1 0 11470 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11708_
timestamp 0
transform -1 0 11890 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11709_
timestamp 0
transform -1 0 11610 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11710_
timestamp 0
transform 1 0 9590 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11711_
timestamp 0
transform 1 0 10770 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11712_
timestamp 0
transform -1 0 10910 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11713_
timestamp 0
transform 1 0 11050 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11714_
timestamp 0
transform 1 0 11390 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__11715_
timestamp 0
transform 1 0 11190 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11716_
timestamp 0
transform -1 0 13770 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11717_
timestamp 0
transform -1 0 13470 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11718_
timestamp 0
transform -1 0 13630 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11719_
timestamp 0
transform -1 0 13530 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11720_
timestamp 0
transform -1 0 13110 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11721_
timestamp 0
transform 1 0 12950 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11722_
timestamp 0
transform -1 0 12910 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11723_
timestamp 0
transform -1 0 12410 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11724_
timestamp 0
transform 1 0 12830 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11725_
timestamp 0
transform -1 0 13350 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11726_
timestamp 0
transform 1 0 13150 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11727_
timestamp 0
transform 1 0 13310 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11728_
timestamp 0
transform 1 0 12430 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11729_
timestamp 0
transform 1 0 12810 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11730_
timestamp 0
transform 1 0 12670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11731_
timestamp 0
transform -1 0 12750 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11732_
timestamp 0
transform 1 0 12550 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11733_
timestamp 0
transform 1 0 12710 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11734_
timestamp 0
transform -1 0 13190 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11735_
timestamp 0
transform -1 0 13010 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11736_
timestamp 0
transform -1 0 13030 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11737_
timestamp 0
transform -1 0 13390 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11738_
timestamp 0
transform -1 0 12330 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11739_
timestamp 0
transform -1 0 12470 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11740_
timestamp 0
transform -1 0 12610 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11741_
timestamp 0
transform 1 0 12950 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__11742_
timestamp 0
transform -1 0 12910 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11743_
timestamp 0
transform -1 0 14550 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11744_
timestamp 0
transform 1 0 12870 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11745_
timestamp 0
transform -1 0 12950 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__11746_
timestamp 0
transform 1 0 12730 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11747_
timestamp 0
transform -1 0 12750 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11748_
timestamp 0
transform -1 0 12570 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11749_
timestamp 0
transform -1 0 14230 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11750_
timestamp 0
transform 1 0 12450 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__11751_
timestamp 0
transform 1 0 12730 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__11752_
timestamp 0
transform 1 0 16190 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11753_
timestamp 0
transform -1 0 16130 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__11754_
timestamp 0
transform -1 0 14750 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11755_
timestamp 0
transform 1 0 14970 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11756_
timestamp 0
transform 1 0 14830 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11757_
timestamp 0
transform -1 0 16290 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__11758_
timestamp 0
transform -1 0 15690 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__11759_
timestamp 0
transform 1 0 15790 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__11760_
timestamp 0
transform 1 0 14810 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__11761_
timestamp 0
transform 1 0 13190 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__11762_
timestamp 0
transform 1 0 13290 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__11763_
timestamp 0
transform 1 0 13050 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__11764_
timestamp 0
transform 1 0 13110 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__11765_
timestamp 0
transform 1 0 13350 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__11766_
timestamp 0
transform 1 0 13210 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__11767_
timestamp 0
transform -1 0 12890 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__11768_
timestamp 0
transform 1 0 12710 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__11769_
timestamp 0
transform 1 0 13110 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__11770_
timestamp 0
transform -1 0 12630 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11771_
timestamp 0
transform 1 0 12870 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11772_
timestamp 0
transform 1 0 14850 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__11773_
timestamp 0
transform -1 0 12430 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11774_
timestamp 0
transform -1 0 13270 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__11775_
timestamp 0
transform -1 0 12990 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__11776_
timestamp 0
transform 1 0 12570 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__11777_
timestamp 0
transform -1 0 12150 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__11778_
timestamp 0
transform -1 0 12410 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__11779_
timestamp 0
transform -1 0 13930 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__11780_
timestamp 0
transform -1 0 15210 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__11781_
timestamp 0
transform 1 0 15270 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__11782_
timestamp 0
transform -1 0 15050 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__11783_
timestamp 0
transform 1 0 12430 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__11784_
timestamp 0
transform -1 0 13150 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__11785_
timestamp 0
transform 1 0 13270 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__11786_
timestamp 0
transform -1 0 12850 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__11787_
timestamp 0
transform -1 0 13010 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__11788_
timestamp 0
transform 1 0 12810 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__11789_
timestamp 0
transform -1 0 13130 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__11790_
timestamp 0
transform -1 0 12290 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11791_
timestamp 0
transform -1 0 11990 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11792_
timestamp 0
transform 1 0 15590 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__11793_
timestamp 0
transform -1 0 15410 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__11794_
timestamp 0
transform -1 0 15550 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__11795_
timestamp 0
transform -1 0 15610 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__11796_
timestamp 0
transform -1 0 15130 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11797_
timestamp 0
transform 1 0 15250 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__11798_
timestamp 0
transform 1 0 15610 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__11799_
timestamp 0
transform -1 0 14790 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__11800_
timestamp 0
transform 1 0 15330 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__11801_
timestamp 0
transform -1 0 15490 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__11802_
timestamp 0
transform 1 0 13430 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__11803_
timestamp 0
transform -1 0 14890 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__11804_
timestamp 0
transform 1 0 15010 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__11805_
timestamp 0
transform -1 0 15170 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__11806_
timestamp 0
transform -1 0 15130 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__11807_
timestamp 0
transform -1 0 13390 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__11808_
timestamp 0
transform 1 0 15350 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__11809_
timestamp 0
transform -1 0 15470 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__11810_
timestamp 0
transform -1 0 15530 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__11811_
timestamp 0
transform 1 0 14610 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__11812_
timestamp 0
transform 1 0 13410 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__11813_
timestamp 0
transform -1 0 14530 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__11814_
timestamp 0
transform -1 0 14610 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__11815_
timestamp 0
transform 1 0 13250 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11816_
timestamp 0
transform -1 0 12990 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11817_
timestamp 0
transform -1 0 12350 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__11818_
timestamp 0
transform -1 0 13130 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11819_
timestamp 0
transform 1 0 12450 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__11820_
timestamp 0
transform -1 0 12630 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__11821_
timestamp 0
transform 1 0 12810 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__11822_
timestamp 0
transform -1 0 12670 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__11823_
timestamp 0
transform -1 0 12530 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__11824_
timestamp 0
transform 1 0 9330 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11825_
timestamp 0
transform -1 0 8710 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11826_
timestamp 0
transform -1 0 8830 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__11827_
timestamp 0
transform 1 0 12470 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11828_
timestamp 0
transform 1 0 12730 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11829_
timestamp 0
transform 1 0 15290 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__11830_
timestamp 0
transform 1 0 15130 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__11831_
timestamp 0
transform 1 0 14670 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__11832_
timestamp 0
transform 1 0 14910 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__11833_
timestamp 0
transform -1 0 14770 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__11834_
timestamp 0
transform -1 0 14790 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11835_
timestamp 0
transform -1 0 13750 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__11836_
timestamp 0
transform 1 0 13590 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__11837_
timestamp 0
transform 1 0 13530 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11838_
timestamp 0
transform 1 0 13530 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__11839_
timestamp 0
transform -1 0 13430 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11840_
timestamp 0
transform -1 0 13010 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__11841_
timestamp 0
transform 1 0 13130 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__11842_
timestamp 0
transform -1 0 13130 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__11843_
timestamp 0
transform 1 0 13210 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__11844_
timestamp 0
transform 1 0 13210 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11845_
timestamp 0
transform -1 0 13130 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11846_
timestamp 0
transform -1 0 12970 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__11847_
timestamp 0
transform -1 0 12990 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11848_
timestamp 0
transform 1 0 15330 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11849_
timestamp 0
transform -1 0 12770 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11850_
timestamp 0
transform -1 0 12610 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11851_
timestamp 0
transform 1 0 13050 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11852_
timestamp 0
transform 1 0 12890 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11853_
timestamp 0
transform 1 0 13370 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__11854_
timestamp 0
transform -1 0 13390 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11855_
timestamp 0
transform 1 0 16130 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__11856_
timestamp 0
transform 1 0 13870 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__11857_
timestamp 0
transform -1 0 14710 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__11858_
timestamp 0
transform 1 0 14350 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__11859_
timestamp 0
transform 1 0 14470 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__11860_
timestamp 0
transform -1 0 15610 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__11861_
timestamp 0
transform 1 0 15610 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11862_
timestamp 0
transform 1 0 16990 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__11863_
timestamp 0
transform 1 0 16410 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__11864_
timestamp 0
transform 1 0 15950 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__11865_
timestamp 0
transform 1 0 15890 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11866_
timestamp 0
transform 1 0 15750 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11867_
timestamp 0
transform 1 0 17050 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__11868_
timestamp 0
transform 1 0 16670 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11869_
timestamp 0
transform 1 0 16750 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__11870_
timestamp 0
transform -1 0 15790 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11871_
timestamp 0
transform -1 0 15650 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11872_
timestamp 0
transform -1 0 14890 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11873_
timestamp 0
transform 1 0 14750 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11874_
timestamp 0
transform -1 0 13630 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11875_
timestamp 0
transform -1 0 13490 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11876_
timestamp 0
transform 1 0 13210 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11877_
timestamp 0
transform 1 0 15130 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11878_
timestamp 0
transform -1 0 17050 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11879_
timestamp 0
transform 1 0 14390 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__11880_
timestamp 0
transform 1 0 14650 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__11881_
timestamp 0
transform 1 0 14430 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__11882_
timestamp 0
transform -1 0 15490 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__11883_
timestamp 0
transform -1 0 15750 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__11884_
timestamp 0
transform -1 0 15770 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11885_
timestamp 0
transform -1 0 16070 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11886_
timestamp 0
transform -1 0 16790 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11887_
timestamp 0
transform 1 0 16830 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11888_
timestamp 0
transform 1 0 16930 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11889_
timestamp 0
transform 1 0 16710 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11890_
timestamp 0
transform 1 0 16710 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11891_
timestamp 0
transform 1 0 16770 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11892_
timestamp 0
transform -1 0 16870 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11893_
timestamp 0
transform -1 0 16990 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11894_
timestamp 0
transform 1 0 16970 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11895_
timestamp 0
transform 1 0 17030 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11896_
timestamp 0
transform -1 0 15450 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11897_
timestamp 0
transform -1 0 15310 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11898_
timestamp 0
transform 1 0 13970 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11899_
timestamp 0
transform 1 0 16290 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11900_
timestamp 0
transform -1 0 16910 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__11901_
timestamp 0
transform 1 0 16910 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__11902_
timestamp 0
transform -1 0 14670 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11903_
timestamp 0
transform 1 0 14930 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11904_
timestamp 0
transform 1 0 15330 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11905_
timestamp 0
transform 1 0 15470 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11906_
timestamp 0
transform 1 0 15550 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__11907_
timestamp 0
transform 1 0 16570 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11908_
timestamp 0
transform -1 0 16530 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__11909_
timestamp 0
transform 1 0 16470 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11910_
timestamp 0
transform -1 0 16330 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11911_
timestamp 0
transform -1 0 16330 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11912_
timestamp 0
transform 1 0 16450 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11913_
timestamp 0
transform 1 0 16770 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11914_
timestamp 0
transform 1 0 16650 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11915_
timestamp 0
transform -1 0 15150 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11916_
timestamp 0
transform -1 0 15010 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11917_
timestamp 0
transform -1 0 14690 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11918_
timestamp 0
transform 1 0 12530 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11919_
timestamp 0
transform 1 0 14390 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11920_
timestamp 0
transform -1 0 16390 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__11921_
timestamp 0
transform 1 0 16570 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11922_
timestamp 0
transform -1 0 15190 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11923_
timestamp 0
transform -1 0 15190 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__11924_
timestamp 0
transform 1 0 15250 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__11925_
timestamp 0
transform -1 0 16050 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11926_
timestamp 0
transform 1 0 16050 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11927_
timestamp 0
transform 1 0 16410 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11928_
timestamp 0
transform 1 0 16150 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11929_
timestamp 0
transform -1 0 16170 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11930_
timestamp 0
transform -1 0 15910 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11931_
timestamp 0
transform 1 0 16270 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11932_
timestamp 0
transform 1 0 15910 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11933_
timestamp 0
transform 1 0 16050 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11934_
timestamp 0
transform -1 0 16630 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11935_
timestamp 0
transform 1 0 16850 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11936_
timestamp 0
transform 1 0 16870 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11937_
timestamp 0
transform 1 0 16530 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11938_
timestamp 0
transform -1 0 15750 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11939_
timestamp 0
transform -1 0 15610 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11940_
timestamp 0
transform 1 0 14510 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11941_
timestamp 0
transform 1 0 12830 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11942_
timestamp 0
transform -1 0 16030 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11943_
timestamp 0
transform 1 0 16970 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11944_
timestamp 0
transform 1 0 16710 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11945_
timestamp 0
transform -1 0 16590 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11946_
timestamp 0
transform 1 0 16410 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11947_
timestamp 0
transform -1 0 15970 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11948_
timestamp 0
transform -1 0 16270 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__11949_
timestamp 0
transform -1 0 16190 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11950_
timestamp 0
transform 1 0 14530 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__11951_
timestamp 0
transform -1 0 15310 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__11952_
timestamp 0
transform 1 0 15410 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__11953_
timestamp 0
transform 1 0 15850 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__11954_
timestamp 0
transform 1 0 15710 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11955_
timestamp 0
transform 1 0 16550 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11956_
timestamp 0
transform 1 0 16370 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__11957_
timestamp 0
transform 1 0 16290 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11958_
timestamp 0
transform 1 0 15850 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11959_
timestamp 0
transform -1 0 16170 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11960_
timestamp 0
transform -1 0 16430 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11961_
timestamp 0
transform -1 0 16030 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__11962_
timestamp 0
transform 1 0 15810 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11963_
timestamp 0
transform 1 0 15590 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11964_
timestamp 0
transform 1 0 15690 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11965_
timestamp 0
transform 1 0 15890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11966_
timestamp 0
transform -1 0 15470 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11967_
timestamp 0
transform -1 0 13230 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__11968_
timestamp 0
transform 1 0 13770 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11969_
timestamp 0
transform -1 0 14330 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11970_
timestamp 0
transform 1 0 12950 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11971_
timestamp 0
transform 1 0 14050 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11972_
timestamp 0
transform 1 0 16090 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11973_
timestamp 0
transform 1 0 16170 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__11974_
timestamp 0
transform 1 0 16250 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11975_
timestamp 0
transform 1 0 15390 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11976_
timestamp 0
transform -1 0 15690 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__11977_
timestamp 0
transform -1 0 15710 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__11978_
timestamp 0
transform -1 0 15550 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__11979_
timestamp 0
transform 1 0 15970 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__11980_
timestamp 0
transform 1 0 15350 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11981_
timestamp 0
transform -1 0 15610 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11982_
timestamp 0
transform -1 0 15230 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11983_
timestamp 0
transform 1 0 15450 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11984_
timestamp 0
transform -1 0 15830 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__11985_
timestamp 0
transform 1 0 15490 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11986_
timestamp 0
transform 1 0 15230 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11987_
timestamp 0
transform 1 0 15230 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11988_
timestamp 0
transform -1 0 15110 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11989_
timestamp 0
transform 1 0 14930 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11990_
timestamp 0
transform 1 0 14150 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__11991_
timestamp 0
transform -1 0 15730 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11992_
timestamp 0
transform -1 0 15450 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11993_
timestamp 0
transform -1 0 15870 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11994_
timestamp 0
transform -1 0 15590 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11995_
timestamp 0
transform -1 0 15310 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11996_
timestamp 0
transform -1 0 15130 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__11997_
timestamp 0
transform -1 0 15010 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__11998_
timestamp 0
transform 1 0 14650 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__11999_
timestamp 0
transform -1 0 15510 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__12000_
timestamp 0
transform -1 0 15290 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__12001_
timestamp 0
transform -1 0 15430 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12002_
timestamp 0
transform -1 0 15150 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__12003_
timestamp 0
transform -1 0 15110 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__12004_
timestamp 0
transform -1 0 15090 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__12005_
timestamp 0
transform 1 0 14770 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__12006_
timestamp 0
transform 1 0 14990 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__12007_
timestamp 0
transform -1 0 15410 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__12008_
timestamp 0
transform 1 0 14670 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__12009_
timestamp 0
transform 1 0 14810 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__12010_
timestamp 0
transform -1 0 14790 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__12011_
timestamp 0
transform -1 0 14650 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__12012_
timestamp 0
transform -1 0 14490 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__12013_
timestamp 0
transform 1 0 13430 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__12014_
timestamp 0
transform 1 0 14630 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__12015_
timestamp 0
transform 1 0 15090 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12016_
timestamp 0
transform -1 0 14750 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__12017_
timestamp 0
transform -1 0 14850 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__12018_
timestamp 0
transform -1 0 14850 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__12019_
timestamp 0
transform 1 0 14550 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__12020_
timestamp 0
transform 1 0 14490 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__12021_
timestamp 0
transform -1 0 14430 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__12022_
timestamp 0
transform 1 0 14270 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__12023_
timestamp 0
transform -1 0 14270 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__12024_
timestamp 0
transform -1 0 14510 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__12025_
timestamp 0
transform -1 0 14150 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__12026_
timestamp 0
transform -1 0 14370 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__12027_
timestamp 0
transform -1 0 14330 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__12028_
timestamp 0
transform 1 0 14930 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__12029_
timestamp 0
transform -1 0 14970 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__12030_
timestamp 0
transform -1 0 14630 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__12031_
timestamp 0
transform -1 0 14470 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__12032_
timestamp 0
transform 1 0 14370 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__12033_
timestamp 0
transform -1 0 14690 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__12034_
timestamp 0
transform -1 0 14530 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__12035_
timestamp 0
transform 1 0 14230 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__12036_
timestamp 0
transform -1 0 14050 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__12037_
timestamp 0
transform 1 0 13870 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__12038_
timestamp 0
transform -1 0 13010 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__12039_
timestamp 0
transform -1 0 14210 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__12040_
timestamp 0
transform 1 0 14650 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12041_
timestamp 0
transform 1 0 14770 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12042_
timestamp 0
transform -1 0 14410 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12043_
timestamp 0
transform -1 0 14530 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12044_
timestamp 0
transform 1 0 14190 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12045_
timestamp 0
transform -1 0 14170 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__12046_
timestamp 0
transform -1 0 14030 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__12047_
timestamp 0
transform -1 0 13910 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__12048_
timestamp 0
transform 1 0 13790 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__12049_
timestamp 0
transform -1 0 13930 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__12050_
timestamp 0
transform -1 0 14110 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__12051_
timestamp 0
transform -1 0 13650 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__12052_
timestamp 0
transform -1 0 13510 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__12053_
timestamp 0
transform 1 0 13350 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__12054_
timestamp 0
transform 1 0 12830 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12055_
timestamp 0
transform -1 0 15810 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12056_
timestamp 0
transform 1 0 16010 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12057_
timestamp 0
transform 1 0 15910 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12058_
timestamp 0
transform -1 0 16010 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12059_
timestamp 0
transform -1 0 12550 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12060_
timestamp 0
transform 1 0 12830 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12061_
timestamp 0
transform -1 0 12590 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12062_
timestamp 0
transform 1 0 16130 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12063_
timestamp 0
transform 1 0 16470 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12064_
timestamp 0
transform -1 0 16610 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12065_
timestamp 0
transform -1 0 17030 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12066_
timestamp 0
transform 1 0 17010 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12067_
timestamp 0
transform 1 0 16690 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12068_
timestamp 0
transform 1 0 16650 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12069_
timestamp 0
transform -1 0 16230 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12070_
timestamp 0
transform 1 0 12830 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12071_
timestamp 0
transform 1 0 17010 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12072_
timestamp 0
transform -1 0 16890 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12073_
timestamp 0
transform 1 0 17050 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12074_
timestamp 0
transform -1 0 16910 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12075_
timestamp 0
transform -1 0 12990 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12076_
timestamp 0
transform -1 0 12710 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12077_
timestamp 0
transform -1 0 12550 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12078_
timestamp 0
transform -1 0 13130 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12079_
timestamp 0
transform 1 0 15550 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__12080_
timestamp 0
transform 1 0 16970 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12081_
timestamp 0
transform 1 0 13770 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12082_
timestamp 0
transform 1 0 13630 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12083_
timestamp 0
transform -1 0 16710 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12084_
timestamp 0
transform 1 0 16550 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12085_
timestamp 0
transform -1 0 16070 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12086_
timestamp 0
transform -1 0 16190 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12087_
timestamp 0
transform -1 0 16690 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12088_
timestamp 0
transform 1 0 16450 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12089_
timestamp 0
transform 1 0 16730 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12090_
timestamp 0
transform 1 0 16950 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12091_
timestamp 0
transform 1 0 16770 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12092_
timestamp 0
transform 1 0 16530 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12093_
timestamp 0
transform -1 0 15410 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12094_
timestamp 0
transform 1 0 16690 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12095_
timestamp 0
transform -1 0 16550 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12096_
timestamp 0
transform 1 0 16350 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12097_
timestamp 0
transform -1 0 15130 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12098_
timestamp 0
transform -1 0 15150 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12099_
timestamp 0
transform 1 0 15250 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12100_
timestamp 0
transform -1 0 15010 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12101_
timestamp 0
transform 1 0 13770 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12102_
timestamp 0
transform -1 0 13650 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12103_
timestamp 0
transform -1 0 13490 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12104_
timestamp 0
transform -1 0 12690 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12105_
timestamp 0
transform -1 0 13150 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12106_
timestamp 0
transform 1 0 15250 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12107_
timestamp 0
transform -1 0 16810 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12108_
timestamp 0
transform -1 0 15530 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12109_
timestamp 0
transform -1 0 15670 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12110_
timestamp 0
transform 1 0 16550 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12111_
timestamp 0
transform 1 0 16130 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12112_
timestamp 0
transform -1 0 16310 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12113_
timestamp 0
transform 1 0 16870 0 1 250
box -6 -8 26 248
use FILL  FILL_0__12114_
timestamp 0
transform -1 0 16450 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12115_
timestamp 0
transform 1 0 16350 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12116_
timestamp 0
transform 1 0 16910 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12117_
timestamp 0
transform -1 0 16770 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12118_
timestamp 0
transform 1 0 16510 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12119_
timestamp 0
transform 1 0 16610 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12120_
timestamp 0
transform 1 0 16450 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12121_
timestamp 0
transform -1 0 16070 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12122_
timestamp 0
transform 1 0 16290 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12123_
timestamp 0
transform -1 0 15950 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12124_
timestamp 0
transform -1 0 15670 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12125_
timestamp 0
transform 1 0 15810 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12126_
timestamp 0
transform -1 0 15530 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12127_
timestamp 0
transform -1 0 13290 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12128_
timestamp 0
transform 1 0 16150 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12129_
timestamp 0
transform 1 0 17010 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12130_
timestamp 0
transform -1 0 14990 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__12131_
timestamp 0
transform 1 0 15350 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__12132_
timestamp 0
transform -1 0 16230 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12133_
timestamp 0
transform -1 0 16790 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12134_
timestamp 0
transform 1 0 16850 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12135_
timestamp 0
transform 1 0 16990 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12136_
timestamp 0
transform 1 0 16850 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12137_
timestamp 0
transform 1 0 16890 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12138_
timestamp 0
transform 1 0 17010 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12139_
timestamp 0
transform 1 0 17030 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12140_
timestamp 0
transform 1 0 16750 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12141_
timestamp 0
transform -1 0 16530 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12142_
timestamp 0
transform 1 0 16510 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12143_
timestamp 0
transform 1 0 16670 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12144_
timestamp 0
transform 1 0 16610 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12145_
timestamp 0
transform 1 0 16870 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12146_
timestamp 0
transform 1 0 16730 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12147_
timestamp 0
transform 1 0 16830 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12148_
timestamp 0
transform 1 0 14350 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12149_
timestamp 0
transform 1 0 16370 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12150_
timestamp 0
transform -1 0 14910 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12151_
timestamp 0
transform 1 0 15010 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12152_
timestamp 0
transform -1 0 15630 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12153_
timestamp 0
transform -1 0 15850 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12154_
timestamp 0
transform -1 0 16530 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12155_
timestamp 0
transform 1 0 16630 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12156_
timestamp 0
transform 1 0 17070 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12157_
timestamp 0
transform 1 0 16910 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12158_
timestamp 0
transform 1 0 16970 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12159_
timestamp 0
transform -1 0 16850 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12160_
timestamp 0
transform 1 0 16830 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12161_
timestamp 0
transform 1 0 16690 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12162_
timestamp 0
transform 1 0 16690 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12163_
timestamp 0
transform 1 0 16970 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12164_
timestamp 0
transform -1 0 16570 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12165_
timestamp 0
transform -1 0 16550 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12166_
timestamp 0
transform -1 0 16130 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12167_
timestamp 0
transform -1 0 15330 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12168_
timestamp 0
transform 1 0 15470 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12169_
timestamp 0
transform 1 0 15190 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12170_
timestamp 0
transform 1 0 13770 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12171_
timestamp 0
transform 1 0 13950 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12172_
timestamp 0
transform 1 0 15830 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12173_
timestamp 0
transform -1 0 16110 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12174_
timestamp 0
transform -1 0 15950 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12175_
timestamp 0
transform 1 0 16070 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12176_
timestamp 0
transform 1 0 16430 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12177_
timestamp 0
transform 1 0 16270 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12178_
timestamp 0
transform 1 0 16130 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12179_
timestamp 0
transform 1 0 16210 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12180_
timestamp 0
transform -1 0 16650 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12181_
timestamp 0
transform -1 0 16510 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12182_
timestamp 0
transform -1 0 16370 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12183_
timestamp 0
transform -1 0 16250 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12184_
timestamp 0
transform -1 0 16250 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12185_
timestamp 0
transform -1 0 15990 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12186_
timestamp 0
transform -1 0 16410 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12187_
timestamp 0
transform -1 0 15450 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12188_
timestamp 0
transform 1 0 15070 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12189_
timestamp 0
transform -1 0 14930 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12190_
timestamp 0
transform -1 0 14790 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12191_
timestamp 0
transform 1 0 14050 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12192_
timestamp 0
transform 1 0 12630 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12193_
timestamp 0
transform -1 0 15950 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12194_
timestamp 0
transform 1 0 15990 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12195_
timestamp 0
transform -1 0 16110 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12196_
timestamp 0
transform -1 0 16210 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12197_
timestamp 0
transform 1 0 15630 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12198_
timestamp 0
transform -1 0 16270 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12199_
timestamp 0
transform 1 0 15890 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12200_
timestamp 0
transform -1 0 16010 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12201_
timestamp 0
transform 1 0 15370 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12202_
timestamp 0
transform 1 0 15250 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12203_
timestamp 0
transform 1 0 15090 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12204_
timestamp 0
transform -1 0 14990 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12205_
timestamp 0
transform -1 0 16390 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12206_
timestamp 0
transform -1 0 16010 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12207_
timestamp 0
transform 1 0 15690 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12208_
timestamp 0
transform 1 0 15550 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12209_
timestamp 0
transform 1 0 15310 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12210_
timestamp 0
transform -1 0 15170 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12211_
timestamp 0
transform -1 0 16250 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12212_
timestamp 0
transform -1 0 15850 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12213_
timestamp 0
transform -1 0 16090 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12214_
timestamp 0
transform -1 0 15710 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12215_
timestamp 0
transform -1 0 15030 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12216_
timestamp 0
transform -1 0 14890 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12217_
timestamp 0
transform 1 0 13110 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12218_
timestamp 0
transform 1 0 12970 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12219_
timestamp 0
transform 1 0 13950 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12220_
timestamp 0
transform -1 0 14770 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12221_
timestamp 0
transform 1 0 16130 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12222_
timestamp 0
transform 1 0 15790 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12223_
timestamp 0
transform -1 0 15750 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12224_
timestamp 0
transform -1 0 15950 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12225_
timestamp 0
transform 1 0 15450 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12226_
timestamp 0
transform 1 0 15790 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12227_
timestamp 0
transform -1 0 15790 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12228_
timestamp 0
transform -1 0 15570 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12229_
timestamp 0
transform -1 0 15410 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12230_
timestamp 0
transform -1 0 15870 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12231_
timestamp 0
transform -1 0 15690 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12232_
timestamp 0
transform -1 0 15710 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12233_
timestamp 0
transform 1 0 15510 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12234_
timestamp 0
transform -1 0 14490 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12235_
timestamp 0
transform 1 0 14630 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12236_
timestamp 0
transform -1 0 14370 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12237_
timestamp 0
transform -1 0 14230 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12238_
timestamp 0
transform 1 0 14050 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__12239_
timestamp 0
transform 1 0 14810 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12240_
timestamp 0
transform -1 0 14710 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12241_
timestamp 0
transform -1 0 14550 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12242_
timestamp 0
transform -1 0 14410 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12243_
timestamp 0
transform 1 0 15990 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12244_
timestamp 0
transform -1 0 16090 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12245_
timestamp 0
transform -1 0 15950 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12246_
timestamp 0
transform -1 0 15190 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12247_
timestamp 0
transform -1 0 14810 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12248_
timestamp 0
transform -1 0 15310 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12249_
timestamp 0
transform -1 0 15070 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12250_
timestamp 0
transform -1 0 14510 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12251_
timestamp 0
transform -1 0 15210 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12252_
timestamp 0
transform 1 0 14930 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12253_
timestamp 0
transform -1 0 14650 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12254_
timestamp 0
transform -1 0 14130 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12255_
timestamp 0
transform -1 0 13730 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12256_
timestamp 0
transform -1 0 14270 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12257_
timestamp 0
transform -1 0 13850 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12258_
timestamp 0
transform 1 0 13530 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12259_
timestamp 0
transform -1 0 13470 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12260_
timestamp 0
transform -1 0 13990 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12261_
timestamp 0
transform -1 0 14070 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12262_
timestamp 0
transform 1 0 15790 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12263_
timestamp 0
transform 1 0 14870 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12264_
timestamp 0
transform -1 0 15070 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12265_
timestamp 0
transform 1 0 14910 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12266_
timestamp 0
transform -1 0 14790 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12267_
timestamp 0
transform -1 0 14510 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12268_
timestamp 0
transform 1 0 14650 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12269_
timestamp 0
transform 1 0 14610 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12270_
timestamp 0
transform 1 0 14250 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12271_
timestamp 0
transform -1 0 13970 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12272_
timestamp 0
transform 1 0 14090 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12273_
timestamp 0
transform -1 0 13830 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12274_
timestamp 0
transform 1 0 13370 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12275_
timestamp 0
transform -1 0 14190 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12276_
timestamp 0
transform 1 0 14290 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12277_
timestamp 0
transform -1 0 14410 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12278_
timestamp 0
transform 1 0 14590 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12279_
timestamp 0
transform -1 0 14450 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12280_
timestamp 0
transform 1 0 15650 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12281_
timestamp 0
transform -1 0 15570 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12282_
timestamp 0
transform 1 0 15350 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12283_
timestamp 0
transform -1 0 14750 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12284_
timestamp 0
transform 1 0 14470 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12285_
timestamp 0
transform -1 0 14570 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12286_
timestamp 0
transform 1 0 14390 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12287_
timestamp 0
transform -1 0 14230 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12288_
timestamp 0
transform 1 0 14350 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12289_
timestamp 0
transform -1 0 14070 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12290_
timestamp 0
transform 1 0 14250 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12291_
timestamp 0
transform -1 0 13790 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12292_
timestamp 0
transform 1 0 13930 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12293_
timestamp 0
transform -1 0 13670 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12294_
timestamp 0
transform 1 0 13470 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12295_
timestamp 0
transform -1 0 13110 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12296_
timestamp 0
transform -1 0 14390 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12297_
timestamp 0
transform -1 0 14130 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12298_
timestamp 0
transform 1 0 14250 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12299_
timestamp 0
transform 1 0 14130 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12300_
timestamp 0
transform 1 0 14250 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12301_
timestamp 0
transform -1 0 14130 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12302_
timestamp 0
transform -1 0 13990 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12303_
timestamp 0
transform -1 0 13830 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12304_
timestamp 0
transform -1 0 13690 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12305_
timestamp 0
transform -1 0 11870 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12306_
timestamp 0
transform 1 0 10670 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12307_
timestamp 0
transform 1 0 10810 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12308_
timestamp 0
transform -1 0 10930 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12309_
timestamp 0
transform 1 0 11050 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12310_
timestamp 0
transform 1 0 11170 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12311_
timestamp 0
transform 1 0 11490 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12312_
timestamp 0
transform 1 0 11250 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12313_
timestamp 0
transform -1 0 11250 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12314_
timestamp 0
transform -1 0 10930 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12315_
timestamp 0
transform 1 0 10710 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12316_
timestamp 0
transform -1 0 10590 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12317_
timestamp 0
transform -1 0 10030 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12318_
timestamp 0
transform -1 0 10310 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12319_
timestamp 0
transform -1 0 10170 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12320_
timestamp 0
transform 1 0 10230 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12321_
timestamp 0
transform -1 0 10190 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12322_
timestamp 0
transform -1 0 10090 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12323_
timestamp 0
transform -1 0 10070 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12324_
timestamp 0
transform -1 0 10850 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12325_
timestamp 0
transform -1 0 10710 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12326_
timestamp 0
transform -1 0 10970 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12327_
timestamp 0
transform 1 0 11070 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12328_
timestamp 0
transform 1 0 10430 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12329_
timestamp 0
transform 1 0 10530 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12330_
timestamp 0
transform -1 0 12450 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12331_
timestamp 0
transform -1 0 11510 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12332_
timestamp 0
transform -1 0 11650 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12333_
timestamp 0
transform 1 0 11210 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12334_
timestamp 0
transform -1 0 11070 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12335_
timestamp 0
transform 1 0 10930 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12336_
timestamp 0
transform -1 0 10830 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12337_
timestamp 0
transform -1 0 10330 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12338_
timestamp 0
transform -1 0 10390 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12339_
timestamp 0
transform 1 0 10230 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12340_
timestamp 0
transform 1 0 10070 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12341_
timestamp 0
transform 1 0 11130 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12342_
timestamp 0
transform -1 0 10630 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12343_
timestamp 0
transform 1 0 10990 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12344_
timestamp 0
transform 1 0 11630 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12345_
timestamp 0
transform 1 0 12590 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12346_
timestamp 0
transform -1 0 12310 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12347_
timestamp 0
transform 1 0 11910 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12348_
timestamp 0
transform -1 0 12010 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12349_
timestamp 0
transform 1 0 11510 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12350_
timestamp 0
transform -1 0 11410 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12351_
timestamp 0
transform -1 0 10610 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12352_
timestamp 0
transform -1 0 10730 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12353_
timestamp 0
transform 1 0 11090 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12354_
timestamp 0
transform 1 0 11110 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12355_
timestamp 0
transform -1 0 11030 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12356_
timestamp 0
transform 1 0 10630 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12357_
timestamp 0
transform -1 0 9930 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12358_
timestamp 0
transform -1 0 10450 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12359_
timestamp 0
transform -1 0 10310 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12360_
timestamp 0
transform -1 0 10010 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12361_
timestamp 0
transform -1 0 9670 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12362_
timestamp 0
transform -1 0 9810 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12363_
timestamp 0
transform -1 0 9750 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12364_
timestamp 0
transform -1 0 10870 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12365_
timestamp 0
transform 1 0 9930 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12366_
timestamp 0
transform 1 0 10090 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12367_
timestamp 0
transform 1 0 10230 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12368_
timestamp 0
transform -1 0 9530 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12369_
timestamp 0
transform -1 0 9910 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12370_
timestamp 0
transform 1 0 12650 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12371_
timestamp 0
transform 1 0 12010 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12372_
timestamp 0
transform 1 0 12150 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12373_
timestamp 0
transform -1 0 12330 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12374_
timestamp 0
transform -1 0 10170 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12375_
timestamp 0
transform -1 0 10210 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12376_
timestamp 0
transform 1 0 10250 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12377_
timestamp 0
transform 1 0 9870 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12378_
timestamp 0
transform -1 0 9270 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12379_
timestamp 0
transform -1 0 9390 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12380_
timestamp 0
transform -1 0 9490 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12381_
timestamp 0
transform -1 0 9330 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12382_
timestamp 0
transform 1 0 10630 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12383_
timestamp 0
transform 1 0 9650 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12384_
timestamp 0
transform 1 0 9750 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12385_
timestamp 0
transform 1 0 10010 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12386_
timestamp 0
transform -1 0 9910 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12387_
timestamp 0
transform -1 0 9730 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12388_
timestamp 0
transform -1 0 12470 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12389_
timestamp 0
transform 1 0 12450 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12390_
timestamp 0
transform 1 0 12170 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12391_
timestamp 0
transform -1 0 12310 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12392_
timestamp 0
transform -1 0 12070 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12393_
timestamp 0
transform 1 0 10990 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12394_
timestamp 0
transform -1 0 10850 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12395_
timestamp 0
transform 1 0 10830 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12396_
timestamp 0
transform -1 0 10010 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12397_
timestamp 0
transform -1 0 10030 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12398_
timestamp 0
transform -1 0 9890 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12399_
timestamp 0
transform -1 0 10150 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12400_
timestamp 0
transform 1 0 10250 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12401_
timestamp 0
transform 1 0 10350 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12402_
timestamp 0
transform 1 0 10710 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12403_
timestamp 0
transform 1 0 11290 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12404_
timestamp 0
transform -1 0 10530 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12405_
timestamp 0
transform -1 0 10390 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12406_
timestamp 0
transform 1 0 10630 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12407_
timestamp 0
transform -1 0 10790 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12408_
timestamp 0
transform -1 0 10590 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12409_
timestamp 0
transform -1 0 10910 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12410_
timestamp 0
transform -1 0 10450 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12411_
timestamp 0
transform 1 0 10570 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12412_
timestamp 0
transform -1 0 10450 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12413_
timestamp 0
transform 1 0 10470 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12414_
timestamp 0
transform 1 0 11110 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12415_
timestamp 0
transform 1 0 11850 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12416_
timestamp 0
transform -1 0 11770 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12417_
timestamp 0
transform -1 0 11630 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12418_
timestamp 0
transform 1 0 11610 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12419_
timestamp 0
transform 1 0 11770 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12420_
timestamp 0
transform -1 0 11730 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12421_
timestamp 0
transform -1 0 10310 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12422_
timestamp 0
transform -1 0 10310 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12423_
timestamp 0
transform 1 0 10150 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12424_
timestamp 0
transform 1 0 9990 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12425_
timestamp 0
transform 1 0 10130 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12426_
timestamp 0
transform 1 0 11230 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12427_
timestamp 0
transform -1 0 11070 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12428_
timestamp 0
transform -1 0 10950 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12429_
timestamp 0
transform 1 0 10950 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12430_
timestamp 0
transform -1 0 11630 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12431_
timestamp 0
transform -1 0 11730 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12432_
timestamp 0
transform -1 0 11590 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12433_
timestamp 0
transform -1 0 11210 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12434_
timestamp 0
transform -1 0 11210 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12435_
timestamp 0
transform 1 0 11350 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12436_
timestamp 0
transform -1 0 11330 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12437_
timestamp 0
transform -1 0 11770 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12438_
timestamp 0
transform 1 0 11470 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12439_
timestamp 0
transform -1 0 11330 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12440_
timestamp 0
transform -1 0 11370 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12441_
timestamp 0
transform 1 0 11450 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12442_
timestamp 0
transform -1 0 12130 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12443_
timestamp 0
transform 1 0 12170 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12444_
timestamp 0
transform -1 0 11990 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12445_
timestamp 0
transform 1 0 12350 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12446_
timestamp 0
transform -1 0 12070 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12447_
timestamp 0
transform -1 0 12010 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12448_
timestamp 0
transform -1 0 11910 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12449_
timestamp 0
transform 1 0 12170 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12450_
timestamp 0
transform 1 0 12210 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__12451_
timestamp 0
transform 1 0 12010 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__12452_
timestamp 0
transform 1 0 11750 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__12453_
timestamp 0
transform -1 0 11670 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__12454_
timestamp 0
transform 1 0 11790 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__12455_
timestamp 0
transform -1 0 13850 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12456_
timestamp 0
transform -1 0 13970 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12457_
timestamp 0
transform -1 0 13930 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12458_
timestamp 0
transform -1 0 14050 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12459_
timestamp 0
transform 1 0 14010 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12460_
timestamp 0
transform -1 0 11690 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__12461_
timestamp 0
transform 1 0 13970 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12462_
timestamp 0
transform 1 0 13830 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12463_
timestamp 0
transform 1 0 14110 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12464_
timestamp 0
transform 1 0 13690 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12465_
timestamp 0
transform -1 0 13530 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12466_
timestamp 0
transform 1 0 12270 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12467_
timestamp 0
transform -1 0 14790 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12468_
timestamp 0
transform 1 0 14230 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12469_
timestamp 0
transform 1 0 14310 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12470_
timestamp 0
transform 1 0 13910 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12471_
timestamp 0
transform 1 0 12150 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12472_
timestamp 0
transform 1 0 16390 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__12473_
timestamp 0
transform -1 0 16550 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__12474_
timestamp 0
transform 1 0 15150 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__12475_
timestamp 0
transform -1 0 15530 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__12476_
timestamp 0
transform 1 0 13530 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12477_
timestamp 0
transform -1 0 13690 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12478_
timestamp 0
transform 1 0 13590 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12479_
timestamp 0
transform -1 0 13750 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__12480_
timestamp 0
transform -1 0 12870 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12481_
timestamp 0
transform 1 0 12970 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12482_
timestamp 0
transform 1 0 13630 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12483_
timestamp 0
transform 1 0 13490 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12484_
timestamp 0
transform -1 0 13990 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__12485_
timestamp 0
transform -1 0 14130 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__12486_
timestamp 0
transform 1 0 14130 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12487_
timestamp 0
transform -1 0 14270 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12488_
timestamp 0
transform -1 0 13890 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__12489_
timestamp 0
transform -1 0 13730 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__12490_
timestamp 0
transform 1 0 13570 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__12491_
timestamp 0
transform -1 0 14030 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12492_
timestamp 0
transform 1 0 13370 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__12493_
timestamp 0
transform -1 0 13530 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__12494_
timestamp 0
transform -1 0 14450 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12495_
timestamp 0
transform 1 0 14050 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12496_
timestamp 0
transform -1 0 14730 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12497_
timestamp 0
transform 1 0 14570 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12498_
timestamp 0
transform 1 0 16330 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12499_
timestamp 0
transform -1 0 16590 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12500_
timestamp 0
transform 1 0 16490 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12501_
timestamp 0
transform -1 0 16630 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12502_
timestamp 0
transform -1 0 13310 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12503_
timestamp 0
transform -1 0 13450 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12504_
timestamp 0
transform 1 0 13530 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12505_
timestamp 0
transform -1 0 13690 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12506_
timestamp 0
transform -1 0 12070 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12507_
timestamp 0
transform -1 0 12210 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12508_
timestamp 0
transform -1 0 11770 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12509_
timestamp 0
transform -1 0 11910 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12510_
timestamp 0
transform 1 0 12430 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12511_
timestamp 0
transform 1 0 12290 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__12512_
timestamp 0
transform 1 0 11850 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12513_
timestamp 0
transform -1 0 11930 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__12514_
timestamp 0
transform 1 0 12030 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12515_
timestamp 0
transform -1 0 12290 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12516_
timestamp 0
transform 1 0 12130 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12517_
timestamp 0
transform 1 0 11650 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12518_
timestamp 0
transform -1 0 12130 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12519_
timestamp 0
transform 1 0 11970 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12520_
timestamp 0
transform 1 0 10970 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12521_
timestamp 0
transform -1 0 11130 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__12522_
timestamp 0
transform 1 0 11370 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12523_
timestamp 0
transform -1 0 11530 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__12524_
timestamp 0
transform -1 0 9390 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12525_
timestamp 0
transform -1 0 9510 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__12526_
timestamp 0
transform -1 0 9630 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12527_
timestamp 0
transform -1 0 9750 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__12528_
timestamp 0
transform 1 0 11330 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12529_
timestamp 0
transform -1 0 11730 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__12530_
timestamp 0
transform -1 0 11570 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12531_
timestamp 0
transform -1 0 11730 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__12532_
timestamp 0
transform 1 0 11150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12533_
timestamp 0
transform 1 0 11010 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12534_
timestamp 0
transform 1 0 10770 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12535_
timestamp 0
transform -1 0 10650 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__12616_
timestamp 0
transform 1 0 11250 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12617_
timestamp 0
transform -1 0 11370 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12618_
timestamp 0
transform 1 0 12330 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12619_
timestamp 0
transform 1 0 11470 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12620_
timestamp 0
transform -1 0 11070 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12621_
timestamp 0
transform -1 0 10810 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12622_
timestamp 0
transform 1 0 10910 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12623_
timestamp 0
transform -1 0 11030 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12624_
timestamp 0
transform -1 0 11510 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12625_
timestamp 0
transform -1 0 11690 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12626_
timestamp 0
transform -1 0 11530 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12627_
timestamp 0
transform -1 0 10590 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__12628_
timestamp 0
transform -1 0 11490 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12629_
timestamp 0
transform 1 0 11310 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12630_
timestamp 0
transform -1 0 11190 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12631_
timestamp 0
transform 1 0 11170 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12632_
timestamp 0
transform 1 0 11130 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12633_
timestamp 0
transform 1 0 11610 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12634_
timestamp 0
transform -1 0 11130 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12635_
timestamp 0
transform -1 0 11270 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12636_
timestamp 0
transform -1 0 11610 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12637_
timestamp 0
transform -1 0 11790 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12638_
timestamp 0
transform 1 0 11610 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12639_
timestamp 0
transform -1 0 11230 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12640_
timestamp 0
transform -1 0 11630 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__12641_
timestamp 0
transform -1 0 11290 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12642_
timestamp 0
transform 1 0 10930 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__12643_
timestamp 0
transform -1 0 11290 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__12644_
timestamp 0
transform -1 0 10990 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__12645_
timestamp 0
transform -1 0 11130 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12646_
timestamp 0
transform -1 0 11510 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12647_
timestamp 0
transform 1 0 11350 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12648_
timestamp 0
transform 1 0 11050 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12649_
timestamp 0
transform 1 0 11390 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12650_
timestamp 0
transform -1 0 10910 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12651_
timestamp 0
transform -1 0 10430 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__12652_
timestamp 0
transform 1 0 11110 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__12653_
timestamp 0
transform 1 0 11170 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12654_
timestamp 0
transform -1 0 11470 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__12655_
timestamp 0
transform 1 0 11170 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__12656_
timestamp 0
transform -1 0 11330 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__12657_
timestamp 0
transform 1 0 11310 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12658_
timestamp 0
transform 1 0 12070 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12659_
timestamp 0
transform -1 0 11370 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12660_
timestamp 0
transform -1 0 12490 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12661_
timestamp 0
transform 1 0 12110 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__12662_
timestamp 0
transform -1 0 12350 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__12663_
timestamp 0
transform -1 0 11970 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__12664_
timestamp 0
transform -1 0 12070 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__12665_
timestamp 0
transform 1 0 11930 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__12666_
timestamp 0
transform -1 0 11810 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__12667_
timestamp 0
transform -1 0 11990 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12668_
timestamp 0
transform -1 0 13310 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__12669_
timestamp 0
transform -1 0 16990 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12670_
timestamp 0
transform 1 0 16010 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__12671_
timestamp 0
transform 1 0 16670 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12672_
timestamp 0
transform -1 0 16530 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12673_
timestamp 0
transform -1 0 16650 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12674_
timestamp 0
transform 1 0 16850 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12675_
timestamp 0
transform 1 0 17050 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__12676_
timestamp 0
transform 1 0 16890 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__12677_
timestamp 0
transform -1 0 16570 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__12678_
timestamp 0
transform 1 0 16410 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__12679_
timestamp 0
transform -1 0 16150 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__12680_
timestamp 0
transform -1 0 16290 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__12681_
timestamp 0
transform 1 0 15910 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__12682_
timestamp 0
transform 1 0 16670 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__12683_
timestamp 0
transform 1 0 16510 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__12684_
timestamp 0
transform 1 0 16330 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__12685_
timestamp 0
transform -1 0 16230 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__12686_
timestamp 0
transform -1 0 13090 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12687_
timestamp 0
transform -1 0 13230 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12688_
timestamp 0
transform -1 0 12630 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12689_
timestamp 0
transform -1 0 14890 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__12690_
timestamp 0
transform -1 0 12750 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__12691_
timestamp 0
transform 1 0 12870 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__12692_
timestamp 0
transform -1 0 12490 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12693_
timestamp 0
transform 1 0 12030 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12694_
timestamp 0
transform -1 0 11550 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12695_
timestamp 0
transform 1 0 11330 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__12696_
timestamp 0
transform -1 0 12850 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12697_
timestamp 0
transform -1 0 16030 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12698_
timestamp 0
transform -1 0 16390 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__12699_
timestamp 0
transform -1 0 15870 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12700_
timestamp 0
transform 1 0 16150 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__12701_
timestamp 0
transform 1 0 16010 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__12702_
timestamp 0
transform -1 0 15870 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__12703_
timestamp 0
transform -1 0 15770 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__12704_
timestamp 0
transform -1 0 16510 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__12705_
timestamp 0
transform -1 0 16190 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__12706_
timestamp 0
transform -1 0 15610 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__12707_
timestamp 0
transform 1 0 14450 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__12708_
timestamp 0
transform 1 0 14430 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12709_
timestamp 0
transform 1 0 16350 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12710_
timestamp 0
transform 1 0 15730 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12711_
timestamp 0
transform 1 0 15870 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12712_
timestamp 0
transform -1 0 16650 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__12713_
timestamp 0
transform 1 0 16790 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12714_
timestamp 0
transform 1 0 16630 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12715_
timestamp 0
transform 1 0 16290 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12716_
timestamp 0
transform 1 0 17010 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__12717_
timestamp 0
transform 1 0 17050 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12718_
timestamp 0
transform 1 0 16910 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12719_
timestamp 0
transform 1 0 16670 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__12720_
timestamp 0
transform 1 0 16770 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__12721_
timestamp 0
transform 1 0 16970 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__12722_
timestamp 0
transform 1 0 16910 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12723_
timestamp 0
transform 1 0 16510 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12724_
timestamp 0
transform -1 0 14410 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12725_
timestamp 0
transform -1 0 15750 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12726_
timestamp 0
transform -1 0 16950 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12727_
timestamp 0
transform 1 0 16350 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12728_
timestamp 0
transform -1 0 16470 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__12729_
timestamp 0
transform 1 0 16710 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__12730_
timestamp 0
transform -1 0 16790 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12731_
timestamp 0
transform -1 0 16190 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12732_
timestamp 0
transform 1 0 14090 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__12733_
timestamp 0
transform -1 0 13890 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12734_
timestamp 0
transform -1 0 13790 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12735_
timestamp 0
transform -1 0 14050 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12736_
timestamp 0
transform -1 0 13630 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12737_
timestamp 0
transform -1 0 13550 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__12738_
timestamp 0
transform -1 0 13010 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12739_
timestamp 0
transform -1 0 12750 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12740_
timestamp 0
transform -1 0 11490 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__12741_
timestamp 0
transform -1 0 8990 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12742_
timestamp 0
transform 1 0 9210 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__12743_
timestamp 0
transform 1 0 9090 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__12744_
timestamp 0
transform -1 0 11710 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12745_
timestamp 0
transform -1 0 13350 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12746_
timestamp 0
transform 1 0 15530 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12747_
timestamp 0
transform -1 0 15710 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12748_
timestamp 0
transform -1 0 15670 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__12749_
timestamp 0
transform -1 0 15370 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__12750_
timestamp 0
transform 1 0 15470 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__12751_
timestamp 0
transform 1 0 15210 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__12752_
timestamp 0
transform -1 0 13810 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__12753_
timestamp 0
transform 1 0 13670 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__12754_
timestamp 0
transform 1 0 14170 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12755_
timestamp 0
transform -1 0 14570 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12756_
timestamp 0
transform 1 0 14270 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__12757_
timestamp 0
transform -1 0 13430 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12758_
timestamp 0
transform -1 0 13590 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12759_
timestamp 0
transform -1 0 13190 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12760_
timestamp 0
transform -1 0 12890 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12761_
timestamp 0
transform -1 0 12890 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12762_
timestamp 0
transform -1 0 12370 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12763_
timestamp 0
transform 1 0 13030 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12764_
timestamp 0
transform -1 0 12210 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12765_
timestamp 0
transform 1 0 12470 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12766_
timestamp 0
transform -1 0 12230 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12767_
timestamp 0
transform -1 0 12070 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12768_
timestamp 0
transform 1 0 11790 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12769_
timestamp 0
transform 1 0 12350 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12770_
timestamp 0
transform 1 0 13270 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12771_
timestamp 0
transform -1 0 12750 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12772_
timestamp 0
transform 1 0 14950 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12773_
timestamp 0
transform -1 0 13970 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__12774_
timestamp 0
transform 1 0 15130 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12775_
timestamp 0
transform -1 0 15330 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12776_
timestamp 0
transform 1 0 15430 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12777_
timestamp 0
transform 1 0 15610 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12778_
timestamp 0
transform 1 0 15470 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12779_
timestamp 0
transform 1 0 16990 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12780_
timestamp 0
transform 1 0 16790 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12781_
timestamp 0
transform 1 0 16450 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12782_
timestamp 0
transform 1 0 15210 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12783_
timestamp 0
transform -1 0 13170 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12784_
timestamp 0
transform -1 0 12970 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12785_
timestamp 0
transform -1 0 13230 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12786_
timestamp 0
transform 1 0 13050 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12787_
timestamp 0
transform -1 0 13210 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12788_
timestamp 0
transform 1 0 13330 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12789_
timestamp 0
transform -1 0 12970 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12790_
timestamp 0
transform -1 0 12850 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12791_
timestamp 0
transform -1 0 12590 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12792_
timestamp 0
transform -1 0 12450 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12793_
timestamp 0
transform 1 0 11890 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12794_
timestamp 0
transform -1 0 13070 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12795_
timestamp 0
transform -1 0 14050 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12796_
timestamp 0
transform 1 0 14950 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12797_
timestamp 0
transform 1 0 15370 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12798_
timestamp 0
transform 1 0 15210 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12799_
timestamp 0
transform -1 0 15370 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12800_
timestamp 0
transform -1 0 15370 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12801_
timestamp 0
transform 1 0 15570 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12802_
timestamp 0
transform -1 0 15090 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12803_
timestamp 0
transform -1 0 13470 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12804_
timestamp 0
transform -1 0 13630 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12805_
timestamp 0
transform -1 0 13470 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12806_
timestamp 0
transform 1 0 13910 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12807_
timestamp 0
transform 1 0 12770 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__12808_
timestamp 0
transform 1 0 13370 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12809_
timestamp 0
transform 1 0 13490 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12810_
timestamp 0
transform 1 0 13610 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12811_
timestamp 0
transform 1 0 13770 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12812_
timestamp 0
transform 1 0 12710 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12813_
timestamp 0
transform -1 0 12850 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12814_
timestamp 0
transform 1 0 12670 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12815_
timestamp 0
transform 1 0 11950 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12816_
timestamp 0
transform -1 0 12590 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12817_
timestamp 0
transform -1 0 14530 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__12818_
timestamp 0
transform 1 0 13310 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12819_
timestamp 0
transform 1 0 15630 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12820_
timestamp 0
transform 1 0 15790 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12821_
timestamp 0
transform 1 0 15650 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12822_
timestamp 0
transform 1 0 16370 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12823_
timestamp 0
transform -1 0 15510 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12824_
timestamp 0
transform -1 0 13770 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12825_
timestamp 0
transform 1 0 13570 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__12826_
timestamp 0
transform -1 0 14070 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12827_
timestamp 0
transform -1 0 13550 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__12828_
timestamp 0
transform -1 0 13250 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__12829_
timestamp 0
transform -1 0 13090 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__12830_
timestamp 0
transform -1 0 13290 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12831_
timestamp 0
transform 1 0 13090 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12832_
timestamp 0
transform -1 0 12550 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12833_
timestamp 0
transform -1 0 12410 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12834_
timestamp 0
transform -1 0 12250 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12835_
timestamp 0
transform 1 0 11470 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12836_
timestamp 0
transform 1 0 12130 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12837_
timestamp 0
transform -1 0 13530 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12838_
timestamp 0
transform 1 0 13370 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__12839_
timestamp 0
transform -1 0 15530 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12840_
timestamp 0
transform 1 0 15310 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12841_
timestamp 0
transform -1 0 15310 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__12842_
timestamp 0
transform -1 0 13470 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12843_
timestamp 0
transform -1 0 14090 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12844_
timestamp 0
transform 1 0 13910 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12845_
timestamp 0
transform 1 0 13790 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12846_
timestamp 0
transform -1 0 13250 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12847_
timestamp 0
transform -1 0 13670 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12848_
timestamp 0
transform 1 0 13930 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12849_
timestamp 0
transform -1 0 13530 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12850_
timestamp 0
transform -1 0 12730 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12851_
timestamp 0
transform -1 0 12950 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__12852_
timestamp 0
transform 1 0 12990 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12853_
timestamp 0
transform 1 0 12850 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12854_
timestamp 0
transform -1 0 12990 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12855_
timestamp 0
transform -1 0 12410 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12856_
timestamp 0
transform -1 0 12450 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12857_
timestamp 0
transform 1 0 12250 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12858_
timestamp 0
transform 1 0 11850 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12859_
timestamp 0
transform 1 0 13370 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12860_
timestamp 0
transform -1 0 13310 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12861_
timestamp 0
transform -1 0 13170 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12862_
timestamp 0
transform 1 0 13110 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12863_
timestamp 0
transform 1 0 13010 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12864_
timestamp 0
transform -1 0 13110 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12865_
timestamp 0
transform -1 0 13910 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12866_
timestamp 0
transform 1 0 13670 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__12867_
timestamp 0
transform 1 0 15190 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12868_
timestamp 0
transform -1 0 15330 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12869_
timestamp 0
transform -1 0 15230 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12870_
timestamp 0
transform 1 0 14690 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12871_
timestamp 0
transform -1 0 13770 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12872_
timestamp 0
transform -1 0 14310 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12873_
timestamp 0
transform 1 0 13590 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12874_
timestamp 0
transform 1 0 13730 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12875_
timestamp 0
transform -1 0 13630 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12876_
timestamp 0
transform 1 0 14010 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12877_
timestamp 0
transform 1 0 14170 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12878_
timestamp 0
transform -1 0 13890 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12879_
timestamp 0
transform -1 0 12990 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12880_
timestamp 0
transform -1 0 12870 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12881_
timestamp 0
transform 1 0 12950 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12882_
timestamp 0
transform 1 0 12570 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12883_
timestamp 0
transform -1 0 12270 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12884_
timestamp 0
transform -1 0 12050 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12885_
timestamp 0
transform -1 0 11950 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12886_
timestamp 0
transform -1 0 12110 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12887_
timestamp 0
transform 1 0 11950 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12888_
timestamp 0
transform -1 0 11410 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12889_
timestamp 0
transform 1 0 12830 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12890_
timestamp 0
transform -1 0 12570 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12891_
timestamp 0
transform -1 0 12690 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12892_
timestamp 0
transform 1 0 13550 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12893_
timestamp 0
transform -1 0 13830 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12894_
timestamp 0
transform 1 0 14650 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12895_
timestamp 0
transform -1 0 13670 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12896_
timestamp 0
transform 1 0 13970 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12897_
timestamp 0
transform 1 0 14130 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12898_
timestamp 0
transform 1 0 13970 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12899_
timestamp 0
transform -1 0 13430 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12900_
timestamp 0
transform -1 0 13830 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12901_
timestamp 0
transform -1 0 13690 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12902_
timestamp 0
transform -1 0 13550 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12903_
timestamp 0
transform -1 0 13350 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12904_
timestamp 0
transform -1 0 12510 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12905_
timestamp 0
transform -1 0 12350 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12906_
timestamp 0
transform -1 0 12210 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12907_
timestamp 0
transform 1 0 11750 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12908_
timestamp 0
transform 1 0 13550 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12909_
timestamp 0
transform -1 0 13430 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12910_
timestamp 0
transform 1 0 13250 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12911_
timestamp 0
transform -1 0 13290 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12912_
timestamp 0
transform 1 0 13110 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12913_
timestamp 0
transform -1 0 13330 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12914_
timestamp 0
transform 1 0 13190 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12915_
timestamp 0
transform 1 0 14230 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12916_
timestamp 0
transform 1 0 13990 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12917_
timestamp 0
transform 1 0 14650 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12918_
timestamp 0
transform 1 0 14930 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12919_
timestamp 0
transform -1 0 14510 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12920_
timestamp 0
transform 1 0 14770 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12921_
timestamp 0
transform 1 0 14530 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12922_
timestamp 0
transform 1 0 14370 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12923_
timestamp 0
transform 1 0 14350 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12924_
timestamp 0
transform 1 0 14490 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12925_
timestamp 0
transform -1 0 14110 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__12926_
timestamp 0
transform -1 0 13510 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12927_
timestamp 0
transform -1 0 12070 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12928_
timestamp 0
transform -1 0 12210 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12929_
timestamp 0
transform -1 0 11910 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12930_
timestamp 0
transform 1 0 11030 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__12931_
timestamp 0
transform 1 0 15050 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12932_
timestamp 0
transform -1 0 15190 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12933_
timestamp 0
transform -1 0 15090 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12934_
timestamp 0
transform 1 0 14910 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12935_
timestamp 0
transform 1 0 14770 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12936_
timestamp 0
transform -1 0 13970 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12937_
timestamp 0
transform 1 0 15170 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12938_
timestamp 0
transform -1 0 14510 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12939_
timestamp 0
transform 1 0 14370 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12940_
timestamp 0
transform 1 0 14670 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12941_
timestamp 0
transform -1 0 13810 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12942_
timestamp 0
transform -1 0 14110 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12943_
timestamp 0
transform -1 0 14230 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12944_
timestamp 0
transform -1 0 12890 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12945_
timestamp 0
transform -1 0 14250 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__12946_
timestamp 0
transform -1 0 13170 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12947_
timestamp 0
transform -1 0 13070 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12948_
timestamp 0
transform -1 0 12910 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12949_
timestamp 0
transform -1 0 12750 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12950_
timestamp 0
transform -1 0 13010 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12951_
timestamp 0
transform -1 0 12610 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12952_
timestamp 0
transform -1 0 12510 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12953_
timestamp 0
transform -1 0 12350 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12954_
timestamp 0
transform 1 0 11730 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12955_
timestamp 0
transform 1 0 11910 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__12956_
timestamp 0
transform -1 0 12810 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12957_
timestamp 0
transform 1 0 15070 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12958_
timestamp 0
transform 1 0 15430 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12959_
timestamp 0
transform -1 0 14850 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12960_
timestamp 0
transform -1 0 14810 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__12961_
timestamp 0
transform 1 0 13770 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12962_
timestamp 0
transform 1 0 13870 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12963_
timestamp 0
transform -1 0 13690 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__12964_
timestamp 0
transform -1 0 13670 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12965_
timestamp 0
transform 1 0 13150 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__12966_
timestamp 0
transform -1 0 12810 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__12967_
timestamp 0
transform 1 0 12630 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__12968_
timestamp 0
transform -1 0 13030 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__12969_
timestamp 0
transform -1 0 12650 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__12970_
timestamp 0
transform 1 0 12210 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__12971_
timestamp 0
transform -1 0 12890 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12972_
timestamp 0
transform 1 0 15690 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12973_
timestamp 0
transform -1 0 15830 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12974_
timestamp 0
transform -1 0 15950 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12975_
timestamp 0
transform 1 0 16250 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12976_
timestamp 0
transform 1 0 14030 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__12977_
timestamp 0
transform -1 0 14050 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__12978_
timestamp 0
transform 1 0 14150 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__12979_
timestamp 0
transform -1 0 16110 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12980_
timestamp 0
transform -1 0 14430 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12981_
timestamp 0
transform 1 0 14530 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12982_
timestamp 0
transform -1 0 14730 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12983_
timestamp 0
transform -1 0 14850 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12984_
timestamp 0
transform 1 0 16190 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12985_
timestamp 0
transform -1 0 16390 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12986_
timestamp 0
transform 1 0 16610 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__12987_
timestamp 0
transform -1 0 15790 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__12988_
timestamp 0
transform -1 0 15830 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12989_
timestamp 0
transform 1 0 16070 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12990_
timestamp 0
transform 1 0 15950 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__12991_
timestamp 0
transform 1 0 16010 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12992_
timestamp 0
transform -1 0 15770 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12993_
timestamp 0
transform -1 0 15610 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12994_
timestamp 0
transform 1 0 12330 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__12995_
timestamp 0
transform -1 0 15910 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__12996_
timestamp 0
transform -1 0 15090 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12997_
timestamp 0
transform -1 0 15230 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__12998_
timestamp 0
transform -1 0 15450 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__12999_
timestamp 0
transform 1 0 15170 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13000_
timestamp 0
transform -1 0 16450 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13001_
timestamp 0
transform 1 0 16570 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13002_
timestamp 0
transform 1 0 14370 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13003_
timestamp 0
transform 1 0 14210 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13004_
timestamp 0
transform 1 0 16010 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13005_
timestamp 0
transform -1 0 14190 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13006_
timestamp 0
transform -1 0 14330 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13007_
timestamp 0
transform 1 0 16410 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13008_
timestamp 0
transform 1 0 16270 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13009_
timestamp 0
transform 1 0 16430 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13010_
timestamp 0
transform -1 0 16970 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13011_
timestamp 0
transform 1 0 16110 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13012_
timestamp 0
transform -1 0 16690 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13013_
timestamp 0
transform 1 0 16490 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13014_
timestamp 0
transform -1 0 16170 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13015_
timestamp 0
transform 1 0 15890 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13016_
timestamp 0
transform -1 0 16310 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13017_
timestamp 0
transform -1 0 15750 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13018_
timestamp 0
transform 1 0 15610 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13019_
timestamp 0
transform -1 0 15470 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13020_
timestamp 0
transform 1 0 14370 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13021_
timestamp 0
transform -1 0 12470 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13022_
timestamp 0
transform -1 0 12250 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13023_
timestamp 0
transform 1 0 16010 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13024_
timestamp 0
transform 1 0 16610 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13025_
timestamp 0
transform 1 0 15010 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13026_
timestamp 0
transform 1 0 14870 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13027_
timestamp 0
transform 1 0 16090 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13028_
timestamp 0
transform 1 0 15950 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13029_
timestamp 0
transform -1 0 16170 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13030_
timestamp 0
transform 1 0 16310 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13031_
timestamp 0
transform -1 0 16190 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13032_
timestamp 0
transform -1 0 16170 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13033_
timestamp 0
transform 1 0 17050 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13034_
timestamp 0
transform -1 0 16770 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13035_
timestamp 0
transform 1 0 16770 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13036_
timestamp 0
transform 1 0 16910 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13037_
timestamp 0
transform 1 0 16730 0 1 250
box -6 -8 26 248
use FILL  FILL_0__13038_
timestamp 0
transform 1 0 16810 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13039_
timestamp 0
transform 1 0 16930 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13040_
timestamp 0
transform -1 0 16710 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13041_
timestamp 0
transform -1 0 16350 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13042_
timestamp 0
transform 1 0 15010 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13043_
timestamp 0
transform -1 0 16190 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13044_
timestamp 0
transform -1 0 12750 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13045_
timestamp 0
transform 1 0 16630 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13046_
timestamp 0
transform -1 0 16670 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13047_
timestamp 0
transform -1 0 15310 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13048_
timestamp 0
transform -1 0 15430 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13049_
timestamp 0
transform -1 0 15490 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13050_
timestamp 0
transform 1 0 16010 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13051_
timestamp 0
transform 1 0 16610 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13052_
timestamp 0
transform -1 0 16750 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13053_
timestamp 0
transform -1 0 16870 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13054_
timestamp 0
transform 1 0 16930 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13055_
timestamp 0
transform 1 0 16910 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13056_
timestamp 0
transform -1 0 16490 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13057_
timestamp 0
transform 1 0 16990 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__13058_
timestamp 0
transform 1 0 16990 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13059_
timestamp 0
transform 1 0 16910 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13060_
timestamp 0
transform -1 0 16850 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13061_
timestamp 0
transform 1 0 17010 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13062_
timestamp 0
transform -1 0 16570 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13063_
timestamp 0
transform 1 0 16710 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13064_
timestamp 0
transform 1 0 16430 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13065_
timestamp 0
transform 1 0 12590 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13066_
timestamp 0
transform 1 0 16770 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13067_
timestamp 0
transform -1 0 15350 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13068_
timestamp 0
transform 1 0 15250 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13069_
timestamp 0
transform -1 0 15690 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13070_
timestamp 0
transform -1 0 15830 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13071_
timestamp 0
transform 1 0 16370 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13072_
timestamp 0
transform 1 0 16490 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13073_
timestamp 0
transform 1 0 17030 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13074_
timestamp 0
transform 1 0 16490 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13075_
timestamp 0
transform -1 0 16890 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13076_
timestamp 0
transform -1 0 16910 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13077_
timestamp 0
transform -1 0 17030 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13078_
timestamp 0
transform -1 0 16770 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13079_
timestamp 0
transform -1 0 16610 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13080_
timestamp 0
transform -1 0 16890 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13081_
timestamp 0
transform -1 0 16730 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13082_
timestamp 0
transform -1 0 16690 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13083_
timestamp 0
transform -1 0 16570 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13084_
timestamp 0
transform 1 0 14430 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13085_
timestamp 0
transform -1 0 16290 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13086_
timestamp 0
transform -1 0 16150 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13087_
timestamp 0
transform 1 0 11790 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13088_
timestamp 0
transform -1 0 12250 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13089_
timestamp 0
transform 1 0 16390 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13090_
timestamp 0
transform 1 0 17010 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13091_
timestamp 0
transform -1 0 15550 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13092_
timestamp 0
transform -1 0 15410 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13093_
timestamp 0
transform 1 0 16290 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13094_
timestamp 0
transform 1 0 16230 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13095_
timestamp 0
transform -1 0 16470 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13096_
timestamp 0
transform 1 0 16970 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13097_
timestamp 0
transform -1 0 16830 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13098_
timestamp 0
transform 1 0 16650 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13099_
timestamp 0
transform 1 0 16730 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13100_
timestamp 0
transform 1 0 16590 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13101_
timestamp 0
transform -1 0 16570 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13102_
timestamp 0
transform -1 0 16050 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13103_
timestamp 0
transform 1 0 16690 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13104_
timestamp 0
transform 1 0 15910 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13105_
timestamp 0
transform 1 0 15770 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13106_
timestamp 0
transform -1 0 15650 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13107_
timestamp 0
transform -1 0 15510 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13108_
timestamp 0
transform 1 0 12570 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13109_
timestamp 0
transform 1 0 9510 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13110_
timestamp 0
transform 1 0 16550 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13111_
timestamp 0
transform 1 0 15530 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13112_
timestamp 0
transform -1 0 16090 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13113_
timestamp 0
transform 1 0 16210 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13114_
timestamp 0
transform -1 0 16230 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13115_
timestamp 0
transform -1 0 16370 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13116_
timestamp 0
transform 1 0 16350 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13117_
timestamp 0
transform 1 0 16190 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13118_
timestamp 0
transform -1 0 15970 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13119_
timestamp 0
transform 1 0 15930 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13120_
timestamp 0
transform -1 0 16090 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13121_
timestamp 0
transform 1 0 13610 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13122_
timestamp 0
transform 1 0 16810 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13123_
timestamp 0
transform 1 0 14890 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13124_
timestamp 0
transform -1 0 14290 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13125_
timestamp 0
transform -1 0 14010 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13126_
timestamp 0
transform 1 0 13730 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13127_
timestamp 0
transform -1 0 13050 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13128_
timestamp 0
transform -1 0 16430 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13129_
timestamp 0
transform -1 0 14610 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13130_
timestamp 0
transform -1 0 14770 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13131_
timestamp 0
transform -1 0 14130 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13132_
timestamp 0
transform -1 0 12930 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13133_
timestamp 0
transform -1 0 12110 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13134_
timestamp 0
transform 1 0 9750 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13135_
timestamp 0
transform 1 0 9610 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13136_
timestamp 0
transform 1 0 11270 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13137_
timestamp 0
transform -1 0 12410 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13138_
timestamp 0
transform 1 0 15950 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13139_
timestamp 0
transform -1 0 15690 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13140_
timestamp 0
transform 1 0 15630 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13141_
timestamp 0
transform 1 0 15510 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13142_
timestamp 0
transform -1 0 15610 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13143_
timestamp 0
transform 1 0 16070 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13144_
timestamp 0
transform -1 0 16290 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13145_
timestamp 0
transform 1 0 16150 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13146_
timestamp 0
transform -1 0 15350 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13147_
timestamp 0
transform -1 0 15750 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13148_
timestamp 0
transform -1 0 16030 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13149_
timestamp 0
transform 1 0 15870 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13150_
timestamp 0
transform 1 0 13850 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13151_
timestamp 0
transform -1 0 11850 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13152_
timestamp 0
transform 1 0 11970 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13153_
timestamp 0
transform -1 0 11730 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13154_
timestamp 0
transform -1 0 11590 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13155_
timestamp 0
transform 1 0 11390 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13156_
timestamp 0
transform 1 0 13350 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13157_
timestamp 0
transform -1 0 13510 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13158_
timestamp 0
transform -1 0 13210 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13159_
timestamp 0
transform -1 0 15090 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13160_
timestamp 0
transform -1 0 15810 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13161_
timestamp 0
transform -1 0 15850 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13162_
timestamp 0
transform -1 0 15690 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13163_
timestamp 0
transform -1 0 15090 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13164_
timestamp 0
transform 1 0 15170 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13165_
timestamp 0
transform -1 0 15450 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13166_
timestamp 0
transform 1 0 15310 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13167_
timestamp 0
transform -1 0 15190 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13168_
timestamp 0
transform -1 0 14950 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13169_
timestamp 0
transform -1 0 14970 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13170_
timestamp 0
transform -1 0 14810 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13171_
timestamp 0
transform -1 0 12510 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13172_
timestamp 0
transform -1 0 10930 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13173_
timestamp 0
transform 1 0 12630 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13174_
timestamp 0
transform -1 0 12250 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13175_
timestamp 0
transform 1 0 10750 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13176_
timestamp 0
transform -1 0 13290 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13177_
timestamp 0
transform 1 0 12770 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13178_
timestamp 0
transform -1 0 13830 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13179_
timestamp 0
transform -1 0 15230 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13180_
timestamp 0
transform 1 0 15410 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13181_
timestamp 0
transform 1 0 15630 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13182_
timestamp 0
transform 1 0 15510 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13183_
timestamp 0
transform -1 0 15290 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13184_
timestamp 0
transform -1 0 15010 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13185_
timestamp 0
transform 1 0 15150 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13186_
timestamp 0
transform 1 0 14790 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13187_
timestamp 0
transform -1 0 14450 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13188_
timestamp 0
transform -1 0 13790 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13189_
timestamp 0
transform 1 0 13910 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13190_
timestamp 0
transform -1 0 13650 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13191_
timestamp 0
transform -1 0 10150 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13192_
timestamp 0
transform -1 0 14570 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13193_
timestamp 0
transform -1 0 14530 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13194_
timestamp 0
transform 1 0 14670 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13195_
timestamp 0
transform -1 0 14670 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13196_
timestamp 0
transform 1 0 14350 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13197_
timestamp 0
transform -1 0 15710 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13198_
timestamp 0
transform -1 0 15590 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13199_
timestamp 0
transform -1 0 15390 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13200_
timestamp 0
transform -1 0 15090 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13201_
timestamp 0
transform 1 0 14850 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13202_
timestamp 0
transform -1 0 14730 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13203_
timestamp 0
transform -1 0 14570 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13204_
timestamp 0
transform -1 0 14810 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13205_
timestamp 0
transform 1 0 14930 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13206_
timestamp 0
transform -1 0 14670 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13207_
timestamp 0
transform 1 0 14310 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13208_
timestamp 0
transform -1 0 14090 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13209_
timestamp 0
transform 1 0 14230 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13210_
timestamp 0
transform -1 0 13950 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13211_
timestamp 0
transform 1 0 10250 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13212_
timestamp 0
transform -1 0 13010 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13213_
timestamp 0
transform -1 0 14230 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13214_
timestamp 0
transform -1 0 14090 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13215_
timestamp 0
transform -1 0 14430 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13216_
timestamp 0
transform 1 0 14290 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13217_
timestamp 0
transform -1 0 14150 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13218_
timestamp 0
transform -1 0 14030 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13219_
timestamp 0
transform -1 0 13690 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13220_
timestamp 0
transform -1 0 13530 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13221_
timestamp 0
transform -1 0 13390 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13222_
timestamp 0
transform -1 0 13330 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13223_
timestamp 0
transform -1 0 13250 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13224_
timestamp 0
transform -1 0 12730 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13225_
timestamp 0
transform 1 0 11570 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13226_
timestamp 0
transform -1 0 13210 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13227_
timestamp 0
transform -1 0 13050 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13228_
timestamp 0
transform 1 0 13310 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13229_
timestamp 0
transform -1 0 13630 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13230_
timestamp 0
transform -1 0 13190 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13231_
timestamp 0
transform -1 0 12890 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13232_
timestamp 0
transform -1 0 11610 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13233_
timestamp 0
transform 1 0 11170 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13234_
timestamp 0
transform -1 0 11450 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13235_
timestamp 0
transform -1 0 11330 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13236_
timestamp 0
transform -1 0 11390 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13237_
timestamp 0
transform -1 0 11270 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13238_
timestamp 0
transform -1 0 11150 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13239_
timestamp 0
transform 1 0 11510 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13240_
timestamp 0
transform -1 0 10970 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13241_
timestamp 0
transform 1 0 10930 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13242_
timestamp 0
transform -1 0 13770 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13243_
timestamp 0
transform 1 0 11730 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13244_
timestamp 0
transform -1 0 11910 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13245_
timestamp 0
transform -1 0 11270 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13246_
timestamp 0
transform -1 0 11110 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13247_
timestamp 0
transform 1 0 10510 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13248_
timestamp 0
transform -1 0 10410 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13249_
timestamp 0
transform -1 0 10290 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13250_
timestamp 0
transform 1 0 11210 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13251_
timestamp 0
transform -1 0 10150 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13252_
timestamp 0
transform -1 0 10050 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13253_
timestamp 0
transform -1 0 12070 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13254_
timestamp 0
transform 1 0 14470 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13255_
timestamp 0
transform -1 0 14330 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13256_
timestamp 0
transform 1 0 13390 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13257_
timestamp 0
transform 1 0 13470 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13258_
timestamp 0
transform -1 0 11150 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13259_
timestamp 0
transform 1 0 11270 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13260_
timestamp 0
transform -1 0 10870 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13261_
timestamp 0
transform -1 0 10750 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13262_
timestamp 0
transform -1 0 10570 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13263_
timestamp 0
transform 1 0 10630 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13264_
timestamp 0
transform -1 0 11030 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13265_
timestamp 0
transform -1 0 12010 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13266_
timestamp 0
transform 1 0 13830 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13267_
timestamp 0
transform -1 0 13990 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13268_
timestamp 0
transform 1 0 13690 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13269_
timestamp 0
transform -1 0 11870 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13270_
timestamp 0
transform 1 0 12010 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13271_
timestamp 0
transform -1 0 11770 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13272_
timestamp 0
transform 1 0 10970 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13273_
timestamp 0
transform -1 0 11230 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13274_
timestamp 0
transform 1 0 13410 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13275_
timestamp 0
transform -1 0 13910 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13276_
timestamp 0
transform 1 0 13890 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13277_
timestamp 0
transform -1 0 13750 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13278_
timestamp 0
transform -1 0 13630 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13279_
timestamp 0
transform -1 0 12370 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13280_
timestamp 0
transform 1 0 12510 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13281_
timestamp 0
transform 1 0 11730 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13282_
timestamp 0
transform -1 0 11470 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13283_
timestamp 0
transform 1 0 11090 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13284_
timestamp 0
transform -1 0 10710 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13285_
timestamp 0
transform 1 0 10570 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13286_
timestamp 0
transform 1 0 10910 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13287_
timestamp 0
transform -1 0 11370 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13288_
timestamp 0
transform 1 0 10830 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13289_
timestamp 0
transform 1 0 11570 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13290_
timestamp 0
transform -1 0 11130 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13291_
timestamp 0
transform 1 0 10950 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13292_
timestamp 0
transform -1 0 14610 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13293_
timestamp 0
transform 1 0 14390 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13294_
timestamp 0
transform 1 0 14270 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13295_
timestamp 0
transform -1 0 14190 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13296_
timestamp 0
transform -1 0 14150 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13297_
timestamp 0
transform 1 0 12410 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13298_
timestamp 0
transform -1 0 12270 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13299_
timestamp 0
transform 1 0 12150 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13300_
timestamp 0
transform -1 0 11370 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13301_
timestamp 0
transform -1 0 11230 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13302_
timestamp 0
transform -1 0 11430 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13303_
timestamp 0
transform -1 0 12130 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13304_
timestamp 0
transform 1 0 12530 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13305_
timestamp 0
transform -1 0 13190 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13306_
timestamp 0
transform -1 0 13050 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13307_
timestamp 0
transform -1 0 12930 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13308_
timestamp 0
transform 1 0 12770 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13309_
timestamp 0
transform 1 0 12810 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13310_
timestamp 0
transform 1 0 12630 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13311_
timestamp 0
transform 1 0 12690 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13312_
timestamp 0
transform 1 0 11970 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13313_
timestamp 0
transform -1 0 11830 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13314_
timestamp 0
transform 1 0 11650 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13315_
timestamp 0
transform 1 0 13050 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13316_
timestamp 0
transform -1 0 12750 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13317_
timestamp 0
transform -1 0 12590 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13318_
timestamp 0
transform 1 0 12190 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13319_
timestamp 0
transform -1 0 12450 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13320_
timestamp 0
transform -1 0 12310 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13321_
timestamp 0
transform 1 0 12270 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13322_
timestamp 0
transform 1 0 11870 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13323_
timestamp 0
transform 1 0 11610 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13324_
timestamp 0
transform 1 0 11450 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13325_
timestamp 0
transform 1 0 11510 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13326_
timestamp 0
transform 1 0 11670 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13327_
timestamp 0
transform -1 0 12070 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13328_
timestamp 0
transform 1 0 12210 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13329_
timestamp 0
transform 1 0 11910 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13330_
timestamp 0
transform -1 0 11710 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13331_
timestamp 0
transform 1 0 11770 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13332_
timestamp 0
transform 1 0 11590 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13333_
timestamp 0
transform 1 0 11830 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13334_
timestamp 0
transform 1 0 11970 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13335_
timestamp 0
transform -1 0 11990 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13336_
timestamp 0
transform 1 0 11810 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13337_
timestamp 0
transform 1 0 12950 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13338_
timestamp 0
transform -1 0 12850 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13339_
timestamp 0
transform 1 0 12930 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13340_
timestamp 0
transform -1 0 12830 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13341_
timestamp 0
transform -1 0 11610 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13342_
timestamp 0
transform -1 0 12150 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13343_
timestamp 0
transform -1 0 11770 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13344_
timestamp 0
transform 1 0 11930 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13345_
timestamp 0
transform 1 0 12190 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13346_
timestamp 0
transform 1 0 12050 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13347_
timestamp 0
transform -1 0 14690 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13348_
timestamp 0
transform 1 0 14910 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13349_
timestamp 0
transform -1 0 15070 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13350_
timestamp 0
transform -1 0 15170 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13351_
timestamp 0
transform 1 0 14990 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13352_
timestamp 0
transform 1 0 14710 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13353_
timestamp 0
transform 1 0 14850 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13354_
timestamp 0
transform -1 0 14970 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13355_
timestamp 0
transform -1 0 15110 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13356_
timestamp 0
transform 1 0 15010 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13357_
timestamp 0
transform 1 0 15150 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13358_
timestamp 0
transform -1 0 11630 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13359_
timestamp 0
transform -1 0 15290 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13360_
timestamp 0
transform 1 0 15110 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13361_
timestamp 0
transform -1 0 15250 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13362_
timestamp 0
transform 1 0 15090 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13363_
timestamp 0
transform 1 0 12310 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13364_
timestamp 0
transform 1 0 16550 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13365_
timestamp 0
transform -1 0 16810 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13366_
timestamp 0
transform 1 0 16790 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13367_
timestamp 0
transform 1 0 16750 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13368_
timestamp 0
transform 1 0 15230 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13369_
timestamp 0
transform 1 0 15090 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13370_
timestamp 0
transform 1 0 14790 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13371_
timestamp 0
transform -1 0 14970 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13372_
timestamp 0
transform -1 0 15650 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13373_
timestamp 0
transform -1 0 15790 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13374_
timestamp 0
transform -1 0 16050 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13375_
timestamp 0
transform 1 0 16170 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13376_
timestamp 0
transform 1 0 14090 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13377_
timestamp 0
transform -1 0 14230 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13378_
timestamp 0
transform -1 0 14650 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13379_
timestamp 0
transform -1 0 14770 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13380_
timestamp 0
transform 1 0 14030 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13381_
timestamp 0
transform 1 0 14910 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13382_
timestamp 0
transform 1 0 14750 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13383_
timestamp 0
transform 1 0 14230 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13384_
timestamp 0
transform 1 0 14290 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13385_
timestamp 0
transform 1 0 14370 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13386_
timestamp 0
transform -1 0 13810 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13387_
timestamp 0
transform -1 0 13850 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13388_
timestamp 0
transform -1 0 13950 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13389_
timestamp 0
transform -1 0 14230 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13390_
timestamp 0
transform 1 0 14150 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13391_
timestamp 0
transform 1 0 14270 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13392_
timestamp 0
transform -1 0 14610 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13393_
timestamp 0
transform 1 0 14450 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13394_
timestamp 0
transform -1 0 13510 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13395_
timestamp 0
transform -1 0 13670 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13396_
timestamp 0
transform 1 0 14510 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13397_
timestamp 0
transform 1 0 14330 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13398_
timestamp 0
transform 1 0 12970 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13399_
timestamp 0
transform -1 0 13130 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13400_
timestamp 0
transform -1 0 14830 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13401_
timestamp 0
transform -1 0 14950 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13402_
timestamp 0
transform -1 0 11930 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13403_
timestamp 0
transform -1 0 12050 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13404_
timestamp 0
transform 1 0 12950 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13405_
timestamp 0
transform -1 0 13090 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13406_
timestamp 0
transform -1 0 11930 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13407_
timestamp 0
transform -1 0 12690 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13408_
timestamp 0
transform 1 0 12510 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13409_
timestamp 0
transform -1 0 12550 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13410_
timestamp 0
transform -1 0 12730 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13411_
timestamp 0
transform 1 0 12570 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13412_
timestamp 0
transform -1 0 11650 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13413_
timestamp 0
transform -1 0 11770 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13414_
timestamp 0
transform 1 0 12410 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13415_
timestamp 0
transform -1 0 12270 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13416_
timestamp 0
transform 1 0 12570 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13417_
timestamp 0
transform 1 0 12410 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13418_
timestamp 0
transform 1 0 12910 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13419_
timestamp 0
transform -1 0 13050 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13420_
timestamp 0
transform -1 0 11630 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13421_
timestamp 0
transform -1 0 11790 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13422_
timestamp 0
transform -1 0 12190 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13423_
timestamp 0
transform -1 0 12350 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13424_
timestamp 0
transform -1 0 12450 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13425_
timestamp 0
transform -1 0 12570 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13426_
timestamp 0
transform 1 0 11050 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13427_
timestamp 0
transform -1 0 10790 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13502_
timestamp 0
transform -1 0 7630 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13503_
timestamp 0
transform -1 0 7490 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13504_
timestamp 0
transform -1 0 7770 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13505_
timestamp 0
transform 1 0 7930 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13506_
timestamp 0
transform 1 0 8330 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13507_
timestamp 0
transform 1 0 8570 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13508_
timestamp 0
transform 1 0 8410 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13509_
timestamp 0
transform -1 0 7730 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13510_
timestamp 0
transform -1 0 7130 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13511_
timestamp 0
transform 1 0 7170 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13512_
timestamp 0
transform -1 0 7050 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13513_
timestamp 0
transform 1 0 6350 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13514_
timestamp 0
transform 1 0 7390 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13515_
timestamp 0
transform -1 0 7650 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13516_
timestamp 0
transform 1 0 7790 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13517_
timestamp 0
transform -1 0 7130 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13518_
timestamp 0
transform 1 0 7910 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13519_
timestamp 0
transform 1 0 7530 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13520_
timestamp 0
transform 1 0 8050 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13521_
timestamp 0
transform -1 0 7810 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13522_
timestamp 0
transform 1 0 7790 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13523_
timestamp 0
transform 1 0 7510 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13524_
timestamp 0
transform -1 0 7670 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13525_
timestamp 0
transform -1 0 7650 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13526_
timestamp 0
transform -1 0 6970 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13527_
timestamp 0
transform 1 0 7550 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__13528_
timestamp 0
transform -1 0 10090 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13529_
timestamp 0
transform 1 0 9030 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13530_
timestamp 0
transform -1 0 8890 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13531_
timestamp 0
transform -1 0 9470 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13532_
timestamp 0
transform -1 0 8710 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13533_
timestamp 0
transform 1 0 8670 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13534_
timestamp 0
transform -1 0 8730 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13535_
timestamp 0
transform -1 0 7870 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13536_
timestamp 0
transform 1 0 8210 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13537_
timestamp 0
transform 1 0 8650 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13538_
timestamp 0
transform 1 0 8890 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13539_
timestamp 0
transform -1 0 9190 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13540_
timestamp 0
transform -1 0 8550 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13541_
timestamp 0
transform -1 0 8830 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__13542_
timestamp 0
transform 1 0 8250 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13543_
timestamp 0
transform -1 0 8290 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13544_
timestamp 0
transform -1 0 7130 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13545_
timestamp 0
transform 1 0 6690 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13546_
timestamp 0
transform -1 0 7870 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13547_
timestamp 0
transform -1 0 7550 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13548_
timestamp 0
transform 1 0 10230 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13549_
timestamp 0
transform -1 0 9870 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13550_
timestamp 0
transform -1 0 9990 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13551_
timestamp 0
transform 1 0 10190 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13552_
timestamp 0
transform -1 0 9730 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13553_
timestamp 0
transform -1 0 10010 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13554_
timestamp 0
transform 1 0 9830 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13555_
timestamp 0
transform -1 0 7750 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13556_
timestamp 0
transform -1 0 8150 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13557_
timestamp 0
transform 1 0 7830 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13558_
timestamp 0
transform 1 0 8110 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13559_
timestamp 0
transform -1 0 8450 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13560_
timestamp 0
transform 1 0 8270 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13561_
timestamp 0
transform 1 0 7970 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13562_
timestamp 0
transform -1 0 7590 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13563_
timestamp 0
transform 1 0 7090 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13564_
timestamp 0
transform -1 0 6590 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13565_
timestamp 0
transform 1 0 7270 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13566_
timestamp 0
transform -1 0 8850 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13567_
timestamp 0
transform 1 0 9370 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13568_
timestamp 0
transform 1 0 9890 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13569_
timestamp 0
transform 1 0 7390 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13570_
timestamp 0
transform 1 0 7230 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13571_
timestamp 0
transform -1 0 8170 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13572_
timestamp 0
transform -1 0 6190 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13573_
timestamp 0
transform 1 0 8430 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13574_
timestamp 0
transform -1 0 9250 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13575_
timestamp 0
transform -1 0 9430 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13576_
timestamp 0
transform -1 0 8570 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13577_
timestamp 0
transform -1 0 7410 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13578_
timestamp 0
transform -1 0 7710 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13579_
timestamp 0
transform 1 0 7810 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13580_
timestamp 0
transform 1 0 8110 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13581_
timestamp 0
transform -1 0 8450 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13582_
timestamp 0
transform 1 0 8270 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13583_
timestamp 0
transform 1 0 7950 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13584_
timestamp 0
transform -1 0 7050 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13585_
timestamp 0
transform 1 0 10310 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13586_
timestamp 0
transform -1 0 9650 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13587_
timestamp 0
transform -1 0 9370 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13588_
timestamp 0
transform -1 0 9510 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13589_
timestamp 0
transform -1 0 9610 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13590_
timestamp 0
transform -1 0 9310 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13591_
timestamp 0
transform 1 0 9230 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13592_
timestamp 0
transform -1 0 8950 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13593_
timestamp 0
transform -1 0 8350 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13594_
timestamp 0
transform 1 0 9290 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13595_
timestamp 0
transform 1 0 9150 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13596_
timestamp 0
transform 1 0 8870 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13597_
timestamp 0
transform 1 0 8590 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13598_
timestamp 0
transform -1 0 8330 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13599_
timestamp 0
transform 1 0 7710 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13600_
timestamp 0
transform -1 0 7130 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13601_
timestamp 0
transform 1 0 6270 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13602_
timestamp 0
transform 1 0 9190 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13603_
timestamp 0
transform -1 0 9290 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13604_
timestamp 0
transform 1 0 9030 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13605_
timestamp 0
transform 1 0 9130 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13606_
timestamp 0
transform 1 0 8790 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13607_
timestamp 0
transform -1 0 8990 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13608_
timestamp 0
transform -1 0 7410 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13609_
timestamp 0
transform 1 0 6790 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13610_
timestamp 0
transform -1 0 6390 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13611_
timestamp 0
transform -1 0 6130 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13612_
timestamp 0
transform 1 0 6510 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13613_
timestamp 0
transform 1 0 6210 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13614_
timestamp 0
transform -1 0 6570 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13615_
timestamp 0
transform 1 0 6270 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13616_
timestamp 0
transform -1 0 6450 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13617_
timestamp 0
transform -1 0 6330 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13618_
timestamp 0
transform 1 0 9090 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__13619_
timestamp 0
transform 1 0 9370 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__13620_
timestamp 0
transform 1 0 9210 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__13621_
timestamp 0
transform 1 0 6990 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13622_
timestamp 0
transform -1 0 6070 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13623_
timestamp 0
transform -1 0 9270 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13624_
timestamp 0
transform 1 0 9210 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13625_
timestamp 0
transform -1 0 8390 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13626_
timestamp 0
transform -1 0 8090 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13627_
timestamp 0
transform 1 0 8190 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13628_
timestamp 0
transform -1 0 7950 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13629_
timestamp 0
transform -1 0 6670 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13630_
timestamp 0
transform -1 0 5530 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13631_
timestamp 0
transform -1 0 6030 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13632_
timestamp 0
transform -1 0 6130 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13633_
timestamp 0
transform -1 0 5910 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13634_
timestamp 0
transform -1 0 5230 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13635_
timestamp 0
transform -1 0 5390 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13636_
timestamp 0
transform -1 0 4750 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13637_
timestamp 0
transform -1 0 4590 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13638_
timestamp 0
transform -1 0 5270 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13639_
timestamp 0
transform 1 0 5370 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13640_
timestamp 0
transform 1 0 4830 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13641_
timestamp 0
transform 1 0 5490 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13642_
timestamp 0
transform 1 0 6730 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13643_
timestamp 0
transform 1 0 6550 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13644_
timestamp 0
transform 1 0 6690 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13645_
timestamp 0
transform 1 0 6850 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13646_
timestamp 0
transform -1 0 6650 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13647_
timestamp 0
transform -1 0 5090 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13648_
timestamp 0
transform -1 0 4990 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13649_
timestamp 0
transform -1 0 5790 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13650_
timestamp 0
transform 1 0 6790 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13651_
timestamp 0
transform 1 0 9870 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13652_
timestamp 0
transform 1 0 10090 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13653_
timestamp 0
transform 1 0 9930 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13654_
timestamp 0
transform 1 0 8970 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13655_
timestamp 0
transform 1 0 8830 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13656_
timestamp 0
transform 1 0 7270 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13657_
timestamp 0
transform 1 0 6310 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13658_
timestamp 0
transform -1 0 7550 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13659_
timestamp 0
transform 1 0 7630 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13660_
timestamp 0
transform -1 0 5990 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13661_
timestamp 0
transform -1 0 5870 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13662_
timestamp 0
transform 1 0 6030 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13663_
timestamp 0
transform -1 0 5710 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13664_
timestamp 0
transform -1 0 5630 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13665_
timestamp 0
transform 1 0 5750 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13666_
timestamp 0
transform -1 0 4370 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13667_
timestamp 0
transform -1 0 4470 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13668_
timestamp 0
transform 1 0 4950 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13669_
timestamp 0
transform 1 0 5110 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13670_
timestamp 0
transform -1 0 5590 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13671_
timestamp 0
transform 1 0 5630 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13672_
timestamp 0
transform -1 0 5590 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13673_
timestamp 0
transform 1 0 10230 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13674_
timestamp 0
transform 1 0 9930 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13675_
timestamp 0
transform 1 0 9770 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13676_
timestamp 0
transform 1 0 9270 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13677_
timestamp 0
transform 1 0 9110 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13678_
timestamp 0
transform 1 0 7810 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13679_
timestamp 0
transform -1 0 7690 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13680_
timestamp 0
transform -1 0 7050 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13681_
timestamp 0
transform 1 0 6250 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13682_
timestamp 0
transform -1 0 5950 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13683_
timestamp 0
transform -1 0 6550 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13684_
timestamp 0
transform -1 0 6390 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13685_
timestamp 0
transform -1 0 6110 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13686_
timestamp 0
transform 1 0 6130 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13687_
timestamp 0
transform -1 0 5990 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13688_
timestamp 0
transform -1 0 5850 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13689_
timestamp 0
transform 1 0 6010 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13690_
timestamp 0
transform -1 0 6070 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13691_
timestamp 0
transform 1 0 5910 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13692_
timestamp 0
transform -1 0 5950 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13693_
timestamp 0
transform -1 0 6210 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13694_
timestamp 0
transform -1 0 6970 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13695_
timestamp 0
transform 1 0 6130 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13696_
timestamp 0
transform 1 0 9630 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13697_
timestamp 0
transform -1 0 9410 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13698_
timestamp 0
transform -1 0 8710 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13699_
timestamp 0
transform 1 0 7450 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13700_
timestamp 0
transform -1 0 7330 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13701_
timestamp 0
transform 1 0 6250 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13702_
timestamp 0
transform -1 0 6830 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13703_
timestamp 0
transform 1 0 6570 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13704_
timestamp 0
transform -1 0 6730 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13705_
timestamp 0
transform 1 0 6450 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13706_
timestamp 0
transform -1 0 6430 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13707_
timestamp 0
transform -1 0 5750 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13708_
timestamp 0
transform 1 0 6830 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13709_
timestamp 0
transform 1 0 6270 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13710_
timestamp 0
transform 1 0 6410 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13711_
timestamp 0
transform 1 0 6470 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13712_
timestamp 0
transform -1 0 7290 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__13713_
timestamp 0
transform -1 0 5770 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13714_
timestamp 0
transform 1 0 7650 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13715_
timestamp 0
transform 1 0 6650 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13716_
timestamp 0
transform -1 0 8990 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13717_
timestamp 0
transform 1 0 8310 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13718_
timestamp 0
transform 1 0 8150 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13719_
timestamp 0
transform -1 0 6650 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13720_
timestamp 0
transform 1 0 7390 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13721_
timestamp 0
transform -1 0 6130 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13722_
timestamp 0
transform -1 0 6610 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13723_
timestamp 0
transform -1 0 6350 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13724_
timestamp 0
transform -1 0 7130 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13725_
timestamp 0
transform 1 0 6990 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13726_
timestamp 0
transform -1 0 6990 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13727_
timestamp 0
transform -1 0 6190 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13728_
timestamp 0
transform 1 0 6230 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13729_
timestamp 0
transform -1 0 5850 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13730_
timestamp 0
transform 1 0 6550 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13731_
timestamp 0
transform -1 0 6730 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13732_
timestamp 0
transform -1 0 6030 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13733_
timestamp 0
transform -1 0 6050 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13734_
timestamp 0
transform 1 0 5870 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13735_
timestamp 0
transform -1 0 6830 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13736_
timestamp 0
transform -1 0 6510 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13737_
timestamp 0
transform 1 0 6150 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13738_
timestamp 0
transform 1 0 6310 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13739_
timestamp 0
transform -1 0 5970 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13740_
timestamp 0
transform 1 0 6410 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13741_
timestamp 0
transform 1 0 6430 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13742_
timestamp 0
transform -1 0 7330 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13743_
timestamp 0
transform 1 0 6850 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13744_
timestamp 0
transform -1 0 9670 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13745_
timestamp 0
transform 1 0 9630 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13746_
timestamp 0
transform -1 0 9530 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13747_
timestamp 0
transform 1 0 8690 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13748_
timestamp 0
transform 1 0 7250 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13749_
timestamp 0
transform -1 0 7070 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13750_
timestamp 0
transform 1 0 6770 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13751_
timestamp 0
transform -1 0 6930 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13752_
timestamp 0
transform -1 0 7190 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13753_
timestamp 0
transform 1 0 7150 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13754_
timestamp 0
transform -1 0 6890 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13755_
timestamp 0
transform -1 0 7030 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13756_
timestamp 0
transform -1 0 6730 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13757_
timestamp 0
transform 1 0 7010 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13758_
timestamp 0
transform -1 0 6890 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13759_
timestamp 0
transform 1 0 6430 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13760_
timestamp 0
transform 1 0 6570 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13761_
timestamp 0
transform -1 0 6870 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13762_
timestamp 0
transform -1 0 6870 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13763_
timestamp 0
transform 1 0 6710 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13764_
timestamp 0
transform -1 0 6690 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13765_
timestamp 0
transform -1 0 6930 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13766_
timestamp 0
transform 1 0 6590 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13767_
timestamp 0
transform 1 0 6310 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13768_
timestamp 0
transform 1 0 6430 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13769_
timestamp 0
transform -1 0 8090 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13770_
timestamp 0
transform 1 0 7870 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13771_
timestamp 0
transform 1 0 8550 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13772_
timestamp 0
transform -1 0 8350 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13773_
timestamp 0
transform -1 0 8050 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13774_
timestamp 0
transform 1 0 8310 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13775_
timestamp 0
transform -1 0 8030 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13776_
timestamp 0
transform -1 0 7950 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13777_
timestamp 0
transform -1 0 8190 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13778_
timestamp 0
transform 1 0 8170 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13779_
timestamp 0
transform -1 0 7770 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13780_
timestamp 0
transform 1 0 7490 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13781_
timestamp 0
transform -1 0 7270 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13782_
timestamp 0
transform -1 0 7110 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13783_
timestamp 0
transform -1 0 6970 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13784_
timestamp 0
transform -1 0 6870 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13785_
timestamp 0
transform 1 0 6750 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13786_
timestamp 0
transform -1 0 6630 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13787_
timestamp 0
transform 1 0 6270 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13788_
timestamp 0
transform -1 0 6590 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13789_
timestamp 0
transform 1 0 6450 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13790_
timestamp 0
transform -1 0 7670 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13791_
timestamp 0
transform -1 0 7370 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13792_
timestamp 0
transform -1 0 8950 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13793_
timestamp 0
transform 1 0 8170 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13794_
timestamp 0
transform -1 0 8530 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13795_
timestamp 0
transform 1 0 8550 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13796_
timestamp 0
transform -1 0 8370 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13797_
timestamp 0
transform 1 0 8610 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13798_
timestamp 0
transform 1 0 8470 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13799_
timestamp 0
transform -1 0 8070 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13800_
timestamp 0
transform 1 0 8630 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13801_
timestamp 0
transform -1 0 8730 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13802_
timestamp 0
transform -1 0 8810 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13803_
timestamp 0
transform -1 0 7790 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13804_
timestamp 0
transform -1 0 7290 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13805_
timestamp 0
transform 1 0 7430 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13806_
timestamp 0
transform -1 0 7290 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13807_
timestamp 0
transform -1 0 7410 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__13808_
timestamp 0
transform -1 0 9790 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13809_
timestamp 0
transform -1 0 8850 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13810_
timestamp 0
transform 1 0 8990 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13811_
timestamp 0
transform 1 0 9090 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13812_
timestamp 0
transform 1 0 9050 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13813_
timestamp 0
transform 1 0 9190 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13814_
timestamp 0
transform -1 0 8890 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13815_
timestamp 0
transform -1 0 8910 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13816_
timestamp 0
transform -1 0 8790 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13817_
timestamp 0
transform 1 0 9210 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13818_
timestamp 0
transform 1 0 9330 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13819_
timestamp 0
transform -1 0 9330 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13820_
timestamp 0
transform 1 0 9050 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13821_
timestamp 0
transform 1 0 8510 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13822_
timestamp 0
transform -1 0 8230 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13823_
timestamp 0
transform 1 0 7890 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13824_
timestamp 0
transform 1 0 7630 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13825_
timestamp 0
transform 1 0 8210 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13826_
timestamp 0
transform -1 0 8390 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13827_
timestamp 0
transform 1 0 7910 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13828_
timestamp 0
transform 1 0 8070 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13829_
timestamp 0
transform -1 0 8030 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13830_
timestamp 0
transform -1 0 7610 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13831_
timestamp 0
transform 1 0 7070 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13832_
timestamp 0
transform -1 0 7330 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13833_
timestamp 0
transform -1 0 8330 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13834_
timestamp 0
transform -1 0 10090 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13835_
timestamp 0
transform 1 0 10410 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13836_
timestamp 0
transform 1 0 10010 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13837_
timestamp 0
transform -1 0 9950 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__13838_
timestamp 0
transform 1 0 9750 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13839_
timestamp 0
transform -1 0 9450 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13840_
timestamp 0
transform -1 0 9450 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13841_
timestamp 0
transform 1 0 9310 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13842_
timestamp 0
transform -1 0 7990 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13843_
timestamp 0
transform -1 0 7770 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13844_
timestamp 0
transform 1 0 8150 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13845_
timestamp 0
transform -1 0 7890 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13846_
timestamp 0
transform -1 0 7450 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__13847_
timestamp 0
transform 1 0 7450 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13848_
timestamp 0
transform -1 0 8430 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__13849_
timestamp 0
transform -1 0 5790 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13850_
timestamp 0
transform -1 0 5670 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13851_
timestamp 0
transform -1 0 5910 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13852_
timestamp 0
transform -1 0 6070 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13853_
timestamp 0
transform -1 0 6710 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13854_
timestamp 0
transform 1 0 6970 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13855_
timestamp 0
transform 1 0 6810 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13856_
timestamp 0
transform -1 0 6710 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13857_
timestamp 0
transform -1 0 7770 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13858_
timestamp 0
transform -1 0 7890 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13859_
timestamp 0
transform 1 0 6690 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13860_
timestamp 0
transform 1 0 6650 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13861_
timestamp 0
transform -1 0 7910 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13862_
timestamp 0
transform 1 0 7950 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13863_
timestamp 0
transform 1 0 7790 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13864_
timestamp 0
transform -1 0 8010 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13865_
timestamp 0
transform -1 0 7410 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13866_
timestamp 0
transform 1 0 7890 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13867_
timestamp 0
transform 1 0 7510 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13868_
timestamp 0
transform 1 0 7630 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13869_
timestamp 0
transform 1 0 8570 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13870_
timestamp 0
transform 1 0 8630 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__13871_
timestamp 0
transform -1 0 8150 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13872_
timestamp 0
transform -1 0 8230 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13873_
timestamp 0
transform 1 0 5470 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13874_
timestamp 0
transform -1 0 5930 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13875_
timestamp 0
transform -1 0 6250 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13876_
timestamp 0
transform -1 0 6390 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13877_
timestamp 0
transform -1 0 6530 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13878_
timestamp 0
transform -1 0 7150 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13879_
timestamp 0
transform 1 0 7750 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13880_
timestamp 0
transform 1 0 7590 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13881_
timestamp 0
transform -1 0 7090 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13882_
timestamp 0
transform 1 0 7510 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13883_
timestamp 0
transform 1 0 7270 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13884_
timestamp 0
transform -1 0 6870 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13885_
timestamp 0
transform -1 0 6990 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13886_
timestamp 0
transform -1 0 7270 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13887_
timestamp 0
transform -1 0 8090 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13888_
timestamp 0
transform -1 0 7370 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13889_
timestamp 0
transform 1 0 7170 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13890_
timestamp 0
transform -1 0 8190 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13891_
timestamp 0
transform 1 0 8450 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13892_
timestamp 0
transform 1 0 8750 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13893_
timestamp 0
transform 1 0 8310 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13894_
timestamp 0
transform -1 0 8610 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13895_
timestamp 0
transform 1 0 8190 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13896_
timestamp 0
transform -1 0 8050 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13897_
timestamp 0
transform -1 0 7910 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13898_
timestamp 0
transform 1 0 7990 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13899_
timestamp 0
transform -1 0 7490 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13900_
timestamp 0
transform 1 0 8450 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13901_
timestamp 0
transform 1 0 8390 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13902_
timestamp 0
transform 1 0 9530 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13903_
timestamp 0
transform 1 0 9490 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13904_
timestamp 0
transform -1 0 8770 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13905_
timestamp 0
transform -1 0 9110 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13906_
timestamp 0
transform -1 0 6190 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13907_
timestamp 0
transform -1 0 6590 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13908_
timestamp 0
transform 1 0 6430 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13909_
timestamp 0
transform -1 0 7230 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13910_
timestamp 0
transform 1 0 8530 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13911_
timestamp 0
transform 1 0 8630 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13912_
timestamp 0
transform 1 0 8030 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13913_
timestamp 0
transform 1 0 8870 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13914_
timestamp 0
transform 1 0 9010 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13915_
timestamp 0
transform 1 0 8830 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13916_
timestamp 0
transform -1 0 8870 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13917_
timestamp 0
transform 1 0 8710 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13918_
timestamp 0
transform -1 0 8450 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13919_
timestamp 0
transform -1 0 8610 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13920_
timestamp 0
transform 1 0 8710 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13921_
timestamp 0
transform -1 0 7630 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__13922_
timestamp 0
transform 1 0 8710 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13923_
timestamp 0
transform -1 0 7110 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13924_
timestamp 0
transform -1 0 9510 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13925_
timestamp 0
transform -1 0 9630 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__13926_
timestamp 0
transform 1 0 10010 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13927_
timestamp 0
transform 1 0 9390 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13928_
timestamp 0
transform 1 0 7630 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13929_
timestamp 0
transform 1 0 7510 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13930_
timestamp 0
transform 1 0 7750 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13931_
timestamp 0
transform 1 0 9450 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13932_
timestamp 0
transform 1 0 8790 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13933_
timestamp 0
transform -1 0 8970 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13934_
timestamp 0
transform -1 0 9050 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13935_
timestamp 0
transform -1 0 7890 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13936_
timestamp 0
transform -1 0 7490 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13937_
timestamp 0
transform -1 0 7730 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13938_
timestamp 0
transform -1 0 7370 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13939_
timestamp 0
transform -1 0 6710 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13940_
timestamp 0
transform -1 0 6990 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13941_
timestamp 0
transform -1 0 6870 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13942_
timestamp 0
transform -1 0 8110 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13943_
timestamp 0
transform 1 0 7570 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13944_
timestamp 0
transform 1 0 10270 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13945_
timestamp 0
transform 1 0 10130 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__13946_
timestamp 0
transform -1 0 10310 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13947_
timestamp 0
transform 1 0 10410 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13948_
timestamp 0
transform 1 0 10570 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__13949_
timestamp 0
transform 1 0 10470 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13950_
timestamp 0
transform 1 0 10190 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13951_
timestamp 0
transform 1 0 8230 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13952_
timestamp 0
transform 1 0 9490 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13953_
timestamp 0
transform 1 0 9950 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13954_
timestamp 0
transform 1 0 9350 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13955_
timestamp 0
transform -1 0 10270 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13956_
timestamp 0
transform -1 0 10110 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13957_
timestamp 0
transform 1 0 10710 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13958_
timestamp 0
transform 1 0 10390 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13959_
timestamp 0
transform 1 0 10570 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13960_
timestamp 0
transform 1 0 9750 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13961_
timestamp 0
transform -1 0 8050 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13962_
timestamp 0
transform 1 0 9230 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13963_
timestamp 0
transform -1 0 9110 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13964_
timestamp 0
transform -1 0 9350 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13965_
timestamp 0
transform 1 0 9070 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13966_
timestamp 0
transform 1 0 9590 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13967_
timestamp 0
transform -1 0 9170 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13968_
timestamp 0
transform 1 0 10190 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13969_
timestamp 0
transform 1 0 10050 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13970_
timestamp 0
transform -1 0 9110 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13971_
timestamp 0
transform 1 0 9810 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13972_
timestamp 0
transform -1 0 8810 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13973_
timestamp 0
transform -1 0 8530 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13974_
timestamp 0
transform 1 0 9330 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13975_
timestamp 0
transform 1 0 9170 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13976_
timestamp 0
transform -1 0 9650 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13977_
timestamp 0
transform -1 0 8690 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13978_
timestamp 0
transform -1 0 8210 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13979_
timestamp 0
transform -1 0 9890 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__13980_
timestamp 0
transform 1 0 8350 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0__13981_
timestamp 0
transform 1 0 9830 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13982_
timestamp 0
transform -1 0 9590 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__13983_
timestamp 0
transform 1 0 9670 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13984_
timestamp 0
transform -1 0 9550 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13985_
timestamp 0
transform 1 0 9170 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__13986_
timestamp 0
transform 1 0 9490 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__13987_
timestamp 0
transform 1 0 10290 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__13988_
timestamp 0
transform 1 0 10330 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13989_
timestamp 0
transform 1 0 10470 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__13990_
timestamp 0
transform 1 0 10350 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__13991_
timestamp 0
transform -1 0 10750 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13992_
timestamp 0
transform 1 0 9950 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0__13993_
timestamp 0
transform 1 0 10870 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13994_
timestamp 0
transform 1 0 10650 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__13995_
timestamp 0
transform 1 0 10610 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13996_
timestamp 0
transform 1 0 10330 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13997_
timestamp 0
transform -1 0 10470 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__13998_
timestamp 0
transform -1 0 10130 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__13999_
timestamp 0
transform -1 0 10430 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__14000_
timestamp 0
transform -1 0 9950 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__14001_
timestamp 0
transform 1 0 9770 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__14002_
timestamp 0
transform -1 0 9730 0 1 16090
box -6 -8 26 248
use FILL  FILL_0__14003_
timestamp 0
transform -1 0 9750 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__14004_
timestamp 0
transform -1 0 10250 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__14005_
timestamp 0
transform -1 0 10290 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__14006_
timestamp 0
transform -1 0 10130 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__14007_
timestamp 0
transform -1 0 10070 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__14008_
timestamp 0
transform 1 0 9970 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0__14009_
timestamp 0
transform -1 0 9930 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__14010_
timestamp 0
transform -1 0 9570 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__14011_
timestamp 0
transform -1 0 9630 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__14012_
timestamp 0
transform 1 0 9590 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__14013_
timestamp 0
transform -1 0 8650 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__14014_
timestamp 0
transform -1 0 9830 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__14015_
timestamp 0
transform -1 0 10510 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__14016_
timestamp 0
transform 1 0 10690 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__14017_
timestamp 0
transform -1 0 10630 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__14018_
timestamp 0
transform 1 0 10830 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__14019_
timestamp 0
transform -1 0 10690 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__14020_
timestamp 0
transform -1 0 10790 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__14021_
timestamp 0
transform 1 0 10970 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__14022_
timestamp 0
transform 1 0 11090 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__14023_
timestamp 0
transform -1 0 10530 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__14024_
timestamp 0
transform -1 0 10970 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__14025_
timestamp 0
transform 1 0 11210 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__14026_
timestamp 0
transform -1 0 10830 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__14027_
timestamp 0
transform 1 0 10390 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__14028_
timestamp 0
transform -1 0 9410 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__14029_
timestamp 0
transform -1 0 9710 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__14030_
timestamp 0
transform 1 0 10170 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__14031_
timestamp 0
transform -1 0 9770 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__14032_
timestamp 0
transform 1 0 8890 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__14033_
timestamp 0
transform 1 0 10210 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__14034_
timestamp 0
transform -1 0 10010 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__14035_
timestamp 0
transform 1 0 10050 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__14036_
timestamp 0
transform 1 0 10470 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__14037_
timestamp 0
transform -1 0 10630 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__14038_
timestamp 0
transform -1 0 10590 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__14039_
timestamp 0
transform 1 0 10590 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__14040_
timestamp 0
transform -1 0 10830 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__14041_
timestamp 0
transform 1 0 10830 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__14042_
timestamp 0
transform 1 0 10990 0 1 14650
box -6 -8 26 248
use FILL  FILL_0__14043_
timestamp 0
transform 1 0 10910 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__14044_
timestamp 0
transform -1 0 10870 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__14045_
timestamp 0
transform -1 0 10590 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__14046_
timestamp 0
transform 1 0 10710 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__14047_
timestamp 0
transform -1 0 10430 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__14048_
timestamp 0
transform -1 0 9930 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__14049_
timestamp 0
transform 1 0 9950 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__14050_
timestamp 0
transform -1 0 9750 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__14051_
timestamp 0
transform -1 0 9510 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__14052_
timestamp 0
transform -1 0 9810 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__14053_
timestamp 0
transform -1 0 9630 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__14054_
timestamp 0
transform 1 0 9650 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__14055_
timestamp 0
transform -1 0 9810 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__14056_
timestamp 0
transform 1 0 10430 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__14057_
timestamp 0
transform -1 0 9810 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__14058_
timestamp 0
transform 1 0 10710 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__14059_
timestamp 0
transform -1 0 9910 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__14060_
timestamp 0
transform -1 0 10430 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__14061_
timestamp 0
transform 1 0 10250 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__14062_
timestamp 0
transform 1 0 10130 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__14063_
timestamp 0
transform 1 0 9990 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0__14064_
timestamp 0
transform -1 0 10710 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__14065_
timestamp 0
transform 1 0 10430 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__14066_
timestamp 0
transform -1 0 10290 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__14067_
timestamp 0
transform -1 0 10150 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__14068_
timestamp 0
transform 1 0 9330 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__14069_
timestamp 0
transform 1 0 10810 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__14070_
timestamp 0
transform -1 0 10590 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__14071_
timestamp 0
transform -1 0 10070 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__14072_
timestamp 0
transform -1 0 10190 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__14073_
timestamp 0
transform 1 0 10530 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__14074_
timestamp 0
transform 1 0 10430 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__14075_
timestamp 0
transform 1 0 10450 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__14076_
timestamp 0
transform -1 0 10590 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__14077_
timestamp 0
transform -1 0 10350 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__14078_
timestamp 0
transform 1 0 10090 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__14079_
timestamp 0
transform -1 0 9090 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__14080_
timestamp 0
transform -1 0 9650 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__14081_
timestamp 0
transform 1 0 9350 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__14082_
timestamp 0
transform -1 0 9230 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__14083_
timestamp 0
transform 1 0 9490 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__14084_
timestamp 0
transform 1 0 10410 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__14085_
timestamp 0
transform -1 0 10050 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__14086_
timestamp 0
transform 1 0 10190 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__14087_
timestamp 0
transform -1 0 9910 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__14088_
timestamp 0
transform 1 0 9450 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__14089_
timestamp 0
transform 1 0 9250 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__14090_
timestamp 0
transform 1 0 11050 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__14091_
timestamp 0
transform 1 0 10910 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0__14092_
timestamp 0
transform 1 0 10030 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__14093_
timestamp 0
transform 1 0 9970 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__14094_
timestamp 0
transform -1 0 9890 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__14095_
timestamp 0
transform 1 0 9850 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__14096_
timestamp 0
transform -1 0 9770 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__14097_
timestamp 0
transform -1 0 9750 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__14098_
timestamp 0
transform -1 0 9630 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__14099_
timestamp 0
transform 1 0 8750 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__14100_
timestamp 0
transform 1 0 8410 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__14101_
timestamp 0
transform 1 0 8750 0 1 12730
box -6 -8 26 248
use FILL  FILL_0__14102_
timestamp 0
transform -1 0 10330 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__14103_
timestamp 0
transform 1 0 10290 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__14104_
timestamp 0
transform -1 0 9670 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__14105_
timestamp 0
transform -1 0 9810 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__14106_
timestamp 0
transform -1 0 9550 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__14107_
timestamp 0
transform -1 0 9490 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__14108_
timestamp 0
transform 1 0 9570 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__14109_
timestamp 0
transform 1 0 9710 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__14110_
timestamp 0
transform -1 0 9850 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__14111_
timestamp 0
transform 1 0 9310 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__14112_
timestamp 0
transform 1 0 9170 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__14113_
timestamp 0
transform 1 0 7570 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__14114_
timestamp 0
transform 1 0 9410 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__14115_
timestamp 0
transform 1 0 9270 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__14116_
timestamp 0
transform -1 0 9570 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__14117_
timestamp 0
transform 1 0 9690 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0__14118_
timestamp 0
transform -1 0 7850 0 1 12250
box -6 -8 26 248
use FILL  FILL_0__14119_
timestamp 0
transform -1 0 10130 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__14120_
timestamp 0
transform -1 0 10170 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__14121_
timestamp 0
transform 1 0 9830 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__14122_
timestamp 0
transform 1 0 9690 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__14123_
timestamp 0
transform -1 0 8410 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__14124_
timestamp 0
transform -1 0 8550 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__14125_
timestamp 0
transform 1 0 8090 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__14126_
timestamp 0
transform -1 0 8510 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__14127_
timestamp 0
transform 1 0 8630 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__14128_
timestamp 0
transform -1 0 8490 0 1 15130
box -6 -8 26 248
use FILL  FILL_0__14129_
timestamp 0
transform 1 0 9150 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__14130_
timestamp 0
transform 1 0 8990 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__14131_
timestamp 0
transform -1 0 10210 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__14132_
timestamp 0
transform 1 0 10130 0 1 13690
box -6 -8 26 248
use FILL  FILL_0__14133_
timestamp 0
transform -1 0 10930 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__14134_
timestamp 0
transform 1 0 10770 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__14135_
timestamp 0
transform -1 0 8430 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__14136_
timestamp 0
transform -1 0 9190 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__14137_
timestamp 0
transform 1 0 9010 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__14138_
timestamp 0
transform 1 0 7910 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__14139_
timestamp 0
transform -1 0 9050 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__14140_
timestamp 0
transform 1 0 8870 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0__14141_
timestamp 0
transform 1 0 7670 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__14142_
timestamp 0
transform 1 0 7610 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__14143_
timestamp 0
transform 1 0 7790 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__14144_
timestamp 0
transform -1 0 7790 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__14145_
timestamp 0
transform -1 0 6550 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__14146_
timestamp 0
transform 1 0 6390 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__14147_
timestamp 0
transform 1 0 7530 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__14148_
timestamp 0
transform 1 0 7130 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__14149_
timestamp 0
transform -1 0 7450 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0__14150_
timestamp 0
transform -1 0 7550 0 1 14170
box -6 -8 26 248
use FILL  FILL_0__14151_
timestamp 0
transform -1 0 7590 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__14152_
timestamp 0
transform -1 0 7750 0 1 13210
box -6 -8 26 248
use FILL  FILL_0__14153_
timestamp 0
transform 1 0 7150 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0__14154_
timestamp 0
transform -1 0 6950 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__14155_
timestamp 0
transform 1 0 7410 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0__14156_
timestamp 0
transform 1 0 7230 0 1 15610
box -6 -8 26 248
use FILL  FILL_0__14157_
timestamp 0
transform -1 0 11070 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__14158_
timestamp 0
transform 1 0 10910 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0__14216_
timestamp 0
transform 1 0 7450 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__14217_
timestamp 0
transform 1 0 7670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__14218_
timestamp 0
transform -1 0 7690 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14219_
timestamp 0
transform -1 0 7510 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14220_
timestamp 0
transform 1 0 7630 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14221_
timestamp 0
transform 1 0 7490 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14222_
timestamp 0
transform -1 0 7410 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14223_
timestamp 0
transform -1 0 6890 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14224_
timestamp 0
transform 1 0 7010 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14225_
timestamp 0
transform 1 0 6810 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__14226_
timestamp 0
transform -1 0 7190 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__14227_
timestamp 0
transform 1 0 7150 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14228_
timestamp 0
transform -1 0 8510 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__14229_
timestamp 0
transform 1 0 7930 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__14230_
timestamp 0
transform -1 0 8350 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__14231_
timestamp 0
transform -1 0 10210 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__14232_
timestamp 0
transform -1 0 9930 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__14233_
timestamp 0
transform -1 0 10070 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__14234_
timestamp 0
transform -1 0 8970 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__14235_
timestamp 0
transform 1 0 8510 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__14236_
timestamp 0
transform 1 0 8410 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__14237_
timestamp 0
transform -1 0 8850 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__14238_
timestamp 0
transform -1 0 7870 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__14239_
timestamp 0
transform -1 0 7990 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__14240_
timestamp 0
transform -1 0 8430 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__14241_
timestamp 0
transform -1 0 8310 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__14242_
timestamp 0
transform -1 0 8270 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__14243_
timestamp 0
transform -1 0 8350 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14244_
timestamp 0
transform 1 0 6870 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14245_
timestamp 0
transform -1 0 6750 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14246_
timestamp 0
transform 1 0 9450 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14247_
timestamp 0
transform 1 0 8690 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__14248_
timestamp 0
transform 1 0 8550 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__14249_
timestamp 0
transform 1 0 9790 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__14250_
timestamp 0
transform 1 0 9970 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14251_
timestamp 0
transform 1 0 9810 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14252_
timestamp 0
transform 1 0 7570 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__14253_
timestamp 0
transform 1 0 7790 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__14254_
timestamp 0
transform 1 0 7630 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14255_
timestamp 0
transform 1 0 7490 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14256_
timestamp 0
transform 1 0 7130 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14257_
timestamp 0
transform -1 0 8090 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14258_
timestamp 0
transform 1 0 7030 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__14259_
timestamp 0
transform -1 0 7150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__14260_
timestamp 0
transform 1 0 7290 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14261_
timestamp 0
transform 1 0 7710 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14262_
timestamp 0
transform 1 0 7570 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14263_
timestamp 0
transform -1 0 7790 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14264_
timestamp 0
transform 1 0 6990 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14265_
timestamp 0
transform -1 0 7010 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14266_
timestamp 0
transform -1 0 6910 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__14267_
timestamp 0
transform -1 0 7150 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14268_
timestamp 0
transform -1 0 6870 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14269_
timestamp 0
transform 1 0 7050 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__14270_
timestamp 0
transform 1 0 6890 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__14271_
timestamp 0
transform -1 0 7290 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14272_
timestamp 0
transform -1 0 7430 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14273_
timestamp 0
transform 1 0 7530 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14274_
timestamp 0
transform -1 0 7710 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14275_
timestamp 0
transform 1 0 7250 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14276_
timestamp 0
transform -1 0 7690 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14277_
timestamp 0
transform -1 0 7910 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14278_
timestamp 0
transform -1 0 7950 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14279_
timestamp 0
transform 1 0 9290 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14280_
timestamp 0
transform -1 0 9230 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14281_
timestamp 0
transform 1 0 8010 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14282_
timestamp 0
transform -1 0 9350 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14283_
timestamp 0
transform 1 0 9430 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14284_
timestamp 0
transform 1 0 8250 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14285_
timestamp 0
transform -1 0 8390 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14286_
timestamp 0
transform 1 0 8190 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__14287_
timestamp 0
transform -1 0 9150 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14288_
timestamp 0
transform 1 0 8210 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14289_
timestamp 0
transform 1 0 8050 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14290_
timestamp 0
transform 1 0 7910 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14291_
timestamp 0
transform -1 0 8070 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14292_
timestamp 0
transform -1 0 8170 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14293_
timestamp 0
transform 1 0 9190 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14294_
timestamp 0
transform -1 0 9210 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14295_
timestamp 0
transform 1 0 8950 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14296_
timestamp 0
transform 1 0 9070 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14297_
timestamp 0
transform 1 0 9050 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14298_
timestamp 0
transform -1 0 9110 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14299_
timestamp 0
transform -1 0 8810 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14300_
timestamp 0
transform -1 0 9090 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14301_
timestamp 0
transform 1 0 7810 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__14302_
timestamp 0
transform -1 0 8830 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14303_
timestamp 0
transform -1 0 8870 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14304_
timestamp 0
transform -1 0 8970 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14305_
timestamp 0
transform 1 0 8670 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14306_
timestamp 0
transform -1 0 8810 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14307_
timestamp 0
transform 1 0 8710 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14308_
timestamp 0
transform 1 0 8110 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14309_
timestamp 0
transform 1 0 9350 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14310_
timestamp 0
transform -1 0 8310 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14311_
timestamp 0
transform -1 0 8330 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14312_
timestamp 0
transform 1 0 8450 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14313_
timestamp 0
transform -1 0 9630 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14314_
timestamp 0
transform -1 0 9510 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14315_
timestamp 0
transform 1 0 9550 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14316_
timestamp 0
transform 1 0 8650 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14317_
timestamp 0
transform -1 0 8670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__14318_
timestamp 0
transform 1 0 8410 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14319_
timestamp 0
transform -1 0 9010 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14320_
timestamp 0
transform -1 0 9690 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14321_
timestamp 0
transform -1 0 8730 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14322_
timestamp 0
transform -1 0 8870 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14323_
timestamp 0
transform 1 0 8530 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14324_
timestamp 0
transform 1 0 8890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__14325_
timestamp 0
transform 1 0 8410 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14326_
timestamp 0
transform -1 0 8610 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14327_
timestamp 0
transform 1 0 8690 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14328_
timestamp 0
transform 1 0 8830 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14329_
timestamp 0
transform -1 0 8790 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__14330_
timestamp 0
transform 1 0 8990 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14331_
timestamp 0
transform -1 0 9150 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14332_
timestamp 0
transform -1 0 9270 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14333_
timestamp 0
transform 1 0 8930 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14334_
timestamp 0
transform -1 0 9690 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__14335_
timestamp 0
transform -1 0 8630 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__14336_
timestamp 0
transform 1 0 8490 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__14337_
timestamp 0
transform -1 0 8390 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__14338_
timestamp 0
transform 1 0 8830 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__14339_
timestamp 0
transform 1 0 8990 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__14340_
timestamp 0
transform -1 0 8990 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__14341_
timestamp 0
transform -1 0 8850 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__14342_
timestamp 0
transform 1 0 9110 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__14343_
timestamp 0
transform 1 0 8690 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__14344_
timestamp 0
transform 1 0 8950 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__14345_
timestamp 0
transform 1 0 9270 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__14346_
timestamp 0
transform 1 0 9390 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__14347_
timestamp 0
transform -1 0 9550 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__14348_
timestamp 0
transform 1 0 7990 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14349_
timestamp 0
transform 1 0 7830 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14350_
timestamp 0
transform -1 0 8150 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14351_
timestamp 0
transform -1 0 7670 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14352_
timestamp 0
transform -1 0 7430 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14353_
timestamp 0
transform -1 0 7530 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14354_
timestamp 0
transform -1 0 7990 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14355_
timestamp 0
transform 1 0 7830 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14356_
timestamp 0
transform 1 0 8270 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14357_
timestamp 0
transform -1 0 8290 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14358_
timestamp 0
transform 1 0 8290 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14359_
timestamp 0
transform 1 0 8410 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14360_
timestamp 0
transform -1 0 8410 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14361_
timestamp 0
transform 1 0 8430 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14362_
timestamp 0
transform 1 0 7530 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__14363_
timestamp 0
transform 1 0 8110 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14364_
timestamp 0
transform -1 0 8010 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14365_
timestamp 0
transform -1 0 7870 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14366_
timestamp 0
transform 1 0 8010 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14367_
timestamp 0
transform 1 0 7290 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14368_
timestamp 0
transform -1 0 9390 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14369_
timestamp 0
transform 1 0 8550 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14370_
timestamp 0
transform 1 0 8530 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14371_
timestamp 0
transform -1 0 9630 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14372_
timestamp 0
transform -1 0 10810 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14373_
timestamp 0
transform 1 0 8650 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14374_
timestamp 0
transform 1 0 10330 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14375_
timestamp 0
transform 1 0 10350 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14376_
timestamp 0
transform 1 0 8850 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__14377_
timestamp 0
transform 1 0 9970 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14378_
timestamp 0
transform 1 0 10930 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14379_
timestamp 0
transform 1 0 11250 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14380_
timestamp 0
transform -1 0 11110 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14381_
timestamp 0
transform 1 0 11010 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14382_
timestamp 0
transform 1 0 9490 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14383_
timestamp 0
transform -1 0 10190 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14384_
timestamp 0
transform 1 0 10470 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14385_
timestamp 0
transform 1 0 10690 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14386_
timestamp 0
transform -1 0 10770 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14387_
timestamp 0
transform 1 0 10610 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14388_
timestamp 0
transform -1 0 10530 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14389_
timestamp 0
transform 1 0 9050 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__14390_
timestamp 0
transform -1 0 10310 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14391_
timestamp 0
transform 1 0 10450 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14392_
timestamp 0
transform 1 0 10590 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14393_
timestamp 0
transform 1 0 11030 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14394_
timestamp 0
transform -1 0 10890 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14395_
timestamp 0
transform 1 0 10650 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14396_
timestamp 0
transform 1 0 9550 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14397_
timestamp 0
transform 1 0 9750 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14398_
timestamp 0
transform -1 0 9950 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14399_
timestamp 0
transform 1 0 10550 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14400_
timestamp 0
transform -1 0 9990 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14401_
timestamp 0
transform 1 0 9970 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14402_
timestamp 0
transform 1 0 10050 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14403_
timestamp 0
transform 1 0 10110 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14404_
timestamp 0
transform -1 0 8930 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__14405_
timestamp 0
transform -1 0 9150 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14406_
timestamp 0
transform 1 0 10230 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14407_
timestamp 0
transform 1 0 9830 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__14408_
timestamp 0
transform -1 0 8850 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14409_
timestamp 0
transform -1 0 8990 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14410_
timestamp 0
transform 1 0 8670 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14411_
timestamp 0
transform -1 0 10410 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14412_
timestamp 0
transform 1 0 10110 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14413_
timestamp 0
transform 1 0 10230 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14414_
timestamp 0
transform 1 0 9070 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14415_
timestamp 0
transform 1 0 8870 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__14416_
timestamp 0
transform 1 0 9830 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14417_
timestamp 0
transform 1 0 9410 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14418_
timestamp 0
transform -1 0 9230 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14419_
timestamp 0
transform -1 0 9410 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14420_
timestamp 0
transform 1 0 9770 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14421_
timestamp 0
transform -1 0 8150 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__14422_
timestamp 0
transform -1 0 8270 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__14423_
timestamp 0
transform 1 0 8950 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__14424_
timestamp 0
transform 1 0 9250 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__14425_
timestamp 0
transform 1 0 9570 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14426_
timestamp 0
transform -1 0 8970 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__14427_
timestamp 0
transform 1 0 9690 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__14428_
timestamp 0
transform -1 0 10030 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14429_
timestamp 0
transform -1 0 9890 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__14430_
timestamp 0
transform 1 0 9770 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14431_
timestamp 0
transform -1 0 9930 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14432_
timestamp 0
transform 1 0 9890 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14433_
timestamp 0
transform 1 0 8010 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__14434_
timestamp 0
transform -1 0 8390 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__14435_
timestamp 0
transform 1 0 8470 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__14436_
timestamp 0
transform 1 0 7870 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__14437_
timestamp 0
transform -1 0 8110 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__14438_
timestamp 0
transform -1 0 8350 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__14439_
timestamp 0
transform 1 0 8450 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__14440_
timestamp 0
transform 1 0 9110 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__14441_
timestamp 0
transform -1 0 9130 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__14442_
timestamp 0
transform 1 0 8290 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__14443_
timestamp 0
transform -1 0 8450 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__14444_
timestamp 0
transform 1 0 8990 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__14445_
timestamp 0
transform -1 0 8750 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__14446_
timestamp 0
transform 1 0 8870 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__14447_
timestamp 0
transform 1 0 8630 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__14448_
timestamp 0
transform 1 0 8490 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__14449_
timestamp 0
transform 1 0 7990 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__14450_
timestamp 0
transform 1 0 9050 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__14451_
timestamp 0
transform 1 0 8910 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__14452_
timestamp 0
transform 1 0 8850 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__14453_
timestamp 0
transform 1 0 8270 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__14454_
timestamp 0
transform 1 0 8110 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__14455_
timestamp 0
transform 1 0 8570 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14456_
timestamp 0
transform 1 0 8530 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__14457_
timestamp 0
transform 1 0 8230 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__14458_
timestamp 0
transform 1 0 8330 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__14459_
timestamp 0
transform 1 0 8110 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__14460_
timestamp 0
transform -1 0 7990 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__14461_
timestamp 0
transform 1 0 8150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__14462_
timestamp 0
transform 1 0 8010 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__14463_
timestamp 0
transform 1 0 8190 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__14464_
timestamp 0
transform -1 0 7930 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__14465_
timestamp 0
transform -1 0 8070 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__14466_
timestamp 0
transform -1 0 7710 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__14467_
timestamp 0
transform -1 0 7870 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__14468_
timestamp 0
transform 1 0 7870 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__14469_
timestamp 0
transform 1 0 7730 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__14470_
timestamp 0
transform -1 0 7350 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__14471_
timestamp 0
transform 1 0 7130 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__14472_
timestamp 0
transform 1 0 9330 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__14473_
timestamp 0
transform 1 0 9170 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__14474_
timestamp 0
transform 1 0 7750 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__14475_
timestamp 0
transform -1 0 7990 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__14476_
timestamp 0
transform 1 0 9450 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__14477_
timestamp 0
transform -1 0 9110 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__14478_
timestamp 0
transform -1 0 9230 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__14479_
timestamp 0
transform -1 0 7770 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__14480_
timestamp 0
transform 1 0 9690 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__14481_
timestamp 0
transform 1 0 9550 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__14482_
timestamp 0
transform 1 0 9950 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__14483_
timestamp 0
transform 1 0 9790 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__14484_
timestamp 0
transform 1 0 9890 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__14485_
timestamp 0
transform 1 0 9490 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__14486_
timestamp 0
transform 1 0 9830 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__14487_
timestamp 0
transform 1 0 9850 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__14488_
timestamp 0
transform -1 0 9510 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__14489_
timestamp 0
transform 1 0 9350 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__14490_
timestamp 0
transform 1 0 8370 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__14491_
timestamp 0
transform -1 0 8550 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__14492_
timestamp 0
transform 1 0 8210 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__14493_
timestamp 0
transform 1 0 8070 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__14494_
timestamp 0
transform -1 0 7470 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__14495_
timestamp 0
transform -1 0 7610 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__14496_
timestamp 0
transform 1 0 7390 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__14497_
timestamp 0
transform -1 0 7310 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__14498_
timestamp 0
transform 1 0 9530 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__14499_
timestamp 0
transform -1 0 9550 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__14556_
timestamp 0
transform -1 0 14730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__14557_
timestamp 0
transform -1 0 14470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__14558_
timestamp 0
transform -1 0 14030 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14559_
timestamp 0
transform -1 0 12910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14560_
timestamp 0
transform -1 0 12130 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14561_
timestamp 0
transform -1 0 13050 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14562_
timestamp 0
transform 1 0 11690 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14563_
timestamp 0
transform -1 0 11990 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14564_
timestamp 0
transform -1 0 12510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14565_
timestamp 0
transform -1 0 12630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14566_
timestamp 0
transform -1 0 14550 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14567_
timestamp 0
transform -1 0 14570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__14568_
timestamp 0
transform -1 0 15450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__14569_
timestamp 0
transform 1 0 15050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__14570_
timestamp 0
transform 1 0 15030 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__14571_
timestamp 0
transform 1 0 14050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__14572_
timestamp 0
transform -1 0 14110 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__14573_
timestamp 0
transform -1 0 12490 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14574_
timestamp 0
transform 1 0 11630 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14575_
timestamp 0
transform 1 0 11830 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14576_
timestamp 0
transform -1 0 13310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14577_
timestamp 0
transform -1 0 13150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14578_
timestamp 0
transform 1 0 12990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14579_
timestamp 0
transform -1 0 13390 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14580_
timestamp 0
transform -1 0 12970 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14581_
timestamp 0
transform 1 0 14310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__14582_
timestamp 0
transform -1 0 14190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__14583_
timestamp 0
transform -1 0 13790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__14584_
timestamp 0
transform -1 0 13910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__14585_
timestamp 0
transform -1 0 12350 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14586_
timestamp 0
transform -1 0 9730 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14587_
timestamp 0
transform -1 0 9990 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14588_
timestamp 0
transform 1 0 10010 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14589_
timestamp 0
transform -1 0 9890 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14590_
timestamp 0
transform 1 0 9850 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14591_
timestamp 0
transform -1 0 11970 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14592_
timestamp 0
transform 1 0 11950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14593_
timestamp 0
transform 1 0 13010 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14594_
timestamp 0
transform -1 0 13930 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14595_
timestamp 0
transform 1 0 11270 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14596_
timestamp 0
transform 1 0 14250 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__14597_
timestamp 0
transform -1 0 14910 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__14598_
timestamp 0
transform 1 0 13770 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14599_
timestamp 0
transform -1 0 12790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14600_
timestamp 0
transform -1 0 12930 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14601_
timestamp 0
transform -1 0 11830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14602_
timestamp 0
transform 1 0 14890 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14603_
timestamp 0
transform 1 0 15290 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14604_
timestamp 0
transform 1 0 15150 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14605_
timestamp 0
transform -1 0 15010 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14606_
timestamp 0
transform -1 0 14550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14607_
timestamp 0
transform -1 0 14950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14608_
timestamp 0
transform -1 0 14830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14609_
timestamp 0
transform 1 0 15050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14610_
timestamp 0
transform -1 0 15750 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14611_
timestamp 0
transform 1 0 16010 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14612_
timestamp 0
transform 1 0 16150 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14613_
timestamp 0
transform 1 0 16290 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14614_
timestamp 0
transform 1 0 15890 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14615_
timestamp 0
transform 1 0 15170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14616_
timestamp 0
transform -1 0 15610 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14617_
timestamp 0
transform -1 0 14670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14618_
timestamp 0
transform 1 0 13710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14619_
timestamp 0
transform -1 0 13610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14620_
timestamp 0
transform 1 0 14310 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14621_
timestamp 0
transform -1 0 14190 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14622_
timestamp 0
transform 1 0 13890 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14623_
timestamp 0
transform -1 0 14050 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14624_
timestamp 0
transform -1 0 13770 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14625_
timestamp 0
transform -1 0 13930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14626_
timestamp 0
transform 1 0 13850 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14627_
timestamp 0
transform 1 0 14650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14628_
timestamp 0
transform -1 0 14550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14629_
timestamp 0
transform 1 0 14390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14630_
timestamp 0
transform 1 0 13970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14631_
timestamp 0
transform -1 0 14130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14632_
timestamp 0
transform -1 0 14270 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14633_
timestamp 0
transform -1 0 13870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14634_
timestamp 0
transform -1 0 13710 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14635_
timestamp 0
transform 1 0 14450 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14636_
timestamp 0
transform 1 0 14590 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14637_
timestamp 0
transform 1 0 14710 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14638_
timestamp 0
transform 1 0 14970 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14639_
timestamp 0
transform 1 0 15490 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14640_
timestamp 0
transform -1 0 15390 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14641_
timestamp 0
transform -1 0 15670 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14642_
timestamp 0
transform -1 0 14870 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14643_
timestamp 0
transform 1 0 15810 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14644_
timestamp 0
transform 1 0 15990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14645_
timestamp 0
transform -1 0 15890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14646_
timestamp 0
transform -1 0 15590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14647_
timestamp 0
transform 1 0 15730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14648_
timestamp 0
transform 1 0 16110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14649_
timestamp 0
transform -1 0 17030 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14650_
timestamp 0
transform 1 0 16850 0 1 16570
box -6 -8 26 248
use FILL  FILL_0__14651_
timestamp 0
transform 1 0 16930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14652_
timestamp 0
transform -1 0 16550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14653_
timestamp 0
transform 1 0 16390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14654_
timestamp 0
transform 1 0 16270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14655_
timestamp 0
transform -1 0 16790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14656_
timestamp 0
transform 1 0 16630 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14657_
timestamp 0
transform 1 0 16370 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14658_
timestamp 0
transform 1 0 16650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14659_
timestamp 0
transform -1 0 16490 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14660_
timestamp 0
transform 1 0 16070 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14661_
timestamp 0
transform 1 0 16230 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14662_
timestamp 0
transform -1 0 16870 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14663_
timestamp 0
transform 1 0 16990 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14664_
timestamp 0
transform 1 0 16630 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14665_
timestamp 0
transform 1 0 17010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14666_
timestamp 0
transform 1 0 16750 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14667_
timestamp 0
transform 1 0 16990 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14668_
timestamp 0
transform 1 0 16850 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14669_
timestamp 0
transform 1 0 16890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14670_
timestamp 0
transform -1 0 16610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14671_
timestamp 0
transform -1 0 16770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14672_
timestamp 0
transform -1 0 16710 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14673_
timestamp 0
transform -1 0 16070 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14674_
timestamp 0
transform -1 0 16330 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14675_
timestamp 0
transform 1 0 16190 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14676_
timestamp 0
transform 1 0 16090 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14677_
timestamp 0
transform -1 0 15950 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14678_
timestamp 0
transform 1 0 16250 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14679_
timestamp 0
transform 1 0 16230 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14680_
timestamp 0
transform -1 0 15970 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14681_
timestamp 0
transform 1 0 16470 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14682_
timestamp 0
transform -1 0 15930 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14683_
timestamp 0
transform 1 0 16610 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14684_
timestamp 0
transform -1 0 16550 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14685_
timestamp 0
transform 1 0 15930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14686_
timestamp 0
transform -1 0 16770 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14687_
timestamp 0
transform -1 0 16630 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14688_
timestamp 0
transform -1 0 16410 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14689_
timestamp 0
transform 1 0 16330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14690_
timestamp 0
transform -1 0 16470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14691_
timestamp 0
transform -1 0 15790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14692_
timestamp 0
transform -1 0 14330 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14693_
timestamp 0
transform 1 0 14430 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14694_
timestamp 0
transform -1 0 14750 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14695_
timestamp 0
transform -1 0 14930 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14696_
timestamp 0
transform 1 0 14650 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14697_
timestamp 0
transform 1 0 14790 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14698_
timestamp 0
transform -1 0 14830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14699_
timestamp 0
transform 1 0 14970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14700_
timestamp 0
transform -1 0 14610 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14701_
timestamp 0
transform 1 0 14810 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14702_
timestamp 0
transform -1 0 14530 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14703_
timestamp 0
transform -1 0 14290 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14704_
timestamp 0
transform -1 0 14410 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14705_
timestamp 0
transform 1 0 14950 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14706_
timestamp 0
transform 1 0 14190 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14707_
timestamp 0
transform -1 0 14090 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14708_
timestamp 0
transform -1 0 13950 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14709_
timestamp 0
transform 1 0 13990 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14710_
timestamp 0
transform 1 0 14130 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14711_
timestamp 0
transform -1 0 14630 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14712_
timestamp 0
transform 1 0 15090 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14713_
timestamp 0
transform 1 0 15230 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14714_
timestamp 0
transform 1 0 14970 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14715_
timestamp 0
transform 1 0 15110 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14716_
timestamp 0
transform -1 0 15530 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14717_
timestamp 0
transform 1 0 15650 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14718_
timestamp 0
transform -1 0 15530 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14719_
timestamp 0
transform -1 0 15290 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14720_
timestamp 0
transform 1 0 15510 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14721_
timestamp 0
transform 1 0 15390 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14722_
timestamp 0
transform 1 0 15430 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14723_
timestamp 0
transform -1 0 15310 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14724_
timestamp 0
transform -1 0 15810 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14725_
timestamp 0
transform -1 0 15690 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14726_
timestamp 0
transform -1 0 15650 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14727_
timestamp 0
transform 1 0 15770 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14728_
timestamp 0
transform 1 0 15390 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14729_
timestamp 0
transform 1 0 16070 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14730_
timestamp 0
transform 1 0 15930 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14731_
timestamp 0
transform 1 0 15790 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14732_
timestamp 0
transform 1 0 15970 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14733_
timestamp 0
transform -1 0 15850 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14734_
timestamp 0
transform 1 0 12730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14735_
timestamp 0
transform 1 0 14850 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14736_
timestamp 0
transform -1 0 15370 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14737_
timestamp 0
transform -1 0 15010 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14738_
timestamp 0
transform -1 0 15310 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14739_
timestamp 0
transform -1 0 15150 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14740_
timestamp 0
transform -1 0 14750 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14741_
timestamp 0
transform 1 0 14650 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14742_
timestamp 0
transform 1 0 12150 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14743_
timestamp 0
transform -1 0 12010 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14744_
timestamp 0
transform 1 0 11870 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14745_
timestamp 0
transform -1 0 12430 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14746_
timestamp 0
transform -1 0 12550 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14747_
timestamp 0
transform -1 0 12390 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14748_
timestamp 0
transform -1 0 12590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14749_
timestamp 0
transform -1 0 11650 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14750_
timestamp 0
transform -1 0 11750 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14751_
timestamp 0
transform -1 0 11230 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14752_
timestamp 0
transform 1 0 12130 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14753_
timestamp 0
transform 1 0 12270 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14754_
timestamp 0
transform -1 0 12090 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14755_
timestamp 0
transform 1 0 12210 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14756_
timestamp 0
transform -1 0 11810 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14757_
timestamp 0
transform -1 0 11950 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14758_
timestamp 0
transform 1 0 12690 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14759_
timestamp 0
transform -1 0 11370 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14760_
timestamp 0
transform -1 0 11490 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14761_
timestamp 0
transform 1 0 12690 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14762_
timestamp 0
transform 1 0 12410 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14763_
timestamp 0
transform -1 0 12290 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14764_
timestamp 0
transform 1 0 12550 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14765_
timestamp 0
transform 1 0 13390 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14766_
timestamp 0
transform 1 0 12830 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14767_
timestamp 0
transform 1 0 12970 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14768_
timestamp 0
transform 1 0 12750 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14769_
timestamp 0
transform -1 0 12770 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14770_
timestamp 0
transform 1 0 12830 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14771_
timestamp 0
transform -1 0 13590 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14772_
timestamp 0
transform 1 0 13450 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14773_
timestamp 0
transform -1 0 13850 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14774_
timestamp 0
transform -1 0 13710 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14775_
timestamp 0
transform -1 0 13130 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14776_
timestamp 0
transform -1 0 13270 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14777_
timestamp 0
transform 1 0 13950 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14778_
timestamp 0
transform -1 0 13350 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14779_
timestamp 0
transform -1 0 13190 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14780_
timestamp 0
transform -1 0 12910 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14781_
timestamp 0
transform -1 0 13050 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14782_
timestamp 0
transform 1 0 12970 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14783_
timestamp 0
transform 1 0 13250 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14784_
timestamp 0
transform -1 0 14370 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14785_
timestamp 0
transform 1 0 14870 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14786_
timestamp 0
transform 1 0 13550 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14787_
timestamp 0
transform 1 0 13550 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14788_
timestamp 0
transform 1 0 13110 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14789_
timestamp 0
transform 1 0 13390 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14790_
timestamp 0
transform -1 0 13710 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14791_
timestamp 0
transform 1 0 13950 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14792_
timestamp 0
transform -1 0 14090 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14793_
timestamp 0
transform -1 0 10950 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14794_
timestamp 0
transform 1 0 11070 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14795_
timestamp 0
transform 1 0 11470 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14796_
timestamp 0
transform 1 0 11590 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14797_
timestamp 0
transform 1 0 16130 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14798_
timestamp 0
transform 1 0 16050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14799_
timestamp 0
transform 1 0 16190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14800_
timestamp 0
transform -1 0 15650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14801_
timestamp 0
transform 1 0 14510 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14802_
timestamp 0
transform 1 0 13810 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14803_
timestamp 0
transform -1 0 14130 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14804_
timestamp 0
transform -1 0 14230 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14805_
timestamp 0
transform 1 0 11850 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14806_
timestamp 0
transform -1 0 11750 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14807_
timestamp 0
transform -1 0 11510 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14808_
timestamp 0
transform -1 0 11650 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14809_
timestamp 0
transform 1 0 11170 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14810_
timestamp 0
transform 1 0 10770 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14811_
timestamp 0
transform 1 0 10650 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14812_
timestamp 0
transform -1 0 10550 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14813_
timestamp 0
transform 1 0 11310 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14814_
timestamp 0
transform 1 0 11210 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14815_
timestamp 0
transform -1 0 11070 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14816_
timestamp 0
transform 1 0 11350 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14817_
timestamp 0
transform -1 0 11050 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14818_
timestamp 0
transform -1 0 10410 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14819_
timestamp 0
transform -1 0 10910 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14820_
timestamp 0
transform -1 0 10250 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14821_
timestamp 0
transform 1 0 10110 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14822_
timestamp 0
transform 1 0 10350 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14823_
timestamp 0
transform -1 0 9910 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14824_
timestamp 0
transform 1 0 10770 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14825_
timestamp 0
transform -1 0 10190 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14826_
timestamp 0
transform -1 0 10310 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14827_
timestamp 0
transform -1 0 10030 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14828_
timestamp 0
transform 1 0 9750 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14829_
timestamp 0
transform -1 0 10090 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14830_
timestamp 0
transform 1 0 10610 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14831_
timestamp 0
transform 1 0 10330 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14832_
timestamp 0
transform -1 0 10890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14833_
timestamp 0
transform 1 0 10630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14834_
timestamp 0
transform -1 0 9510 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14835_
timestamp 0
transform -1 0 9630 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14836_
timestamp 0
transform -1 0 9110 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14837_
timestamp 0
transform 1 0 9230 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14838_
timestamp 0
transform -1 0 9390 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14839_
timestamp 0
transform 1 0 10490 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14840_
timestamp 0
transform -1 0 10650 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14841_
timestamp 0
transform 1 0 10210 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14842_
timestamp 0
transform 1 0 10470 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14843_
timestamp 0
transform -1 0 10530 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14844_
timestamp 0
transform -1 0 12230 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14845_
timestamp 0
transform -1 0 12310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14846_
timestamp 0
transform 1 0 12350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14847_
timestamp 0
transform -1 0 11650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14848_
timestamp 0
transform -1 0 13450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14849_
timestamp 0
transform 1 0 11750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14850_
timestamp 0
transform -1 0 15250 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14851_
timestamp 0
transform 1 0 15430 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14852_
timestamp 0
transform -1 0 13630 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14853_
timestamp 0
transform -1 0 13310 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14854_
timestamp 0
transform 1 0 12810 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14855_
timestamp 0
transform 1 0 14370 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__14856_
timestamp 0
transform -1 0 12150 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14857_
timestamp 0
transform 1 0 12430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14858_
timestamp 0
transform 1 0 13010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14859_
timestamp 0
transform 1 0 13770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14860_
timestamp 0
transform -1 0 13470 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14861_
timestamp 0
transform 1 0 13390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__14862_
timestamp 0
transform 1 0 11990 0 1 730
box -6 -8 26 248
use FILL  FILL_0__14863_
timestamp 0
transform 1 0 12130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14864_
timestamp 0
transform 1 0 10750 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14865_
timestamp 0
transform -1 0 10910 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__14866_
timestamp 0
transform 1 0 11570 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14867_
timestamp 0
transform 1 0 10990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__14868_
timestamp 0
transform -1 0 11230 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__14908_
timestamp 0
transform -1 0 7590 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__14909_
timestamp 0
transform -1 0 30 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__14910_
timestamp 0
transform -1 0 8490 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14911_
timestamp 0
transform -1 0 9750 0 1 250
box -6 -8 26 248
use FILL  FILL_0__14912_
timestamp 0
transform -1 0 6770 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14913_
timestamp 0
transform -1 0 30 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__14914_
timestamp 0
transform 1 0 8210 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__14915_
timestamp 0
transform 1 0 16170 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__14916_
timestamp 0
transform 1 0 8410 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__14917_
timestamp 0
transform -1 0 7950 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__14918_
timestamp 0
transform -1 0 8090 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__14919_
timestamp 0
transform -1 0 6290 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__14920_
timestamp 0
transform 1 0 8970 0 -1 250
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert0
timestamp 0
transform 1 0 8190 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert1
timestamp 0
transform 1 0 9470 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert2
timestamp 0
transform -1 0 7830 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert3
timestamp 0
transform 1 0 9430 0 1 8410
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert4
timestamp 0
transform -1 0 9330 0 1 8410
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert5
timestamp 0
transform 1 0 5390 0 1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert6
timestamp 0
transform 1 0 4610 0 1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert7
timestamp 0
transform -1 0 1310 0 1 10810
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert8
timestamp 0
transform -1 0 1150 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert9
timestamp 0
transform 1 0 4510 0 1 6010
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert10
timestamp 0
transform 1 0 4110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert11
timestamp 0
transform 1 0 3570 0 1 6010
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert12
timestamp 0
transform -1 0 3290 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert13
timestamp 0
transform -1 0 4410 0 1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert14
timestamp 0
transform -1 0 4090 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert15
timestamp 0
transform 1 0 6830 0 1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert16
timestamp 0
transform -1 0 4770 0 1 7450
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert17
timestamp 0
transform -1 0 3210 0 1 7450
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert18
timestamp 0
transform -1 0 4510 0 1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert19
timestamp 0
transform -1 0 16130 0 1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert20
timestamp 0
transform -1 0 16250 0 1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert21
timestamp 0
transform -1 0 12870 0 1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert22
timestamp 0
transform -1 0 12090 0 1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert23
timestamp 0
transform -1 0 3010 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert24
timestamp 0
transform 1 0 4650 0 1 10330
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert25
timestamp 0
transform 1 0 1030 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert26
timestamp 0
transform -1 0 30 0 1 10810
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert27
timestamp 0
transform -1 0 1170 0 1 10810
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert28
timestamp 0
transform -1 0 30 0 1 10330
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert108
timestamp 0
transform -1 0 7790 0 1 7450
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert109
timestamp 0
transform 1 0 9270 0 1 7450
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert110
timestamp 0
transform -1 0 9010 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert111
timestamp 0
transform 1 0 8790 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert112
timestamp 0
transform 1 0 8290 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert113
timestamp 0
transform -1 0 13830 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert114
timestamp 0
transform -1 0 13510 0 1 13210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert115
timestamp 0
transform -1 0 14330 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert116
timestamp 0
transform 1 0 15070 0 1 14650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert117
timestamp 0
transform -1 0 6950 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert118
timestamp 0
transform 1 0 8130 0 1 6490
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert119
timestamp 0
transform 1 0 7690 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert120
timestamp 0
transform 1 0 7070 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert121
timestamp 0
transform -1 0 5790 0 1 6490
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert122
timestamp 0
transform -1 0 7570 0 1 6010
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert123
timestamp 0
transform 1 0 7730 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert124
timestamp 0
transform -1 0 6570 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert125
timestamp 0
transform -1 0 5990 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert126
timestamp 0
transform 1 0 5330 0 1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert127
timestamp 0
transform -1 0 4070 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert128
timestamp 0
transform 1 0 4590 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert129
timestamp 0
transform -1 0 4170 0 1 7450
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert130
timestamp 0
transform -1 0 5090 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert131
timestamp 0
transform -1 0 2550 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert132
timestamp 0
transform 1 0 2650 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert133
timestamp 0
transform 1 0 870 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert134
timestamp 0
transform -1 0 410 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert135
timestamp 0
transform 1 0 590 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert136
timestamp 0
transform 1 0 13570 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert137
timestamp 0
transform -1 0 11890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert138
timestamp 0
transform -1 0 12030 0 1 250
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert139
timestamp 0
transform 1 0 15490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert140
timestamp 0
transform 1 0 14530 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert141
timestamp 0
transform -1 0 10950 0 1 11290
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert142
timestamp 0
transform 1 0 12110 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert143
timestamp 0
transform -1 0 11290 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert144
timestamp 0
transform 1 0 12170 0 1 11290
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert145
timestamp 0
transform 1 0 12290 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert146
timestamp 0
transform -1 0 10510 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert147
timestamp 0
transform 1 0 10630 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert148
timestamp 0
transform 1 0 8470 0 1 250
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert149
timestamp 0
transform 1 0 8070 0 -1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert150
timestamp 0
transform -1 0 7910 0 1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert151
timestamp 0
transform -1 0 16050 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert152
timestamp 0
transform 1 0 16030 0 1 13690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert153
timestamp 0
transform -1 0 15910 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert154
timestamp 0
transform -1 0 15910 0 1 12730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert155
timestamp 0
transform -1 0 15970 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert156
timestamp 0
transform -1 0 15710 0 1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert157
timestamp 0
transform -1 0 15010 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert158
timestamp 0
transform 1 0 16930 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert159
timestamp 0
transform 1 0 15870 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert160
timestamp 0
transform 1 0 16390 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert161
timestamp 0
transform 1 0 11930 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert162
timestamp 0
transform 1 0 12710 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert163
timestamp 0
transform 1 0 12710 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert164
timestamp 0
transform -1 0 10510 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert165
timestamp 0
transform -1 0 11670 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert166
timestamp 0
transform -1 0 1170 0 1 9850
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert167
timestamp 0
transform -1 0 1130 0 1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert168
timestamp 0
transform 1 0 3630 0 1 9850
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert169
timestamp 0
transform 1 0 3690 0 1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert170
timestamp 0
transform 1 0 1490 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert171
timestamp 0
transform -1 0 14410 0 1 12730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert172
timestamp 0
transform 1 0 12830 0 1 12730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert173
timestamp 0
transform -1 0 11930 0 1 13690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert174
timestamp 0
transform -1 0 12090 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert175
timestamp 0
transform 1 0 14730 0 1 12250
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert176
timestamp 0
transform -1 0 14010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert177
timestamp 0
transform 1 0 15830 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert178
timestamp 0
transform -1 0 14030 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert179
timestamp 0
transform 1 0 15810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert180
timestamp 0
transform 1 0 15230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert181
timestamp 0
transform 1 0 11470 0 1 6490
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert182
timestamp 0
transform -1 0 10030 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert183
timestamp 0
transform 1 0 11710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert184
timestamp 0
transform 1 0 11790 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert185
timestamp 0
transform -1 0 10310 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert186
timestamp 0
transform -1 0 5990 0 1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert187
timestamp 0
transform 1 0 8210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert188
timestamp 0
transform -1 0 6810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert189
timestamp 0
transform -1 0 5950 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert190
timestamp 0
transform 1 0 9590 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert191
timestamp 0
transform 1 0 12490 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert192
timestamp 0
transform 1 0 12370 0 1 14650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert193
timestamp 0
transform 1 0 12110 0 1 15130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert194
timestamp 0
transform -1 0 11410 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert195
timestamp 0
transform -1 0 11830 0 1 14170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert196
timestamp 0
transform -1 0 1370 0 1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert197
timestamp 0
transform -1 0 1850 0 1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert198
timestamp 0
transform -1 0 710 0 1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert199
timestamp 0
transform 1 0 1870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert200
timestamp 0
transform 1 0 12730 0 1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert201
timestamp 0
transform -1 0 11870 0 1 10810
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert202
timestamp 0
transform 1 0 12810 0 1 10810
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert203
timestamp 0
transform -1 0 12590 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert204
timestamp 0
transform -1 0 12490 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert205
timestamp 0
transform 1 0 12030 0 1 5530
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert206
timestamp 0
transform 1 0 14010 0 1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert207
timestamp 0
transform -1 0 11810 0 1 5530
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert208
timestamp 0
transform 1 0 15470 0 1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert209
timestamp 0
transform 1 0 130 0 1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert210
timestamp 0
transform 1 0 1110 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert211
timestamp 0
transform 1 0 290 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert212
timestamp 0
transform -1 0 770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert213
timestamp 0
transform -1 0 30 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert214
timestamp 0
transform 1 0 6390 0 1 6970
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert215
timestamp 0
transform -1 0 5710 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert216
timestamp 0
transform -1 0 4790 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert217
timestamp 0
transform -1 0 3470 0 1 6970
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert218
timestamp 0
transform 1 0 6670 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert219
timestamp 0
transform -1 0 11550 0 1 5530
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert220
timestamp 0
transform 1 0 11730 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert221
timestamp 0
transform -1 0 12090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert222
timestamp 0
transform -1 0 9950 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert223
timestamp 0
transform 1 0 12270 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert224
timestamp 0
transform -1 0 8930 0 1 14170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert225
timestamp 0
transform 1 0 6930 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert226
timestamp 0
transform -1 0 10550 0 1 15610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert227
timestamp 0
transform -1 0 6830 0 1 15130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert228
timestamp 0
transform -1 0 7530 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert229
timestamp 0
transform 1 0 8950 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert230
timestamp 0
transform 1 0 8710 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert231
timestamp 0
transform -1 0 7430 0 1 16090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert232
timestamp 0
transform -1 0 8910 0 1 15130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert233
timestamp 0
transform -1 0 15130 0 1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert234
timestamp 0
transform 1 0 15350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert235
timestamp 0
transform -1 0 12910 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert236
timestamp 0
transform -1 0 12110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert237
timestamp 0
transform -1 0 13210 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert238
timestamp 0
transform -1 0 2270 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert239
timestamp 0
transform -1 0 4650 0 1 13210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert240
timestamp 0
transform 1 0 5190 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert241
timestamp 0
transform 1 0 5610 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert242
timestamp 0
transform 1 0 5390 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert243
timestamp 0
transform -1 0 1830 0 1 5530
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert244
timestamp 0
transform -1 0 1390 0 1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert245
timestamp 0
transform 1 0 4450 0 1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert246
timestamp 0
transform 1 0 2410 0 1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert247
timestamp 0
transform 1 0 3850 0 1 5530
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert248
timestamp 0
transform 1 0 2250 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert249
timestamp 0
transform 1 0 3230 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert250
timestamp 0
transform -1 0 430 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert251
timestamp 0
transform -1 0 1890 0 -1 15610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert252
timestamp 0
transform 1 0 3030 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert253
timestamp 0
transform 1 0 8610 0 1 6010
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert254
timestamp 0
transform 1 0 11350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert255
timestamp 0
transform -1 0 10210 0 1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert256
timestamp 0
transform 1 0 11090 0 1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert257
timestamp 0
transform 1 0 12030 0 1 6010
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert258
timestamp 0
transform -1 0 13970 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert259
timestamp 0
transform -1 0 13730 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert260
timestamp 0
transform 1 0 16450 0 1 15610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert261
timestamp 0
transform -1 0 15850 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert262
timestamp 0
transform -1 0 13430 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert263
timestamp 0
transform -1 0 13330 0 1 13690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert264
timestamp 0
transform 1 0 4530 0 1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert265
timestamp 0
transform 1 0 5410 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert266
timestamp 0
transform -1 0 4270 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert267
timestamp 0
transform -1 0 4390 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert268
timestamp 0
transform -1 0 4350 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert269
timestamp 0
transform -1 0 7510 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert270
timestamp 0
transform -1 0 7170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert271
timestamp 0
transform 1 0 9830 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert272
timestamp 0
transform 1 0 8050 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert273
timestamp 0
transform 1 0 8990 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert274
timestamp 0
transform -1 0 8250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert275
timestamp 0
transform 1 0 9850 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert276
timestamp 0
transform 1 0 9670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert277
timestamp 0
transform -1 0 7010 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert278
timestamp 0
transform 1 0 7430 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert279
timestamp 0
transform 1 0 9890 0 1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert280
timestamp 0
transform -1 0 15910 0 1 14170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert281
timestamp 0
transform -1 0 15850 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert282
timestamp 0
transform 1 0 15890 0 1 13690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert283
timestamp 0
transform -1 0 16570 0 1 14170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert284
timestamp 0
transform 1 0 16070 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert285
timestamp 0
transform -1 0 15850 0 1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert286
timestamp 0
transform -1 0 16310 0 1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert287
timestamp 0
transform 1 0 16350 0 1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert288
timestamp 0
transform 1 0 15050 0 1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert289
timestamp 0
transform -1 0 12990 0 1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert290
timestamp 0
transform 1 0 6710 0 1 12730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert291
timestamp 0
transform 1 0 6570 0 1 12730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert292
timestamp 0
transform -1 0 6470 0 1 12730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert293
timestamp 0
transform 1 0 8270 0 1 12730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert294
timestamp 0
transform -1 0 11850 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert295
timestamp 0
transform -1 0 11870 0 1 10330
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert296
timestamp 0
transform 1 0 15210 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert297
timestamp 0
transform 1 0 14990 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert298
timestamp 0
transform 1 0 17050 0 1 10330
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert299
timestamp 0
transform 1 0 16890 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert300
timestamp 0
transform 1 0 9090 0 1 14650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert301
timestamp 0
transform -1 0 7970 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert302
timestamp 0
transform -1 0 8050 0 1 14650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert303
timestamp 0
transform -1 0 8030 0 1 12730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert304
timestamp 0
transform -1 0 8550 0 1 6970
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert305
timestamp 0
transform 1 0 8590 0 1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert306
timestamp 0
transform -1 0 9670 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert307
timestamp 0
transform 1 0 9690 0 1 6970
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert308
timestamp 0
transform 1 0 10190 0 1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert309
timestamp 0
transform -1 0 13630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert310
timestamp 0
transform 1 0 13730 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert311
timestamp 0
transform -1 0 15890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert312
timestamp 0
transform -1 0 15970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert313
timestamp 0
transform -1 0 15070 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert314
timestamp 0
transform 1 0 15590 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert315
timestamp 0
transform 1 0 16370 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert316
timestamp 0
transform 1 0 14230 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert317
timestamp 0
transform 1 0 16350 0 1 5530
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert318
timestamp 0
transform -1 0 11670 0 1 5530
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert319
timestamp 0
transform 1 0 11910 0 1 5530
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert320
timestamp 0
transform 1 0 8550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert321
timestamp 0
transform -1 0 6930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert322
timestamp 0
transform 1 0 7010 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert323
timestamp 0
transform 1 0 8630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert324
timestamp 0
transform -1 0 630 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert325
timestamp 0
transform 1 0 2950 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert326
timestamp 0
transform 1 0 2070 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert327
timestamp 0
transform -1 0 2870 0 1 15130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert328
timestamp 0
transform 1 0 1030 0 1 15610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert329
timestamp 0
transform 1 0 2050 0 1 16570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert330
timestamp 0
transform -1 0 2830 0 1 15610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert331
timestamp 0
transform 1 0 3730 0 1 14170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert332
timestamp 0
transform -1 0 2810 0 1 12730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert333
timestamp 0
transform -1 0 1790 0 1 15130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert334
timestamp 0
transform 1 0 2790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert335
timestamp 0
transform 1 0 2550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert336
timestamp 0
transform 1 0 290 0 1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert337
timestamp 0
transform -1 0 1150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert338
timestamp 0
transform -1 0 1510 0 1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert339
timestamp 0
transform -1 0 790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert340
timestamp 0
transform 1 0 290 0 1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert341
timestamp 0
transform -1 0 530 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert342
timestamp 0
transform 1 0 1170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert343
timestamp 0
transform 1 0 170 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert344
timestamp 0
transform -1 0 30 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert345
timestamp 0
transform 1 0 10850 0 -1 16570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert346
timestamp 0
transform -1 0 11050 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert347
timestamp 0
transform 1 0 11470 0 1 15130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert348
timestamp 0
transform -1 0 10910 0 1 13690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert349
timestamp 0
transform 1 0 8070 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert350
timestamp 0
transform -1 0 7790 0 -1 16090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert351
timestamp 0
transform -1 0 7610 0 1 15130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert352
timestamp 0
transform 1 0 7730 0 1 15130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert353
timestamp 0
transform 1 0 10710 0 -1 14650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert354
timestamp 0
transform -1 0 6450 0 1 16090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert355
timestamp 0
transform -1 0 9430 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert356
timestamp 0
transform 1 0 9430 0 1 16090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert357
timestamp 0
transform -1 0 7030 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert358
timestamp 0
transform 1 0 10750 0 1 13690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert359
timestamp 0
transform -1 0 9450 0 1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert360
timestamp 0
transform -1 0 7490 0 1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert361
timestamp 0
transform -1 0 6290 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert362
timestamp 0
transform -1 0 8150 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert363
timestamp 0
transform 1 0 6650 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert364
timestamp 0
transform 1 0 3450 0 1 11770
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert365
timestamp 0
transform -1 0 4790 0 1 13210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert366
timestamp 0
transform -1 0 3650 0 1 13210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert367
timestamp 0
transform -1 0 2950 0 -1 13210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert368
timestamp 0
transform -1 0 4730 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert369
timestamp 0
transform 1 0 13310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert370
timestamp 0
transform -1 0 12890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert371
timestamp 0
transform 1 0 12010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert372
timestamp 0
transform 1 0 13170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert373
timestamp 0
transform -1 0 11170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert374
timestamp 0
transform 1 0 2850 0 1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert375
timestamp 0
transform 1 0 2970 0 1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert376
timestamp 0
transform -1 0 1430 0 1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert377
timestamp 0
transform -1 0 1970 0 1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert378
timestamp 0
transform -1 0 1310 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert379
timestamp 0
transform 1 0 6330 0 1 11770
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert380
timestamp 0
transform 1 0 4910 0 1 13210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert381
timestamp 0
transform -1 0 2850 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert382
timestamp 0
transform 1 0 5730 0 1 11290
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert383
timestamp 0
transform -1 0 4490 0 1 11290
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert29
timestamp 0
transform -1 0 9390 0 1 4570
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert30
timestamp 0
transform 1 0 10450 0 1 16570
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert31
timestamp 0
transform -1 0 1730 0 1 5050
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert32
timestamp 0
transform -1 0 6190 0 1 12250
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert33
timestamp 0
transform -1 0 5770 0 -1 14170
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert34
timestamp 0
transform -1 0 10030 0 1 7450
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert35
timestamp 0
transform -1 0 13170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert36
timestamp 0
transform 1 0 3490 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert37
timestamp 0
transform -1 0 14670 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert38
timestamp 0
transform 1 0 5610 0 1 10810
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert39
timestamp 0
transform -1 0 5850 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert40
timestamp 0
transform 1 0 15870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert41
timestamp 0
transform -1 0 11290 0 1 3130
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert42
timestamp 0
transform 1 0 9450 0 1 11290
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert43
timestamp 0
transform 1 0 7350 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert44
timestamp 0
transform 1 0 2730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert45
timestamp 0
transform 1 0 11030 0 -1 15130
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert46
timestamp 0
transform 1 0 3470 0 1 6490
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert47
timestamp 0
transform 1 0 12970 0 1 7930
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert48
timestamp 0
transform -1 0 2070 0 -1 12730
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert49
timestamp 0
transform 1 0 6090 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert50
timestamp 0
transform -1 0 13470 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert51
timestamp 0
transform 1 0 14690 0 1 13690
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert52
timestamp 0
transform -1 0 7010 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert53
timestamp 0
transform -1 0 4230 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert54
timestamp 0
transform 1 0 13090 0 1 6970
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert55
timestamp 0
transform 1 0 14130 0 1 12730
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert56
timestamp 0
transform -1 0 11170 0 1 7930
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert57
timestamp 0
transform -1 0 14670 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert58
timestamp 0
transform 1 0 7130 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert59
timestamp 0
transform -1 0 5830 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert60
timestamp 0
transform -1 0 8830 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert61
timestamp 0
transform 1 0 6330 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert62
timestamp 0
transform 1 0 11170 0 1 7450
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert63
timestamp 0
transform 1 0 10310 0 1 12250
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert64
timestamp 0
transform 1 0 3770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert65
timestamp 0
transform 1 0 6910 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert66
timestamp 0
transform 1 0 10550 0 1 16090
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert67
timestamp 0
transform -1 0 15190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert68
timestamp 0
transform -1 0 6230 0 1 14170
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert69
timestamp 0
transform 1 0 6910 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert70
timestamp 0
transform 1 0 3010 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert71
timestamp 0
transform -1 0 2590 0 1 11770
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert72
timestamp 0
transform 1 0 9390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert73
timestamp 0
transform 1 0 12370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert74
timestamp 0
transform 1 0 15270 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert75
timestamp 0
transform 1 0 10310 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert76
timestamp 0
transform 1 0 8290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert77
timestamp 0
transform 1 0 11390 0 1 7930
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert78
timestamp 0
transform 1 0 10810 0 1 15610
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert79
timestamp 0
transform 1 0 11350 0 1 4570
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert80
timestamp 0
transform 1 0 4490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert81
timestamp 0
transform -1 0 5310 0 1 13210
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert82
timestamp 0
transform 1 0 11930 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert83
timestamp 0
transform -1 0 1790 0 1 6490
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert84
timestamp 0
transform 1 0 8430 0 1 11290
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert85
timestamp 0
transform -1 0 5270 0 -1 13690
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert86
timestamp 0
transform 1 0 12570 0 1 3130
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert87
timestamp 0
transform -1 0 12030 0 1 7450
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert88
timestamp 0
transform 1 0 8050 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert89
timestamp 0
transform 1 0 6490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert90
timestamp 0
transform -1 0 2770 0 1 13210
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert91
timestamp 0
transform -1 0 2110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert92
timestamp 0
transform 1 0 9350 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert93
timestamp 0
transform -1 0 2110 0 1 7450
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert94
timestamp 0
transform -1 0 4090 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert95
timestamp 0
transform -1 0 3070 0 1 11770
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert96
timestamp 0
transform -1 0 8970 0 1 5050
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert97
timestamp 0
transform -1 0 9230 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert98
timestamp 0
transform -1 0 8090 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert99
timestamp 0
transform -1 0 9890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert100
timestamp 0
transform 1 0 11610 0 1 4570
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert101
timestamp 0
transform -1 0 14910 0 -1 12250
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert102
timestamp 0
transform 1 0 12250 0 1 7450
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert103
timestamp 0
transform -1 0 10110 0 1 6970
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert104
timestamp 0
transform -1 0 6170 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert105
timestamp 0
transform -1 0 6570 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert106
timestamp 0
transform -1 0 2170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert107
timestamp 0
transform 1 0 9690 0 1 11290
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert384
timestamp 0
transform 1 0 8890 0 -1 17050
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert385
timestamp 0
transform -1 0 5550 0 1 6490
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert386
timestamp 0
transform -1 0 4650 0 1 5050
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert387
timestamp 0
transform 1 0 10750 0 1 7450
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert388
timestamp 0
transform -1 0 7830 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert389
timestamp 0
transform 1 0 8350 0 1 6010
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert390
timestamp 0
transform -1 0 10330 0 1 4570
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert391
timestamp 0
transform -1 0 7010 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__7072_
timestamp 0
transform 1 0 6150 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__7073_
timestamp 0
transform 1 0 8810 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7074_
timestamp 0
transform 1 0 6690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7075_
timestamp 0
transform 1 0 7650 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__7076_
timestamp 0
transform -1 0 5830 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7077_
timestamp 0
transform -1 0 8610 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7078_
timestamp 0
transform -1 0 5470 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7079_
timestamp 0
transform -1 0 6790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7080_
timestamp 0
transform -1 0 8610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7081_
timestamp 0
transform -1 0 5410 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7082_
timestamp 0
transform -1 0 6390 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7083_
timestamp 0
transform 1 0 5950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7084_
timestamp 0
transform 1 0 8670 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7085_
timestamp 0
transform 1 0 5830 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7086_
timestamp 0
transform -1 0 5610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7087_
timestamp 0
transform -1 0 5490 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7088_
timestamp 0
transform -1 0 5190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7089_
timestamp 0
transform -1 0 5350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7090_
timestamp 0
transform -1 0 7870 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7091_
timestamp 0
transform -1 0 5430 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7092_
timestamp 0
transform -1 0 5570 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7093_
timestamp 0
transform -1 0 5250 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7094_
timestamp 0
transform 1 0 5310 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7095_
timestamp 0
transform -1 0 5210 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7096_
timestamp 0
transform -1 0 5690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7097_
timestamp 0
transform -1 0 5810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7098_
timestamp 0
transform -1 0 5810 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7099_
timestamp 0
transform 1 0 5630 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7100_
timestamp 0
transform 1 0 5450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7101_
timestamp 0
transform 1 0 5370 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__7102_
timestamp 0
transform -1 0 5250 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__7103_
timestamp 0
transform 1 0 6390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7104_
timestamp 0
transform 1 0 5110 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__7105_
timestamp 0
transform 1 0 5330 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7106_
timestamp 0
transform 1 0 4970 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__7107_
timestamp 0
transform 1 0 4890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7108_
timestamp 0
transform 1 0 5950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7109_
timestamp 0
transform 1 0 5210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7110_
timestamp 0
transform -1 0 5350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7111_
timestamp 0
transform 1 0 5490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7112_
timestamp 0
transform -1 0 6230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7113_
timestamp 0
transform -1 0 5590 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7114_
timestamp 0
transform -1 0 10370 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7115_
timestamp 0
transform -1 0 8970 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__7116_
timestamp 0
transform -1 0 8830 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__7117_
timestamp 0
transform -1 0 10790 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7118_
timestamp 0
transform -1 0 9010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7119_
timestamp 0
transform 1 0 8650 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__7120_
timestamp 0
transform -1 0 8030 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__7121_
timestamp 0
transform -1 0 8090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7122_
timestamp 0
transform -1 0 7890 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__7123_
timestamp 0
transform -1 0 9450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7124_
timestamp 0
transform 1 0 9110 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__7125_
timestamp 0
transform -1 0 9250 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7126_
timestamp 0
transform 1 0 9250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7127_
timestamp 0
transform 1 0 9090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7128_
timestamp 0
transform 1 0 8770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7129_
timestamp 0
transform -1 0 8950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7130_
timestamp 0
transform 1 0 7450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7131_
timestamp 0
transform 1 0 8470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7132_
timestamp 0
transform 1 0 8450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7133_
timestamp 0
transform 1 0 7390 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7134_
timestamp 0
transform 1 0 13050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7135_
timestamp 0
transform 1 0 13270 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7136_
timestamp 0
transform 1 0 13110 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7137_
timestamp 0
transform 1 0 12010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7138_
timestamp 0
transform -1 0 10470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7139_
timestamp 0
transform -1 0 10850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7140_
timestamp 0
transform 1 0 10770 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7141_
timestamp 0
transform -1 0 9290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7142_
timestamp 0
transform -1 0 9010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7143_
timestamp 0
transform -1 0 9130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7144_
timestamp 0
transform -1 0 9270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7145_
timestamp 0
transform 1 0 9710 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7146_
timestamp 0
transform 1 0 9550 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7147_
timestamp 0
transform 1 0 9530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7148_
timestamp 0
transform -1 0 9990 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7149_
timestamp 0
transform 1 0 8350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7150_
timestamp 0
transform 1 0 8890 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7151_
timestamp 0
transform -1 0 7870 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7152_
timestamp 0
transform -1 0 9750 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7153_
timestamp 0
transform 1 0 9730 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7154_
timestamp 0
transform 1 0 11010 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7155_
timestamp 0
transform 1 0 7950 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7156_
timestamp 0
transform 1 0 7550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7157_
timestamp 0
transform -1 0 6490 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7158_
timestamp 0
transform -1 0 6470 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7159_
timestamp 0
transform 1 0 9330 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7160_
timestamp 0
transform -1 0 10170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7161_
timestamp 0
transform -1 0 10010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7162_
timestamp 0
transform 1 0 9190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7163_
timestamp 0
transform 1 0 7970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7164_
timestamp 0
transform -1 0 8610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7165_
timestamp 0
transform 1 0 8650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7166_
timestamp 0
transform 1 0 8830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7167_
timestamp 0
transform -1 0 9190 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7168_
timestamp 0
transform -1 0 9050 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7169_
timestamp 0
transform 1 0 8810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7170_
timestamp 0
transform -1 0 7610 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7171_
timestamp 0
transform -1 0 8630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7172_
timestamp 0
transform 1 0 11130 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7173_
timestamp 0
transform -1 0 9750 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7174_
timestamp 0
transform -1 0 9870 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7175_
timestamp 0
transform 1 0 8310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7176_
timestamp 0
transform 1 0 8490 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7177_
timestamp 0
transform 1 0 8330 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7178_
timestamp 0
transform -1 0 8370 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7179_
timestamp 0
transform 1 0 10330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7180_
timestamp 0
transform 1 0 9290 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7181_
timestamp 0
transform 1 0 9130 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7182_
timestamp 0
transform 1 0 9450 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7183_
timestamp 0
transform 1 0 8850 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7184_
timestamp 0
transform -1 0 8990 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7185_
timestamp 0
transform 1 0 8690 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7186_
timestamp 0
transform 1 0 8510 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7187_
timestamp 0
transform -1 0 8390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7188_
timestamp 0
transform -1 0 7990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7189_
timestamp 0
transform -1 0 8170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7190_
timestamp 0
transform 1 0 7810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7191_
timestamp 0
transform 1 0 10330 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7192_
timestamp 0
transform 1 0 9810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7193_
timestamp 0
transform -1 0 10170 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7194_
timestamp 0
transform 1 0 9570 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7195_
timestamp 0
transform 1 0 8510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7196_
timestamp 0
transform -1 0 7950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7197_
timestamp 0
transform 1 0 8090 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7198_
timestamp 0
transform 1 0 8090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7199_
timestamp 0
transform 1 0 8190 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7200_
timestamp 0
transform 1 0 8450 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7201_
timestamp 0
transform 1 0 8750 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7202_
timestamp 0
transform -1 0 8630 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7203_
timestamp 0
transform -1 0 6610 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7204_
timestamp 0
transform 1 0 7750 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__7205_
timestamp 0
transform 1 0 9390 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7206_
timestamp 0
transform 1 0 7950 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__7207_
timestamp 0
transform -1 0 6350 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7208_
timestamp 0
transform -1 0 7790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7209_
timestamp 0
transform -1 0 9850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7210_
timestamp 0
transform -1 0 8890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7211_
timestamp 0
transform -1 0 9690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7212_
timestamp 0
transform -1 0 9390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7213_
timestamp 0
transform 1 0 9510 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7214_
timestamp 0
transform 1 0 9050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7215_
timestamp 0
transform 1 0 8890 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7216_
timestamp 0
transform 1 0 9050 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7217_
timestamp 0
transform 1 0 9170 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7218_
timestamp 0
transform 1 0 9430 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7219_
timestamp 0
transform 1 0 9290 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7220_
timestamp 0
transform -1 0 8630 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7221_
timestamp 0
transform 1 0 8750 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7222_
timestamp 0
transform -1 0 8350 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7223_
timestamp 0
transform -1 0 7830 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7224_
timestamp 0
transform -1 0 7690 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7225_
timestamp 0
transform -1 0 7590 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7226_
timestamp 0
transform 1 0 7950 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7227_
timestamp 0
transform -1 0 7430 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7228_
timestamp 0
transform -1 0 7730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7229_
timestamp 0
transform -1 0 6130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7230_
timestamp 0
transform 1 0 6370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7231_
timestamp 0
transform -1 0 5910 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7232_
timestamp 0
transform 1 0 6270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7233_
timestamp 0
transform 1 0 8470 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7234_
timestamp 0
transform 1 0 8350 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7235_
timestamp 0
transform -1 0 6950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7236_
timestamp 0
transform -1 0 8730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7237_
timestamp 0
transform 1 0 11250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7238_
timestamp 0
transform -1 0 9330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7239_
timestamp 0
transform -1 0 9450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7240_
timestamp 0
transform 1 0 7790 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7241_
timestamp 0
transform 1 0 7630 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7242_
timestamp 0
transform 1 0 7970 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7243_
timestamp 0
transform -1 0 8090 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7244_
timestamp 0
transform -1 0 8190 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7245_
timestamp 0
transform 1 0 7310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7246_
timestamp 0
transform -1 0 6470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7247_
timestamp 0
transform 1 0 6370 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7248_
timestamp 0
transform 1 0 6510 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7249_
timestamp 0
transform 1 0 6370 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7250_
timestamp 0
transform -1 0 6170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7251_
timestamp 0
transform -1 0 6330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7252_
timestamp 0
transform 1 0 6410 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7253_
timestamp 0
transform 1 0 6410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7254_
timestamp 0
transform 1 0 8210 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7255_
timestamp 0
transform -1 0 8070 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7256_
timestamp 0
transform 1 0 6270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7257_
timestamp 0
transform -1 0 6290 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7258_
timestamp 0
transform -1 0 5770 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7259_
timestamp 0
transform -1 0 9830 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7260_
timestamp 0
transform -1 0 7930 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7261_
timestamp 0
transform -1 0 8050 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7262_
timestamp 0
transform -1 0 8230 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7263_
timestamp 0
transform 1 0 7570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7264_
timestamp 0
transform -1 0 7970 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7265_
timestamp 0
transform -1 0 6670 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7266_
timestamp 0
transform -1 0 6490 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7267_
timestamp 0
transform -1 0 5670 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7268_
timestamp 0
transform -1 0 5030 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7269_
timestamp 0
transform 1 0 5810 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7270_
timestamp 0
transform -1 0 5170 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7271_
timestamp 0
transform 1 0 4870 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7272_
timestamp 0
transform -1 0 5470 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7273_
timestamp 0
transform 1 0 5310 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7274_
timestamp 0
transform 1 0 5590 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7275_
timestamp 0
transform -1 0 5630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7276_
timestamp 0
transform -1 0 5990 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7277_
timestamp 0
transform 1 0 5810 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7278_
timestamp 0
transform 1 0 5730 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7279_
timestamp 0
transform 1 0 6110 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7280_
timestamp 0
transform 1 0 6570 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7281_
timestamp 0
transform -1 0 6230 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7282_
timestamp 0
transform -1 0 7410 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7283_
timestamp 0
transform 1 0 7450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7284_
timestamp 0
transform -1 0 7350 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7285_
timestamp 0
transform 1 0 6810 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7286_
timestamp 0
transform 1 0 6770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7287_
timestamp 0
transform -1 0 6090 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7288_
timestamp 0
transform -1 0 6590 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7289_
timestamp 0
transform -1 0 5550 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7290_
timestamp 0
transform -1 0 5650 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7291_
timestamp 0
transform -1 0 5790 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7292_
timestamp 0
transform 1 0 5930 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7293_
timestamp 0
transform 1 0 5950 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7294_
timestamp 0
transform 1 0 6030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7295_
timestamp 0
transform -1 0 7810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7296_
timestamp 0
transform 1 0 7890 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7297_
timestamp 0
transform -1 0 7290 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7298_
timestamp 0
transform 1 0 6050 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7299_
timestamp 0
transform 1 0 5390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7300_
timestamp 0
transform -1 0 4270 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7301_
timestamp 0
transform -1 0 5130 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7302_
timestamp 0
transform -1 0 7510 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7303_
timestamp 0
transform 1 0 7070 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7304_
timestamp 0
transform 1 0 6930 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7305_
timestamp 0
transform -1 0 4810 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7306_
timestamp 0
transform -1 0 4390 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7307_
timestamp 0
transform -1 0 5410 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7308_
timestamp 0
transform -1 0 4130 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7309_
timestamp 0
transform 1 0 3970 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7310_
timestamp 0
transform -1 0 4650 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7311_
timestamp 0
transform -1 0 4490 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7312_
timestamp 0
transform -1 0 4490 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7313_
timestamp 0
transform -1 0 4630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7314_
timestamp 0
transform -1 0 4750 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7315_
timestamp 0
transform 1 0 5490 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7316_
timestamp 0
transform -1 0 5490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7317_
timestamp 0
transform -1 0 5350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7318_
timestamp 0
transform 1 0 5670 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7319_
timestamp 0
transform 1 0 5530 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7320_
timestamp 0
transform 1 0 5490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7321_
timestamp 0
transform 1 0 5210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7322_
timestamp 0
transform -1 0 3830 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7323_
timestamp 0
transform 1 0 5810 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7324_
timestamp 0
transform -1 0 5890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7325_
timestamp 0
transform 1 0 5670 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7326_
timestamp 0
transform -1 0 5750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7327_
timestamp 0
transform -1 0 4750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7328_
timestamp 0
transform -1 0 6650 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7329_
timestamp 0
transform 1 0 5170 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7330_
timestamp 0
transform -1 0 7350 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7331_
timestamp 0
transform -1 0 7270 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7332_
timestamp 0
transform -1 0 7170 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7333_
timestamp 0
transform -1 0 7050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7334_
timestamp 0
transform -1 0 6230 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7335_
timestamp 0
transform -1 0 5090 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7336_
timestamp 0
transform -1 0 4970 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7337_
timestamp 0
transform -1 0 4970 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7338_
timestamp 0
transform -1 0 6090 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7339_
timestamp 0
transform 1 0 5330 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7340_
timestamp 0
transform 1 0 5550 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7341_
timestamp 0
transform 1 0 5390 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7342_
timestamp 0
transform 1 0 5270 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7343_
timestamp 0
transform -1 0 5010 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7344_
timestamp 0
transform -1 0 4890 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7345_
timestamp 0
transform -1 0 5070 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7346_
timestamp 0
transform 1 0 5130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7347_
timestamp 0
transform -1 0 5270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7348_
timestamp 0
transform 1 0 5310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7349_
timestamp 0
transform 1 0 5270 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7350_
timestamp 0
transform 1 0 5310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7351_
timestamp 0
transform 1 0 6150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7352_
timestamp 0
transform 1 0 5190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7353_
timestamp 0
transform -1 0 5270 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7354_
timestamp 0
transform 1 0 5390 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7355_
timestamp 0
transform -1 0 5430 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7356_
timestamp 0
transform 1 0 5930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7357_
timestamp 0
transform -1 0 6670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7358_
timestamp 0
transform -1 0 5830 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7359_
timestamp 0
transform -1 0 5550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7360_
timestamp 0
transform -1 0 5710 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7361_
timestamp 0
transform -1 0 5670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7362_
timestamp 0
transform 1 0 5530 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7363_
timestamp 0
transform 1 0 5970 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7364_
timestamp 0
transform 1 0 5790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7365_
timestamp 0
transform 1 0 6110 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7366_
timestamp 0
transform 1 0 6810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7367_
timestamp 0
transform -1 0 6830 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7368_
timestamp 0
transform -1 0 6310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7369_
timestamp 0
transform -1 0 6170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7370_
timestamp 0
transform -1 0 5990 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7371_
timestamp 0
transform 1 0 4990 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7372_
timestamp 0
transform -1 0 4910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7373_
timestamp 0
transform 1 0 4810 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7374_
timestamp 0
transform 1 0 5110 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7375_
timestamp 0
transform -1 0 5130 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7376_
timestamp 0
transform 1 0 6950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7377_
timestamp 0
transform -1 0 6670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7378_
timestamp 0
transform 1 0 7930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7379_
timestamp 0
transform 1 0 6070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7380_
timestamp 0
transform -1 0 6330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7381_
timestamp 0
transform 1 0 6510 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7382_
timestamp 0
transform 1 0 6430 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7383_
timestamp 0
transform 1 0 6550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7384_
timestamp 0
transform 1 0 6590 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7385_
timestamp 0
transform -1 0 7510 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7386_
timestamp 0
transform 1 0 6270 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7387_
timestamp 0
transform -1 0 6810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7388_
timestamp 0
transform -1 0 7070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7389_
timestamp 0
transform -1 0 7210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7390_
timestamp 0
transform -1 0 6450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7391_
timestamp 0
transform -1 0 6490 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7392_
timestamp 0
transform -1 0 6350 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7393_
timestamp 0
transform -1 0 5070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7394_
timestamp 0
transform 1 0 7290 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7395_
timestamp 0
transform -1 0 7070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7396_
timestamp 0
transform -1 0 7070 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7397_
timestamp 0
transform 1 0 6910 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7398_
timestamp 0
transform 1 0 6750 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7399_
timestamp 0
transform 1 0 8310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7400_
timestamp 0
transform -1 0 7190 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7401_
timestamp 0
transform -1 0 7310 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7402_
timestamp 0
transform 1 0 7210 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7403_
timestamp 0
transform 1 0 7570 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7404_
timestamp 0
transform 1 0 8430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7405_
timestamp 0
transform 1 0 8170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7406_
timestamp 0
transform 1 0 8030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7407_
timestamp 0
transform 1 0 7770 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7408_
timestamp 0
transform 1 0 7630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7409_
timestamp 0
transform 1 0 7350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7410_
timestamp 0
transform 1 0 7190 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7411_
timestamp 0
transform 1 0 7630 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7412_
timestamp 0
transform 1 0 6950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7413_
timestamp 0
transform 1 0 7350 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7414_
timestamp 0
transform 1 0 7490 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7415_
timestamp 0
transform 1 0 7110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7416_
timestamp 0
transform -1 0 7150 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7417_
timestamp 0
transform 1 0 5930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7418_
timestamp 0
transform -1 0 5450 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7419_
timestamp 0
transform -1 0 6870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7420_
timestamp 0
transform 1 0 7430 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7421_
timestamp 0
transform 1 0 7030 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7422_
timestamp 0
transform 1 0 7650 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7423_
timestamp 0
transform 1 0 7570 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7424_
timestamp 0
transform -1 0 7670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7425_
timestamp 0
transform 1 0 7410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7426_
timestamp 0
transform -1 0 7550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7427_
timestamp 0
transform -1 0 7290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7428_
timestamp 0
transform 1 0 7030 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7429_
timestamp 0
transform -1 0 6810 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7430_
timestamp 0
transform -1 0 6730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7431_
timestamp 0
transform -1 0 6590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7432_
timestamp 0
transform -1 0 6650 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7433_
timestamp 0
transform 1 0 5590 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7434_
timestamp 0
transform 1 0 8210 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7435_
timestamp 0
transform 1 0 7470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7436_
timestamp 0
transform -1 0 7210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7437_
timestamp 0
transform -1 0 7350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7438_
timestamp 0
transform -1 0 7570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7439_
timestamp 0
transform 1 0 8030 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7440_
timestamp 0
transform 1 0 7170 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7441_
timestamp 0
transform -1 0 7710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7442_
timestamp 0
transform 1 0 7670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7443_
timestamp 0
transform 1 0 5250 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7444_
timestamp 0
transform -1 0 4610 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7445_
timestamp 0
transform 1 0 6530 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7446_
timestamp 0
transform 1 0 6370 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7447_
timestamp 0
transform -1 0 7690 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7448_
timestamp 0
transform 1 0 8230 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7449_
timestamp 0
transform 1 0 8770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7450_
timestamp 0
transform -1 0 8730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7451_
timestamp 0
transform -1 0 8070 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7452_
timestamp 0
transform -1 0 7570 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7453_
timestamp 0
transform 1 0 8190 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7454_
timestamp 0
transform 1 0 8310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7455_
timestamp 0
transform -1 0 10050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7456_
timestamp 0
transform -1 0 8610 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7457_
timestamp 0
transform -1 0 8510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7458_
timestamp 0
transform 1 0 10350 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7459_
timestamp 0
transform -1 0 5950 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7460_
timestamp 0
transform -1 0 6630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7461_
timestamp 0
transform -1 0 7710 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7462_
timestamp 0
transform -1 0 7830 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7463_
timestamp 0
transform 1 0 8050 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7464_
timestamp 0
transform 1 0 8410 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7465_
timestamp 0
transform 1 0 6870 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7466_
timestamp 0
transform 1 0 6730 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7467_
timestamp 0
transform 1 0 8490 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7468_
timestamp 0
transform -1 0 6810 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7469_
timestamp 0
transform -1 0 6930 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7470_
timestamp 0
transform -1 0 8230 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7471_
timestamp 0
transform 1 0 8350 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7472_
timestamp 0
transform -1 0 8710 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7473_
timestamp 0
transform -1 0 9190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7474_
timestamp 0
transform -1 0 8250 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7475_
timestamp 0
transform 1 0 8530 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7476_
timestamp 0
transform -1 0 9050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7477_
timestamp 0
transform 1 0 9570 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7478_
timestamp 0
transform -1 0 11090 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7479_
timestamp 0
transform 1 0 9410 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7480_
timestamp 0
transform -1 0 10950 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7481_
timestamp 0
transform -1 0 10150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7482_
timestamp 0
transform -1 0 9990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7483_
timestamp 0
transform -1 0 9410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7484_
timestamp 0
transform -1 0 8630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7485_
timestamp 0
transform -1 0 8750 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7486_
timestamp 0
transform 1 0 11170 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7487_
timestamp 0
transform -1 0 9270 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7488_
timestamp 0
transform -1 0 7650 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7489_
timestamp 0
transform -1 0 7770 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7490_
timestamp 0
transform -1 0 7850 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7491_
timestamp 0
transform 1 0 8330 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7492_
timestamp 0
transform 1 0 7810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7493_
timestamp 0
transform 1 0 7930 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7494_
timestamp 0
transform -1 0 7810 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7495_
timestamp 0
transform 1 0 8630 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7496_
timestamp 0
transform -1 0 9070 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7497_
timestamp 0
transform 1 0 9510 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7498_
timestamp 0
transform 1 0 8850 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7499_
timestamp 0
transform -1 0 8930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7500_
timestamp 0
transform 1 0 10150 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7501_
timestamp 0
transform -1 0 11650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7502_
timestamp 0
transform 1 0 10010 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7503_
timestamp 0
transform 1 0 11610 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7504_
timestamp 0
transform -1 0 11350 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7505_
timestamp 0
transform 1 0 11470 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7506_
timestamp 0
transform -1 0 10930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7507_
timestamp 0
transform -1 0 8870 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7508_
timestamp 0
transform 1 0 11750 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7509_
timestamp 0
transform 1 0 12210 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7510_
timestamp 0
transform -1 0 7710 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7511_
timestamp 0
transform -1 0 7850 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7512_
timestamp 0
transform 1 0 8610 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7513_
timestamp 0
transform 1 0 9030 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7514_
timestamp 0
transform -1 0 8090 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7515_
timestamp 0
transform -1 0 7950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7516_
timestamp 0
transform -1 0 8210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7517_
timestamp 0
transform 1 0 9170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7518_
timestamp 0
transform -1 0 9390 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7519_
timestamp 0
transform 1 0 10150 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7520_
timestamp 0
transform 1 0 9330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7521_
timestamp 0
transform 1 0 11350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7522_
timestamp 0
transform 1 0 12110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7523_
timestamp 0
transform 1 0 11490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7524_
timestamp 0
transform 1 0 12230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7525_
timestamp 0
transform 1 0 12430 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7526_
timestamp 0
transform -1 0 12330 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7527_
timestamp 0
transform 1 0 12570 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7528_
timestamp 0
transform 1 0 9770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7529_
timestamp 0
transform -1 0 11930 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7530_
timestamp 0
transform -1 0 7410 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7531_
timestamp 0
transform -1 0 7530 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7532_
timestamp 0
transform -1 0 7970 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7533_
timestamp 0
transform -1 0 8110 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7534_
timestamp 0
transform 1 0 8750 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7535_
timestamp 0
transform 1 0 8610 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7536_
timestamp 0
transform -1 0 10790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7537_
timestamp 0
transform 1 0 9110 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7538_
timestamp 0
transform 1 0 10810 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7539_
timestamp 0
transform 1 0 11670 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7540_
timestamp 0
transform -1 0 10710 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7541_
timestamp 0
transform -1 0 11150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7542_
timestamp 0
transform 1 0 11830 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7543_
timestamp 0
transform 1 0 11450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7544_
timestamp 0
transform 1 0 11290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7545_
timestamp 0
transform 1 0 12910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7546_
timestamp 0
transform 1 0 12630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7547_
timestamp 0
transform -1 0 12510 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7548_
timestamp 0
transform 1 0 12630 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7549_
timestamp 0
transform -1 0 12470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7550_
timestamp 0
transform 1 0 11130 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7551_
timestamp 0
transform -1 0 9690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7552_
timestamp 0
transform -1 0 11870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7553_
timestamp 0
transform 1 0 11090 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7554_
timestamp 0
transform -1 0 8390 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7555_
timestamp 0
transform 1 0 8770 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7556_
timestamp 0
transform -1 0 8790 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7557_
timestamp 0
transform -1 0 8910 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7558_
timestamp 0
transform 1 0 10410 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7559_
timestamp 0
transform 1 0 10950 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7560_
timestamp 0
transform 1 0 9270 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7561_
timestamp 0
transform 1 0 9130 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7562_
timestamp 0
transform 1 0 10130 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7563_
timestamp 0
transform -1 0 10290 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7564_
timestamp 0
transform 1 0 10990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7565_
timestamp 0
transform 1 0 13690 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7566_
timestamp 0
transform 1 0 10850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7567_
timestamp 0
transform 1 0 13550 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7568_
timestamp 0
transform -1 0 11730 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7569_
timestamp 0
transform -1 0 11750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7570_
timestamp 0
transform -1 0 11570 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7571_
timestamp 0
transform 1 0 10030 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7572_
timestamp 0
transform 1 0 9110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7573_
timestamp 0
transform -1 0 10530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7574_
timestamp 0
transform 1 0 8930 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7575_
timestamp 0
transform 1 0 9470 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7576_
timestamp 0
transform 1 0 9610 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7577_
timestamp 0
transform 1 0 10350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7578_
timestamp 0
transform 1 0 9510 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7579_
timestamp 0
transform -1 0 9630 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7580_
timestamp 0
transform 1 0 9770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7581_
timestamp 0
transform 1 0 12510 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7582_
timestamp 0
transform -1 0 12990 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7583_
timestamp 0
transform -1 0 12390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7584_
timestamp 0
transform -1 0 12010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7585_
timestamp 0
transform -1 0 12790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7586_
timestamp 0
transform -1 0 12650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7587_
timestamp 0
transform 1 0 12250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7588_
timestamp 0
transform -1 0 12150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7589_
timestamp 0
transform 1 0 12070 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7590_
timestamp 0
transform -1 0 11730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7591_
timestamp 0
transform 1 0 13950 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7592_
timestamp 0
transform 1 0 13810 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7593_
timestamp 0
transform 1 0 13410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7594_
timestamp 0
transform 1 0 13390 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7595_
timestamp 0
transform -1 0 11610 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7596_
timestamp 0
transform -1 0 10750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7597_
timestamp 0
transform 1 0 10230 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7598_
timestamp 0
transform 1 0 9230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7599_
timestamp 0
transform 1 0 10170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7600_
timestamp 0
transform 1 0 11870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7601_
timestamp 0
transform -1 0 9650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7602_
timestamp 0
transform 1 0 9070 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7603_
timestamp 0
transform 1 0 9190 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7604_
timestamp 0
transform 1 0 9310 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7605_
timestamp 0
transform 1 0 10410 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7606_
timestamp 0
transform 1 0 10010 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7607_
timestamp 0
transform 1 0 10210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7608_
timestamp 0
transform 1 0 10070 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7609_
timestamp 0
transform 1 0 10470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7610_
timestamp 0
transform 1 0 9910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7611_
timestamp 0
transform -1 0 10310 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7612_
timestamp 0
transform 1 0 10710 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7613_
timestamp 0
transform 1 0 11390 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7614_
timestamp 0
transform -1 0 11010 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7615_
timestamp 0
transform 1 0 11130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7616_
timestamp 0
transform -1 0 10910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7617_
timestamp 0
transform -1 0 10870 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7618_
timestamp 0
transform 1 0 10690 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7619_
timestamp 0
transform -1 0 12090 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7620_
timestamp 0
transform 1 0 12210 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7621_
timestamp 0
transform 1 0 12350 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7622_
timestamp 0
transform 1 0 11890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7623_
timestamp 0
transform -1 0 9750 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7624_
timestamp 0
transform 1 0 8890 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7625_
timestamp 0
transform 1 0 9310 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7626_
timestamp 0
transform -1 0 10630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7627_
timestamp 0
transform 1 0 10310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7628_
timestamp 0
transform 1 0 10550 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7629_
timestamp 0
transform 1 0 11530 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7630_
timestamp 0
transform 1 0 11750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7631_
timestamp 0
transform 1 0 10170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7632_
timestamp 0
transform 1 0 10710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7633_
timestamp 0
transform 1 0 11250 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7634_
timestamp 0
transform 1 0 11910 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7635_
timestamp 0
transform -1 0 10690 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7636_
timestamp 0
transform -1 0 11790 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7637_
timestamp 0
transform -1 0 11330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7638_
timestamp 0
transform 1 0 10570 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7639_
timestamp 0
transform -1 0 10270 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7640_
timestamp 0
transform 1 0 11610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7641_
timestamp 0
transform 1 0 11470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7642_
timestamp 0
transform 1 0 9170 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7643_
timestamp 0
transform 1 0 10050 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7644_
timestamp 0
transform -1 0 10030 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7645_
timestamp 0
transform -1 0 10870 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7646_
timestamp 0
transform 1 0 10970 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7647_
timestamp 0
transform 1 0 11050 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7648_
timestamp 0
transform 1 0 12830 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7649_
timestamp 0
transform -1 0 12730 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__7650_
timestamp 0
transform 1 0 11190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7651_
timestamp 0
transform -1 0 11030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7652_
timestamp 0
transform 1 0 11170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7653_
timestamp 0
transform -1 0 10410 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7654_
timestamp 0
transform 1 0 10130 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7655_
timestamp 0
transform 1 0 11510 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7656_
timestamp 0
transform -1 0 11630 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7657_
timestamp 0
transform 1 0 11470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7658_
timestamp 0
transform 1 0 11310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7659_
timestamp 0
transform 1 0 11370 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7660_
timestamp 0
transform 1 0 9450 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7661_
timestamp 0
transform -1 0 9430 0 1 730
box -6 -8 26 248
use FILL  FILL_1__7662_
timestamp 0
transform -1 0 9510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__7663_
timestamp 0
transform 1 0 9650 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7664_
timestamp 0
transform -1 0 10310 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7665_
timestamp 0
transform 1 0 10410 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7666_
timestamp 0
transform 1 0 10570 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__7667_
timestamp 0
transform -1 0 9610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7668_
timestamp 0
transform 1 0 9890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7669_
timestamp 0
transform -1 0 9770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7670_
timestamp 0
transform 1 0 10770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7671_
timestamp 0
transform -1 0 10750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7672_
timestamp 0
transform 1 0 10870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7673_
timestamp 0
transform -1 0 10570 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7674_
timestamp 0
transform 1 0 10170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7675_
timestamp 0
transform 1 0 9950 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7676_
timestamp 0
transform 1 0 11270 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7677_
timestamp 0
transform 1 0 11110 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7678_
timestamp 0
transform 1 0 10390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7679_
timestamp 0
transform 1 0 10250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7680_
timestamp 0
transform 1 0 10510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7681_
timestamp 0
transform 1 0 10650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__7682_
timestamp 0
transform -1 0 10590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7683_
timestamp 0
transform -1 0 10450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7684_
timestamp 0
transform -1 0 10110 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7685_
timestamp 0
transform 1 0 6830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7686_
timestamp 0
transform 1 0 6210 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7687_
timestamp 0
transform -1 0 6270 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7688_
timestamp 0
transform -1 0 6110 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7689_
timestamp 0
transform -1 0 6130 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7690_
timestamp 0
transform 1 0 5930 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7691_
timestamp 0
transform -1 0 5710 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7692_
timestamp 0
transform -1 0 5810 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7693_
timestamp 0
transform 1 0 5150 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__7694_
timestamp 0
transform -1 0 5490 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7695_
timestamp 0
transform 1 0 5070 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7696_
timestamp 0
transform -1 0 6070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7697_
timestamp 0
transform -1 0 6370 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7698_
timestamp 0
transform -1 0 6370 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7699_
timestamp 0
transform -1 0 6230 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7700_
timestamp 0
transform -1 0 5910 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7701_
timestamp 0
transform -1 0 5810 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__7702_
timestamp 0
transform -1 0 5770 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7703_
timestamp 0
transform -1 0 5670 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__7704_
timestamp 0
transform -1 0 5430 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__7705_
timestamp 0
transform 1 0 5530 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__7706_
timestamp 0
transform -1 0 5290 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__7707_
timestamp 0
transform -1 0 5030 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__7708_
timestamp 0
transform -1 0 6050 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7709_
timestamp 0
transform -1 0 5970 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__7710_
timestamp 0
transform 1 0 7210 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__7711_
timestamp 0
transform 1 0 7430 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__7712_
timestamp 0
transform 1 0 7270 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__7713_
timestamp 0
transform 1 0 7610 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__7714_
timestamp 0
transform -1 0 7490 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__7715_
timestamp 0
transform 1 0 7330 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__7716_
timestamp 0
transform -1 0 6830 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__7717_
timestamp 0
transform -1 0 6470 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__7718_
timestamp 0
transform -1 0 6790 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__7719_
timestamp 0
transform 1 0 6550 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__7720_
timestamp 0
transform 1 0 6270 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__7721_
timestamp 0
transform -1 0 5790 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__7722_
timestamp 0
transform -1 0 6930 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__7723_
timestamp 0
transform -1 0 6690 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__7724_
timestamp 0
transform -1 0 6690 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7725_
timestamp 0
transform -1 0 7690 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7726_
timestamp 0
transform -1 0 7550 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7727_
timestamp 0
transform 1 0 7050 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__7728_
timestamp 0
transform 1 0 7370 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__7729_
timestamp 0
transform -1 0 6530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7730_
timestamp 0
transform 1 0 6650 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7731_
timestamp 0
transform -1 0 6330 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7732_
timestamp 0
transform -1 0 6350 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__7733_
timestamp 0
transform 1 0 6410 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__7734_
timestamp 0
transform -1 0 6270 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__7735_
timestamp 0
transform 1 0 6130 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__7736_
timestamp 0
transform -1 0 6490 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__7737_
timestamp 0
transform -1 0 8090 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7738_
timestamp 0
transform -1 0 7350 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7739_
timestamp 0
transform 1 0 7170 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7740_
timestamp 0
transform 1 0 6770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7741_
timestamp 0
transform 1 0 7690 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7742_
timestamp 0
transform -1 0 7470 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7743_
timestamp 0
transform 1 0 7570 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7744_
timestamp 0
transform -1 0 6550 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7745_
timestamp 0
transform -1 0 6990 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__7746_
timestamp 0
transform 1 0 7110 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__7747_
timestamp 0
transform -1 0 6850 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__7748_
timestamp 0
transform 1 0 7590 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7749_
timestamp 0
transform -1 0 8130 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7750_
timestamp 0
transform 1 0 8170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7751_
timestamp 0
transform 1 0 8830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7752_
timestamp 0
transform -1 0 8710 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7753_
timestamp 0
transform 1 0 8270 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__7754_
timestamp 0
transform -1 0 8150 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7755_
timestamp 0
transform 1 0 8270 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7756_
timestamp 0
transform -1 0 8010 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7757_
timestamp 0
transform -1 0 7750 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7758_
timestamp 0
transform 1 0 7450 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7759_
timestamp 0
transform 1 0 7330 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7760_
timestamp 0
transform 1 0 7150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7761_
timestamp 0
transform 1 0 7290 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7762_
timestamp 0
transform -1 0 6430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7763_
timestamp 0
transform -1 0 7490 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7764_
timestamp 0
transform -1 0 7610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7765_
timestamp 0
transform 1 0 7830 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7766_
timestamp 0
transform 1 0 7850 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7767_
timestamp 0
transform 1 0 7710 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7768_
timestamp 0
transform 1 0 7870 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7769_
timestamp 0
transform 1 0 7950 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7770_
timestamp 0
transform 1 0 7830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7771_
timestamp 0
transform -1 0 7830 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7772_
timestamp 0
transform -1 0 7710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7773_
timestamp 0
transform 1 0 7610 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7774_
timestamp 0
transform -1 0 7490 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7775_
timestamp 0
transform 1 0 6910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7776_
timestamp 0
transform 1 0 7050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7777_
timestamp 0
transform 1 0 7330 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7778_
timestamp 0
transform -1 0 7230 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7779_
timestamp 0
transform 1 0 7070 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7780_
timestamp 0
transform -1 0 6950 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7781_
timestamp 0
transform 1 0 5530 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7782_
timestamp 0
transform 1 0 6630 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7783_
timestamp 0
transform 1 0 5130 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7784_
timestamp 0
transform -1 0 4890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7785_
timestamp 0
transform -1 0 4750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7786_
timestamp 0
transform 1 0 5010 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7787_
timestamp 0
transform -1 0 5150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7788_
timestamp 0
transform 1 0 5190 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7789_
timestamp 0
transform 1 0 5270 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7790_
timestamp 0
transform 1 0 5630 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7791_
timestamp 0
transform -1 0 6070 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7792_
timestamp 0
transform -1 0 5930 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7793_
timestamp 0
transform 1 0 5750 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7794_
timestamp 0
transform -1 0 8470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7795_
timestamp 0
transform -1 0 6990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7796_
timestamp 0
transform 1 0 7090 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7797_
timestamp 0
transform 1 0 7370 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7798_
timestamp 0
transform -1 0 7330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7799_
timestamp 0
transform -1 0 7230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7800_
timestamp 0
transform -1 0 7210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7801_
timestamp 0
transform -1 0 6490 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7802_
timestamp 0
transform 1 0 6770 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7803_
timestamp 0
transform -1 0 6910 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7804_
timestamp 0
transform -1 0 7210 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7805_
timestamp 0
transform -1 0 7070 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__7806_
timestamp 0
transform -1 0 7430 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7807_
timestamp 0
transform -1 0 7750 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7808_
timestamp 0
transform 1 0 8190 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7809_
timestamp 0
transform 1 0 8450 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7810_
timestamp 0
transform -1 0 7050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7811_
timestamp 0
transform -1 0 8030 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7812_
timestamp 0
transform 1 0 8150 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7813_
timestamp 0
transform 1 0 7870 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7814_
timestamp 0
transform -1 0 6550 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7815_
timestamp 0
transform -1 0 6390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7816_
timestamp 0
transform 1 0 6210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7817_
timestamp 0
transform 1 0 5930 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7818_
timestamp 0
transform 1 0 7450 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7819_
timestamp 0
transform -1 0 7750 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7820_
timestamp 0
transform 1 0 7610 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7821_
timestamp 0
transform -1 0 7330 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7822_
timestamp 0
transform 1 0 7050 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7823_
timestamp 0
transform 1 0 6930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7824_
timestamp 0
transform -1 0 6470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7825_
timestamp 0
transform -1 0 6330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7826_
timestamp 0
transform -1 0 6030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7827_
timestamp 0
transform 1 0 6150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7828_
timestamp 0
transform -1 0 5890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7829_
timestamp 0
transform 1 0 6050 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7830_
timestamp 0
transform 1 0 6310 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7831_
timestamp 0
transform -1 0 6190 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7832_
timestamp 0
transform 1 0 6750 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7833_
timestamp 0
transform 1 0 8370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7834_
timestamp 0
transform 1 0 6890 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__7835_
timestamp 0
transform -1 0 8630 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7836_
timestamp 0
transform -1 0 8750 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__7837_
timestamp 0
transform 1 0 6890 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7838_
timestamp 0
transform -1 0 6930 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7839_
timestamp 0
transform -1 0 10510 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7840_
timestamp 0
transform -1 0 7530 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__7841_
timestamp 0
transform 1 0 9590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7842_
timestamp 0
transform -1 0 9910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7843_
timestamp 0
transform -1 0 8810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7844_
timestamp 0
transform 1 0 9270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7845_
timestamp 0
transform 1 0 9130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7846_
timestamp 0
transform -1 0 6650 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7847_
timestamp 0
transform -1 0 10630 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7848_
timestamp 0
transform 1 0 10730 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7849_
timestamp 0
transform 1 0 9750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7850_
timestamp 0
transform 1 0 9570 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7851_
timestamp 0
transform -1 0 6150 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__7852_
timestamp 0
transform 1 0 11130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7853_
timestamp 0
transform 1 0 10970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__7854_
timestamp 0
transform 1 0 8910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7855_
timestamp 0
transform -1 0 8790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__7856_
timestamp 0
transform 1 0 8910 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7857_
timestamp 0
transform -1 0 9090 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7858_
timestamp 0
transform -1 0 8770 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7859_
timestamp 0
transform -1 0 8630 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7860_
timestamp 0
transform -1 0 8990 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7861_
timestamp 0
transform -1 0 9110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7862_
timestamp 0
transform 1 0 10230 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7863_
timestamp 0
transform 1 0 10070 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__7864_
timestamp 0
transform -1 0 7230 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7865_
timestamp 0
transform -1 0 7070 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__7866_
timestamp 0
transform 1 0 7270 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7867_
timestamp 0
transform 1 0 7130 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7868_
timestamp 0
transform -1 0 6790 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7869_
timestamp 0
transform -1 0 6910 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7870_
timestamp 0
transform -1 0 7050 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7871_
timestamp 0
transform -1 0 6970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7872_
timestamp 0
transform -1 0 7930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7873_
timestamp 0
transform 1 0 7530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7874_
timestamp 0
transform 1 0 6490 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7875_
timestamp 0
transform -1 0 6630 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7876_
timestamp 0
transform 1 0 6670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7877_
timestamp 0
transform -1 0 6810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7878_
timestamp 0
transform -1 0 6270 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7879_
timestamp 0
transform 1 0 6110 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__7880_
timestamp 0
transform -1 0 6070 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7881_
timestamp 0
transform -1 0 6210 0 1 250
box -6 -8 26 248
use FILL  FILL_1__7882_
timestamp 0
transform -1 0 7170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7883_
timestamp 0
transform 1 0 7010 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7884_
timestamp 0
transform -1 0 7210 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7885_
timestamp 0
transform -1 0 7370 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7886_
timestamp 0
transform -1 0 8090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7887_
timestamp 0
transform 1 0 8190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__7888_
timestamp 0
transform -1 0 7330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7889_
timestamp 0
transform -1 0 7450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__7890_
timestamp 0
transform 1 0 7330 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7891_
timestamp 0
transform 1 0 7170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__7892_
timestamp 0
transform 1 0 8490 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7893_
timestamp 0
transform 1 0 8350 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__7894_
timestamp 0
transform 1 0 8330 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7895_
timestamp 0
transform 1 0 8050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7896_
timestamp 0
transform -1 0 8210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7897_
timestamp 0
transform -1 0 6950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7898_
timestamp 0
transform 1 0 7910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7899_
timestamp 0
transform 1 0 7510 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__7900_
timestamp 0
transform -1 0 7950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7901_
timestamp 0
transform -1 0 8070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7902_
timestamp 0
transform 1 0 5050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7903_
timestamp 0
transform -1 0 4910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7904_
timestamp 0
transform -1 0 7870 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7905_
timestamp 0
transform -1 0 7990 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7906_
timestamp 0
transform 1 0 8830 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7907_
timestamp 0
transform 1 0 8470 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__7908_
timestamp 0
transform -1 0 8290 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7909_
timestamp 0
transform -1 0 7810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__7910_
timestamp 0
transform 1 0 6770 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7911_
timestamp 0
transform -1 0 6930 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__7912_
timestamp 0
transform 1 0 7050 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7913_
timestamp 0
transform 1 0 6770 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7914_
timestamp 0
transform 1 0 6930 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__7915_
timestamp 0
transform 1 0 6150 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__7996_
timestamp 0
transform -1 0 6230 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__7997_
timestamp 0
transform -1 0 5190 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__7998_
timestamp 0
transform -1 0 4930 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__7999_
timestamp 0
transform 1 0 4990 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8000_
timestamp 0
transform 1 0 4330 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8001_
timestamp 0
transform 1 0 4210 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8002_
timestamp 0
transform -1 0 4490 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8003_
timestamp 0
transform -1 0 4650 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8004_
timestamp 0
transform -1 0 4510 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8005_
timestamp 0
transform -1 0 4350 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8006_
timestamp 0
transform -1 0 5290 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8007_
timestamp 0
transform 1 0 4470 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8008_
timestamp 0
transform 1 0 5050 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8009_
timestamp 0
transform 1 0 4310 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8010_
timestamp 0
transform -1 0 3770 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8011_
timestamp 0
transform -1 0 5450 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__8012_
timestamp 0
transform -1 0 4010 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__8013_
timestamp 0
transform -1 0 4170 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__8014_
timestamp 0
transform 1 0 6550 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8015_
timestamp 0
transform -1 0 5030 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8016_
timestamp 0
transform 1 0 4870 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8017_
timestamp 0
transform 1 0 4850 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8018_
timestamp 0
transform -1 0 4890 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8019_
timestamp 0
transform -1 0 4490 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8020_
timestamp 0
transform 1 0 3290 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8021_
timestamp 0
transform 1 0 4370 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8022_
timestamp 0
transform -1 0 4230 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8023_
timestamp 0
transform 1 0 3330 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8024_
timestamp 0
transform 1 0 2970 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8025_
timestamp 0
transform -1 0 3410 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8026_
timestamp 0
transform -1 0 3550 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8027_
timestamp 0
transform -1 0 4230 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8028_
timestamp 0
transform -1 0 3710 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8029_
timestamp 0
transform 1 0 3350 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8030_
timestamp 0
transform 1 0 3790 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8031_
timestamp 0
transform -1 0 3650 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8032_
timestamp 0
transform 1 0 2870 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8033_
timestamp 0
transform 1 0 3110 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8034_
timestamp 0
transform -1 0 3270 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8035_
timestamp 0
transform -1 0 3370 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8036_
timestamp 0
transform -1 0 4350 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8037_
timestamp 0
transform -1 0 3510 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8038_
timestamp 0
transform 1 0 3070 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8039_
timestamp 0
transform 1 0 4090 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8040_
timestamp 0
transform 1 0 3850 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8041_
timestamp 0
transform 1 0 4430 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8042_
timestamp 0
transform 1 0 4670 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8043_
timestamp 0
transform 1 0 4510 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8044_
timestamp 0
transform -1 0 3730 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8045_
timestamp 0
transform 1 0 3910 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8046_
timestamp 0
transform -1 0 3610 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8047_
timestamp 0
transform 1 0 2770 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8048_
timestamp 0
transform -1 0 3550 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8049_
timestamp 0
transform 1 0 3930 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8050_
timestamp 0
transform 1 0 4550 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8051_
timestamp 0
transform 1 0 3610 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8052_
timestamp 0
transform 1 0 3050 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8053_
timestamp 0
transform 1 0 2890 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8054_
timestamp 0
transform 1 0 4610 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8055_
timestamp 0
transform -1 0 5390 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8056_
timestamp 0
transform -1 0 1290 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8057_
timestamp 0
transform 1 0 1550 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8058_
timestamp 0
transform 1 0 2370 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8059_
timestamp 0
transform 1 0 2630 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8060_
timestamp 0
transform 1 0 2470 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8061_
timestamp 0
transform 1 0 3490 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8062_
timestamp 0
transform -1 0 3930 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8063_
timestamp 0
transform 1 0 3770 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8064_
timestamp 0
transform 1 0 3590 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8065_
timestamp 0
transform 1 0 4150 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8066_
timestamp 0
transform 1 0 3790 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8067_
timestamp 0
transform -1 0 4010 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8068_
timestamp 0
transform -1 0 2830 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8069_
timestamp 0
transform -1 0 2930 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8070_
timestamp 0
transform -1 0 3070 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8071_
timestamp 0
transform 1 0 3830 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8072_
timestamp 0
transform 1 0 3790 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8073_
timestamp 0
transform -1 0 5130 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8074_
timestamp 0
transform 1 0 5230 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8075_
timestamp 0
transform -1 0 5130 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8076_
timestamp 0
transform 1 0 5550 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8077_
timestamp 0
transform -1 0 4490 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8078_
timestamp 0
transform -1 0 4390 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8079_
timestamp 0
transform -1 0 4970 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8080_
timestamp 0
transform 1 0 4710 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8081_
timestamp 0
transform 1 0 6830 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8082_
timestamp 0
transform 1 0 4870 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8083_
timestamp 0
transform 1 0 5230 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8084_
timestamp 0
transform -1 0 2870 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8085_
timestamp 0
transform -1 0 3050 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8086_
timestamp 0
transform -1 0 2610 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8087_
timestamp 0
transform -1 0 3710 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8088_
timestamp 0
transform 1 0 3650 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8089_
timestamp 0
transform -1 0 3530 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8090_
timestamp 0
transform 1 0 3250 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8091_
timestamp 0
transform 1 0 3130 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8092_
timestamp 0
transform 1 0 3290 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8093_
timestamp 0
transform -1 0 3350 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8094_
timestamp 0
transform -1 0 5750 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8095_
timestamp 0
transform -1 0 50 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8096_
timestamp 0
transform -1 0 2750 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8097_
timestamp 0
transform -1 0 2490 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8098_
timestamp 0
transform -1 0 2710 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8099_
timestamp 0
transform 1 0 3110 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8100_
timestamp 0
transform 1 0 3350 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8101_
timestamp 0
transform 1 0 3210 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8102_
timestamp 0
transform 1 0 3010 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8103_
timestamp 0
transform -1 0 3210 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8104_
timestamp 0
transform 1 0 3330 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8105_
timestamp 0
transform 1 0 3170 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8106_
timestamp 0
transform -1 0 2650 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8107_
timestamp 0
transform -1 0 2230 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8108_
timestamp 0
transform -1 0 2370 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8109_
timestamp 0
transform 1 0 3450 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8110_
timestamp 0
transform -1 0 3630 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8111_
timestamp 0
transform 1 0 4770 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8112_
timestamp 0
transform -1 0 2130 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8113_
timestamp 0
transform -1 0 2330 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8114_
timestamp 0
transform 1 0 2130 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8115_
timestamp 0
transform -1 0 3510 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8116_
timestamp 0
transform 1 0 3170 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8117_
timestamp 0
transform -1 0 3330 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8118_
timestamp 0
transform 1 0 3770 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8119_
timestamp 0
transform 1 0 4810 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8120_
timestamp 0
transform 1 0 5070 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8121_
timestamp 0
transform 1 0 5350 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8122_
timestamp 0
transform -1 0 4930 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8123_
timestamp 0
transform -1 0 4990 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8124_
timestamp 0
transform -1 0 4810 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8125_
timestamp 0
transform -1 0 4670 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8126_
timestamp 0
transform -1 0 4510 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8127_
timestamp 0
transform 1 0 4730 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8128_
timestamp 0
transform 1 0 7030 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__8129_
timestamp 0
transform 1 0 7190 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__8130_
timestamp 0
transform 1 0 7050 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__8131_
timestamp 0
transform 1 0 4490 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8132_
timestamp 0
transform 1 0 5210 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8133_
timestamp 0
transform -1 0 1910 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8134_
timestamp 0
transform -1 0 1970 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8135_
timestamp 0
transform 1 0 4070 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8136_
timestamp 0
transform -1 0 4070 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8137_
timestamp 0
transform 1 0 4190 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8138_
timestamp 0
transform 1 0 4350 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8139_
timestamp 0
transform -1 0 4690 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8140_
timestamp 0
transform 1 0 4650 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8141_
timestamp 0
transform -1 0 4270 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8142_
timestamp 0
transform 1 0 4510 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8143_
timestamp 0
transform 1 0 4370 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8144_
timestamp 0
transform 1 0 4950 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8145_
timestamp 0
transform -1 0 4810 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8146_
timestamp 0
transform -1 0 4790 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8147_
timestamp 0
transform 1 0 5030 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8148_
timestamp 0
transform 1 0 5270 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8149_
timestamp 0
transform -1 0 5190 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8150_
timestamp 0
transform 1 0 4870 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8151_
timestamp 0
transform -1 0 5110 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8152_
timestamp 0
transform -1 0 1090 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8153_
timestamp 0
transform 1 0 3910 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8154_
timestamp 0
transform 1 0 4350 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8155_
timestamp 0
transform 1 0 3550 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8156_
timestamp 0
transform -1 0 4270 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8157_
timestamp 0
transform -1 0 4630 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8158_
timestamp 0
transform 1 0 2950 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8159_
timestamp 0
transform -1 0 2570 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8160_
timestamp 0
transform -1 0 4530 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8161_
timestamp 0
transform -1 0 1890 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8162_
timestamp 0
transform -1 0 1550 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8163_
timestamp 0
transform -1 0 1590 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8164_
timestamp 0
transform 1 0 1850 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8165_
timestamp 0
transform 1 0 1550 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8166_
timestamp 0
transform -1 0 1370 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8167_
timestamp 0
transform 1 0 5950 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8168_
timestamp 0
transform -1 0 2870 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8169_
timestamp 0
transform 1 0 1570 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8170_
timestamp 0
transform 1 0 1410 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8171_
timestamp 0
transform 1 0 750 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8172_
timestamp 0
transform 1 0 990 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8173_
timestamp 0
transform 1 0 850 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8174_
timestamp 0
transform 1 0 1970 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8175_
timestamp 0
transform 1 0 2130 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8176_
timestamp 0
transform 1 0 2350 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__8177_
timestamp 0
transform -1 0 2450 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8178_
timestamp 0
transform 1 0 2650 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8179_
timestamp 0
transform -1 0 2810 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8180_
timestamp 0
transform -1 0 3410 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8181_
timestamp 0
transform -1 0 2290 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8182_
timestamp 0
transform 1 0 1730 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__8183_
timestamp 0
transform -1 0 710 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8184_
timestamp 0
transform -1 0 430 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8185_
timestamp 0
transform -1 0 570 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8186_
timestamp 0
transform -1 0 1730 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8187_
timestamp 0
transform 1 0 690 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8188_
timestamp 0
transform 1 0 1650 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8189_
timestamp 0
transform -1 0 710 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8190_
timestamp 0
transform 1 0 730 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8191_
timestamp 0
transform 1 0 790 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8192_
timestamp 0
transform -1 0 290 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__8193_
timestamp 0
transform -1 0 850 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8194_
timestamp 0
transform -1 0 630 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8195_
timestamp 0
transform 1 0 710 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__8196_
timestamp 0
transform 1 0 550 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__8197_
timestamp 0
transform 1 0 410 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__8198_
timestamp 0
transform 1 0 690 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__8199_
timestamp 0
transform 1 0 990 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__8200_
timestamp 0
transform 1 0 1110 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8201_
timestamp 0
transform 1 0 1270 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8202_
timestamp 0
transform -1 0 2810 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8203_
timestamp 0
transform -1 0 970 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8204_
timestamp 0
transform -1 0 1410 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__8205_
timestamp 0
transform -1 0 470 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8206_
timestamp 0
transform -1 0 790 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8207_
timestamp 0
transform 1 0 1010 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8208_
timestamp 0
transform -1 0 770 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8209_
timestamp 0
transform 1 0 1050 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8210_
timestamp 0
transform 1 0 530 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8211_
timestamp 0
transform -1 0 50 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8212_
timestamp 0
transform -1 0 670 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8213_
timestamp 0
transform -1 0 510 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8214_
timestamp 0
transform -1 0 370 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8215_
timestamp 0
transform 1 0 30 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8216_
timestamp 0
transform 1 0 30 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__8217_
timestamp 0
transform 1 0 170 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__8218_
timestamp 0
transform 1 0 170 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8219_
timestamp 0
transform 1 0 1110 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8220_
timestamp 0
transform -1 0 990 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8221_
timestamp 0
transform 1 0 1270 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8222_
timestamp 0
transform -1 0 2490 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8223_
timestamp 0
transform -1 0 2150 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8224_
timestamp 0
transform 1 0 490 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8225_
timestamp 0
transform 1 0 590 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8226_
timestamp 0
transform -1 0 610 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8227_
timestamp 0
transform 1 0 410 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8228_
timestamp 0
transform -1 0 290 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8229_
timestamp 0
transform -1 0 50 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8230_
timestamp 0
transform 1 0 150 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8231_
timestamp 0
transform -1 0 310 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8232_
timestamp 0
transform 1 0 250 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8233_
timestamp 0
transform 1 0 350 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8234_
timestamp 0
transform -1 0 50 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8235_
timestamp 0
transform 1 0 370 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8236_
timestamp 0
transform 1 0 490 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8237_
timestamp 0
transform 1 0 710 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8238_
timestamp 0
transform -1 0 570 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__8239_
timestamp 0
transform -1 0 450 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__8240_
timestamp 0
transform -1 0 670 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8241_
timestamp 0
transform 1 0 510 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8242_
timestamp 0
transform 1 0 1130 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8243_
timestamp 0
transform 1 0 1190 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8244_
timestamp 0
transform -1 0 1990 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8245_
timestamp 0
transform -1 0 2810 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8246_
timestamp 0
transform -1 0 210 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8247_
timestamp 0
transform -1 0 870 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__8248_
timestamp 0
transform 1 0 190 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8249_
timestamp 0
transform -1 0 310 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__8250_
timestamp 0
transform -1 0 370 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8251_
timestamp 0
transform 1 0 430 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8252_
timestamp 0
transform -1 0 190 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8253_
timestamp 0
transform -1 0 210 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8254_
timestamp 0
transform 1 0 670 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8255_
timestamp 0
transform -1 0 790 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8256_
timestamp 0
transform 1 0 890 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8257_
timestamp 0
transform -1 0 850 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8258_
timestamp 0
transform 1 0 370 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8259_
timestamp 0
transform -1 0 50 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8260_
timestamp 0
transform 1 0 150 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8261_
timestamp 0
transform 1 0 130 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8262_
timestamp 0
transform 1 0 510 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8263_
timestamp 0
transform 1 0 30 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8264_
timestamp 0
transform -1 0 270 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8265_
timestamp 0
transform 1 0 170 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8266_
timestamp 0
transform 1 0 790 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8267_
timestamp 0
transform -1 0 810 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8268_
timestamp 0
transform -1 0 690 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8269_
timestamp 0
transform -1 0 850 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8270_
timestamp 0
transform 1 0 910 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8271_
timestamp 0
transform -1 0 2510 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8272_
timestamp 0
transform -1 0 2170 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8273_
timestamp 0
transform 1 0 990 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8274_
timestamp 0
transform -1 0 2650 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8275_
timestamp 0
transform -1 0 2290 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8276_
timestamp 0
transform 1 0 910 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8277_
timestamp 0
transform -1 0 1010 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8278_
timestamp 0
transform 1 0 1050 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8279_
timestamp 0
transform -1 0 390 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8280_
timestamp 0
transform -1 0 50 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8281_
timestamp 0
transform -1 0 550 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8282_
timestamp 0
transform 1 0 170 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8283_
timestamp 0
transform -1 0 50 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8284_
timestamp 0
transform -1 0 50 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8285_
timestamp 0
transform -1 0 50 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8286_
timestamp 0
transform -1 0 230 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8287_
timestamp 0
transform 1 0 150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8288_
timestamp 0
transform 1 0 310 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8289_
timestamp 0
transform 1 0 470 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8290_
timestamp 0
transform 1 0 490 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8291_
timestamp 0
transform 1 0 1030 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8292_
timestamp 0
transform 1 0 1390 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8293_
timestamp 0
transform 1 0 1530 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8294_
timestamp 0
transform -1 0 2010 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8295_
timestamp 0
transform 1 0 310 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8296_
timestamp 0
transform 1 0 330 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8297_
timestamp 0
transform 1 0 570 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8298_
timestamp 0
transform -1 0 650 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8299_
timestamp 0
transform -1 0 510 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8300_
timestamp 0
transform 1 0 610 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8301_
timestamp 0
transform 1 0 630 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8302_
timestamp 0
transform -1 0 1010 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8303_
timestamp 0
transform 1 0 150 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8304_
timestamp 0
transform -1 0 190 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8305_
timestamp 0
transform 1 0 730 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8306_
timestamp 0
transform 1 0 30 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8307_
timestamp 0
transform -1 0 50 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8308_
timestamp 0
transform -1 0 290 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8309_
timestamp 0
transform -1 0 450 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8310_
timestamp 0
transform 1 0 130 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8311_
timestamp 0
transform 1 0 290 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8312_
timestamp 0
transform 1 0 430 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8313_
timestamp 0
transform 1 0 590 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8314_
timestamp 0
transform 1 0 1130 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8315_
timestamp 0
transform 1 0 1270 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8316_
timestamp 0
transform 1 0 1430 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8317_
timestamp 0
transform -1 0 3210 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8318_
timestamp 0
transform 1 0 450 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8319_
timestamp 0
transform 1 0 430 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8320_
timestamp 0
transform 1 0 470 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8321_
timestamp 0
transform -1 0 190 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8322_
timestamp 0
transform 1 0 310 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8323_
timestamp 0
transform -1 0 170 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8324_
timestamp 0
transform -1 0 590 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8325_
timestamp 0
transform 1 0 270 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8326_
timestamp 0
transform -1 0 430 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8327_
timestamp 0
transform -1 0 50 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8328_
timestamp 0
transform -1 0 190 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8329_
timestamp 0
transform -1 0 50 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8330_
timestamp 0
transform -1 0 330 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8331_
timestamp 0
transform -1 0 550 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8332_
timestamp 0
transform 1 0 570 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8333_
timestamp 0
transform 1 0 710 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8334_
timestamp 0
transform 1 0 710 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8335_
timestamp 0
transform 1 0 870 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8336_
timestamp 0
transform 1 0 670 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8337_
timestamp 0
transform 1 0 730 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8338_
timestamp 0
transform 1 0 870 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8339_
timestamp 0
transform 1 0 970 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8340_
timestamp 0
transform 1 0 1110 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8341_
timestamp 0
transform -1 0 2890 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8342_
timestamp 0
transform 1 0 3510 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8343_
timestamp 0
transform -1 0 570 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8344_
timestamp 0
transform -1 0 690 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8345_
timestamp 0
transform 1 0 790 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8346_
timestamp 0
transform 1 0 530 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8347_
timestamp 0
transform -1 0 430 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8348_
timestamp 0
transform -1 0 170 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8349_
timestamp 0
transform -1 0 190 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8350_
timestamp 0
transform -1 0 50 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8351_
timestamp 0
transform 1 0 290 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8352_
timestamp 0
transform -1 0 690 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8353_
timestamp 0
transform 1 0 770 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8354_
timestamp 0
transform -1 0 850 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8355_
timestamp 0
transform 1 0 1250 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8356_
timestamp 0
transform 1 0 1410 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8357_
timestamp 0
transform -1 0 3170 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8358_
timestamp 0
transform 1 0 3370 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8359_
timestamp 0
transform 1 0 4570 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8360_
timestamp 0
transform -1 0 4310 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8361_
timestamp 0
transform -1 0 4450 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8362_
timestamp 0
transform 1 0 4110 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8363_
timestamp 0
transform 1 0 5830 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8364_
timestamp 0
transform -1 0 5230 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8365_
timestamp 0
transform 1 0 5690 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8366_
timestamp 0
transform -1 0 3990 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8367_
timestamp 0
transform 1 0 750 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8368_
timestamp 0
transform 1 0 610 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8369_
timestamp 0
transform 1 0 1250 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__8370_
timestamp 0
transform -1 0 1130 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__8371_
timestamp 0
transform 1 0 1270 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8372_
timestamp 0
transform -1 0 1730 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8373_
timestamp 0
transform -1 0 2730 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8374_
timestamp 0
transform -1 0 2690 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8375_
timestamp 0
transform 1 0 1150 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8376_
timestamp 0
transform -1 0 910 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8377_
timestamp 0
transform -1 0 1030 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8378_
timestamp 0
transform 1 0 2010 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8379_
timestamp 0
transform 1 0 2850 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8380_
timestamp 0
transform 1 0 2950 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8381_
timestamp 0
transform -1 0 2770 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8382_
timestamp 0
transform -1 0 2750 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8383_
timestamp 0
transform 1 0 1830 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__8384_
timestamp 0
transform -1 0 1830 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8385_
timestamp 0
transform -1 0 5370 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8386_
timestamp 0
transform -1 0 5490 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8387_
timestamp 0
transform 1 0 2950 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8388_
timestamp 0
transform 1 0 1890 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8389_
timestamp 0
transform -1 0 310 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8390_
timestamp 0
transform -1 0 410 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8391_
timestamp 0
transform 1 0 830 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8392_
timestamp 0
transform -1 0 910 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8393_
timestamp 0
transform -1 0 1030 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8394_
timestamp 0
transform -1 0 1110 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8395_
timestamp 0
transform -1 0 970 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8396_
timestamp 0
transform 1 0 1730 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8397_
timestamp 0
transform 1 0 2490 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8398_
timestamp 0
transform 1 0 1210 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8399_
timestamp 0
transform -1 0 1810 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8400_
timestamp 0
transform -1 0 2610 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8401_
timestamp 0
transform 1 0 2530 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8402_
timestamp 0
transform 1 0 2630 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8403_
timestamp 0
transform -1 0 2390 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8404_
timestamp 0
transform -1 0 2510 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8405_
timestamp 0
transform -1 0 2390 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8406_
timestamp 0
transform 1 0 2510 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8407_
timestamp 0
transform 1 0 2650 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8408_
timestamp 0
transform -1 0 2610 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8409_
timestamp 0
transform -1 0 3570 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8410_
timestamp 0
transform -1 0 2350 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8411_
timestamp 0
transform 1 0 2310 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8412_
timestamp 0
transform -1 0 1010 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8413_
timestamp 0
transform 1 0 1130 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8414_
timestamp 0
transform -1 0 1290 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8415_
timestamp 0
transform -1 0 1410 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8416_
timestamp 0
transform 1 0 4050 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8417_
timestamp 0
transform 1 0 1430 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8418_
timestamp 0
transform -1 0 1570 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8419_
timestamp 0
transform 1 0 1610 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8420_
timestamp 0
transform 1 0 2030 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8421_
timestamp 0
transform 1 0 2290 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8422_
timestamp 0
transform 1 0 2150 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8423_
timestamp 0
transform -1 0 2590 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8424_
timestamp 0
transform -1 0 2310 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8425_
timestamp 0
transform 1 0 1970 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8426_
timestamp 0
transform 1 0 2450 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8427_
timestamp 0
transform -1 0 2110 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8428_
timestamp 0
transform 1 0 2230 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8429_
timestamp 0
transform -1 0 2070 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8430_
timestamp 0
transform 1 0 2190 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8431_
timestamp 0
transform 1 0 3390 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8432_
timestamp 0
transform -1 0 2090 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8433_
timestamp 0
transform -1 0 1750 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8434_
timestamp 0
transform -1 0 870 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8435_
timestamp 0
transform -1 0 930 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8436_
timestamp 0
transform 1 0 890 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8437_
timestamp 0
transform -1 0 1410 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8438_
timestamp 0
transform -1 0 2850 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8439_
timestamp 0
transform 1 0 1670 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8440_
timestamp 0
transform -1 0 1830 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8441_
timestamp 0
transform -1 0 1950 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8442_
timestamp 0
transform -1 0 2170 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8443_
timestamp 0
transform 1 0 2230 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8444_
timestamp 0
transform 1 0 2090 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8445_
timestamp 0
transform 1 0 2530 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8446_
timestamp 0
transform -1 0 2590 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8447_
timestamp 0
transform -1 0 2410 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8448_
timestamp 0
transform -1 0 2450 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8449_
timestamp 0
transform 1 0 1830 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8450_
timestamp 0
transform 1 0 1830 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8451_
timestamp 0
transform 1 0 1970 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8452_
timestamp 0
transform -1 0 2390 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8453_
timestamp 0
transform 1 0 2670 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8454_
timestamp 0
transform -1 0 1030 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8455_
timestamp 0
transform 1 0 1130 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8456_
timestamp 0
transform -1 0 1450 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8457_
timestamp 0
transform -1 0 1570 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8458_
timestamp 0
transform 1 0 1690 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8459_
timestamp 0
transform 1 0 1570 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8460_
timestamp 0
transform 1 0 2170 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8461_
timestamp 0
transform -1 0 2450 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8462_
timestamp 0
transform -1 0 1870 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8463_
timestamp 0
transform 1 0 2590 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8464_
timestamp 0
transform 1 0 2010 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8465_
timestamp 0
transform 1 0 2430 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8466_
timestamp 0
transform -1 0 3130 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8467_
timestamp 0
transform 1 0 2130 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8468_
timestamp 0
transform -1 0 2310 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8469_
timestamp 0
transform 1 0 2970 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8470_
timestamp 0
transform 1 0 3410 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8471_
timestamp 0
transform 1 0 4230 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8472_
timestamp 0
transform -1 0 4110 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8473_
timestamp 0
transform 1 0 4170 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8474_
timestamp 0
transform -1 0 4270 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8475_
timestamp 0
transform 1 0 4530 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8476_
timestamp 0
transform -1 0 3970 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8477_
timestamp 0
transform -1 0 2310 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8478_
timestamp 0
transform -1 0 1210 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8479_
timestamp 0
transform 1 0 1270 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8480_
timestamp 0
transform -1 0 1310 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8481_
timestamp 0
transform -1 0 1430 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8482_
timestamp 0
transform 1 0 1930 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8483_
timestamp 0
transform 1 0 2430 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8484_
timestamp 0
transform 1 0 1890 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8485_
timestamp 0
transform -1 0 1770 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8486_
timestamp 0
transform -1 0 1570 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8487_
timestamp 0
transform -1 0 1450 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8488_
timestamp 0
transform 1 0 2710 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8489_
timestamp 0
transform 1 0 3430 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8490_
timestamp 0
transform -1 0 2590 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8491_
timestamp 0
transform 1 0 3550 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8492_
timestamp 0
transform -1 0 3990 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8493_
timestamp 0
transform 1 0 4090 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8494_
timestamp 0
transform 1 0 4250 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8495_
timestamp 0
transform -1 0 4410 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8496_
timestamp 0
transform -1 0 4230 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8497_
timestamp 0
transform -1 0 2050 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8498_
timestamp 0
transform 1 0 1310 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8499_
timestamp 0
transform -1 0 1450 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8500_
timestamp 0
transform -1 0 1490 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8501_
timestamp 0
transform 1 0 2210 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8502_
timestamp 0
transform -1 0 1730 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8503_
timestamp 0
transform -1 0 1570 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8504_
timestamp 0
transform 1 0 2070 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8505_
timestamp 0
transform -1 0 2390 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8506_
timestamp 0
transform -1 0 2670 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8507_
timestamp 0
transform 1 0 2510 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8508_
timestamp 0
transform -1 0 3050 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8509_
timestamp 0
transform 1 0 2830 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8510_
timestamp 0
transform -1 0 2870 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8511_
timestamp 0
transform -1 0 3850 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8512_
timestamp 0
transform 1 0 3690 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8513_
timestamp 0
transform 1 0 3430 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8514_
timestamp 0
transform 1 0 3170 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8515_
timestamp 0
transform 1 0 3250 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8516_
timestamp 0
transform -1 0 3310 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8517_
timestamp 0
transform 1 0 2990 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8518_
timestamp 0
transform -1 0 3170 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8519_
timestamp 0
transform 1 0 3310 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8520_
timestamp 0
transform 1 0 3550 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8521_
timestamp 0
transform -1 0 3950 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8522_
timestamp 0
transform -1 0 4070 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8523_
timestamp 0
transform -1 0 4390 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8524_
timestamp 0
transform -1 0 2770 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8525_
timestamp 0
transform 1 0 1810 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8526_
timestamp 0
transform -1 0 1110 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8527_
timestamp 0
transform 1 0 1210 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8528_
timestamp 0
transform 1 0 1170 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8529_
timestamp 0
transform 1 0 1210 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8530_
timestamp 0
transform 1 0 1110 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8531_
timestamp 0
transform -1 0 1950 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8532_
timestamp 0
transform -1 0 1510 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8533_
timestamp 0
transform 1 0 1630 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8534_
timestamp 0
transform 1 0 1770 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8535_
timestamp 0
transform 1 0 1370 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8536_
timestamp 0
transform -1 0 1950 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8537_
timestamp 0
transform -1 0 2110 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8538_
timestamp 0
transform -1 0 2890 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8539_
timestamp 0
transform 1 0 3010 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8540_
timestamp 0
transform 1 0 3710 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8541_
timestamp 0
transform 1 0 3810 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8542_
timestamp 0
transform -1 0 3990 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8543_
timestamp 0
transform -1 0 2230 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__8544_
timestamp 0
transform -1 0 2930 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8545_
timestamp 0
transform -1 0 2790 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8546_
timestamp 0
transform -1 0 2150 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8547_
timestamp 0
transform 1 0 1670 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8548_
timestamp 0
transform -1 0 1630 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8549_
timestamp 0
transform -1 0 1490 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8550_
timestamp 0
transform -1 0 1650 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8551_
timestamp 0
transform 1 0 1690 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8552_
timestamp 0
transform 1 0 1410 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__8553_
timestamp 0
transform 1 0 1850 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8554_
timestamp 0
transform 1 0 1990 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8555_
timestamp 0
transform 1 0 1730 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8556_
timestamp 0
transform 1 0 1730 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8557_
timestamp 0
transform 1 0 1850 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8558_
timestamp 0
transform 1 0 2010 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8559_
timestamp 0
transform 1 0 2170 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8560_
timestamp 0
transform 1 0 1850 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8561_
timestamp 0
transform 1 0 2530 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8562_
timestamp 0
transform -1 0 2690 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8563_
timestamp 0
transform 1 0 3010 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8564_
timestamp 0
transform 1 0 2410 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8565_
timestamp 0
transform 1 0 2270 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8566_
timestamp 0
transform -1 0 1510 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8567_
timestamp 0
transform 1 0 1690 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8568_
timestamp 0
transform -1 0 1750 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8569_
timestamp 0
transform -1 0 1830 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8570_
timestamp 0
transform 1 0 1930 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8571_
timestamp 0
transform 1 0 2230 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8572_
timestamp 0
transform 1 0 2090 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8573_
timestamp 0
transform -1 0 1730 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8574_
timestamp 0
transform -1 0 2210 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8575_
timestamp 0
transform 1 0 2330 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8576_
timestamp 0
transform 1 0 2470 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8577_
timestamp 0
transform 1 0 2610 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8578_
timestamp 0
transform -1 0 4010 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8579_
timestamp 0
transform -1 0 2090 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8580_
timestamp 0
transform -1 0 1810 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8581_
timestamp 0
transform -1 0 1850 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8582_
timestamp 0
transform -1 0 1970 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8583_
timestamp 0
transform -1 0 1950 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8584_
timestamp 0
transform -1 0 1350 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8585_
timestamp 0
transform -1 0 1310 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8586_
timestamp 0
transform -1 0 1590 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8587_
timestamp 0
transform -1 0 1570 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8588_
timestamp 0
transform 1 0 1310 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8589_
timestamp 0
transform 1 0 1570 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8590_
timestamp 0
transform 1 0 1430 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8591_
timestamp 0
transform -1 0 1050 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8592_
timestamp 0
transform 1 0 1190 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8593_
timestamp 0
transform 1 0 1190 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8594_
timestamp 0
transform 1 0 1350 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8595_
timestamp 0
transform 1 0 1730 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8596_
timestamp 0
transform 1 0 1870 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8597_
timestamp 0
transform 1 0 2010 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8598_
timestamp 0
transform -1 0 3690 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8599_
timestamp 0
transform 1 0 2810 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8600_
timestamp 0
transform 1 0 1470 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8601_
timestamp 0
transform -1 0 1590 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8602_
timestamp 0
transform 1 0 550 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8603_
timestamp 0
transform 1 0 410 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8604_
timestamp 0
transform -1 0 290 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8605_
timestamp 0
transform 1 0 270 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8606_
timestamp 0
transform 1 0 2130 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8607_
timestamp 0
transform 1 0 2270 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8608_
timestamp 0
transform 1 0 2410 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8609_
timestamp 0
transform 1 0 5970 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8610_
timestamp 0
transform -1 0 6030 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8611_
timestamp 0
transform -1 0 5630 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8612_
timestamp 0
transform 1 0 5850 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8613_
timestamp 0
transform 1 0 5710 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8614_
timestamp 0
transform 1 0 5690 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8615_
timestamp 0
transform -1 0 4610 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8616_
timestamp 0
transform -1 0 4750 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8617_
timestamp 0
transform 1 0 6610 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8618_
timestamp 0
transform 1 0 6450 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8619_
timestamp 0
transform 1 0 6790 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8620_
timestamp 0
transform 1 0 6630 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8621_
timestamp 0
transform 1 0 6330 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8622_
timestamp 0
transform 1 0 6170 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8623_
timestamp 0
transform 1 0 6410 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8624_
timestamp 0
transform -1 0 6130 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8625_
timestamp 0
transform 1 0 6170 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8626_
timestamp 0
transform -1 0 6290 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8627_
timestamp 0
transform 1 0 6310 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8628_
timestamp 0
transform -1 0 6390 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8629_
timestamp 0
transform 1 0 6230 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8630_
timestamp 0
transform 1 0 6970 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8631_
timestamp 0
transform -1 0 6850 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8632_
timestamp 0
transform -1 0 6070 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8633_
timestamp 0
transform 1 0 6090 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8634_
timestamp 0
transform 1 0 5250 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8635_
timestamp 0
transform -1 0 5570 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8636_
timestamp 0
transform 1 0 5370 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8637_
timestamp 0
transform 1 0 5090 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8638_
timestamp 0
transform -1 0 5050 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8639_
timestamp 0
transform -1 0 5190 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8640_
timestamp 0
transform 1 0 6070 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8641_
timestamp 0
transform -1 0 6590 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8642_
timestamp 0
transform 1 0 6710 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8643_
timestamp 0
transform -1 0 6750 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8644_
timestamp 0
transform 1 0 6550 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8645_
timestamp 0
transform 1 0 6090 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8646_
timestamp 0
transform 1 0 6430 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8647_
timestamp 0
transform -1 0 6290 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8648_
timestamp 0
transform 1 0 5790 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8649_
timestamp 0
transform 1 0 5690 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8650_
timestamp 0
transform -1 0 5490 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8651_
timestamp 0
transform 1 0 6050 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8652_
timestamp 0
transform 1 0 5350 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8653_
timestamp 0
transform 1 0 6030 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8654_
timestamp 0
transform -1 0 5930 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8655_
timestamp 0
transform -1 0 6190 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8656_
timestamp 0
transform 1 0 6150 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8657_
timestamp 0
transform 1 0 6010 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8658_
timestamp 0
transform -1 0 5870 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8659_
timestamp 0
transform -1 0 5990 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8660_
timestamp 0
transform -1 0 7250 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8661_
timestamp 0
transform 1 0 7130 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8662_
timestamp 0
transform 1 0 6450 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8663_
timestamp 0
transform 1 0 6590 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8664_
timestamp 0
transform 1 0 6750 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8665_
timestamp 0
transform 1 0 6950 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8666_
timestamp 0
transform 1 0 6830 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8667_
timestamp 0
transform -1 0 6790 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8668_
timestamp 0
transform 1 0 6290 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8669_
timestamp 0
transform 1 0 7330 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8670_
timestamp 0
transform 1 0 7170 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8671_
timestamp 0
transform 1 0 7370 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8672_
timestamp 0
transform 1 0 7350 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8673_
timestamp 0
transform 1 0 7410 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8674_
timestamp 0
transform 1 0 5870 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8675_
timestamp 0
transform -1 0 6250 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8676_
timestamp 0
transform -1 0 6110 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8677_
timestamp 0
transform 1 0 6110 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8678_
timestamp 0
transform 1 0 7450 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8679_
timestamp 0
transform -1 0 7330 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8680_
timestamp 0
transform -1 0 7250 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8681_
timestamp 0
transform 1 0 7270 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8682_
timestamp 0
transform 1 0 6750 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8683_
timestamp 0
transform 1 0 7470 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8684_
timestamp 0
transform -1 0 7570 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8685_
timestamp 0
transform 1 0 6590 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8686_
timestamp 0
transform -1 0 6910 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8687_
timestamp 0
transform -1 0 6670 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8688_
timestamp 0
transform -1 0 6770 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8689_
timestamp 0
transform 1 0 7110 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8690_
timestamp 0
transform 1 0 6810 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8691_
timestamp 0
transform 1 0 6850 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8692_
timestamp 0
transform -1 0 5230 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8693_
timestamp 0
transform 1 0 5610 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8694_
timestamp 0
transform -1 0 5890 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8695_
timestamp 0
transform 1 0 5730 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8696_
timestamp 0
transform 1 0 6010 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8697_
timestamp 0
transform 1 0 6170 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8698_
timestamp 0
transform 1 0 6150 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8699_
timestamp 0
transform -1 0 6330 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8700_
timestamp 0
transform -1 0 6310 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8701_
timestamp 0
transform 1 0 6390 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8702_
timestamp 0
transform 1 0 6530 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8703_
timestamp 0
transform 1 0 7090 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8704_
timestamp 0
transform -1 0 7050 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8705_
timestamp 0
transform 1 0 6190 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8706_
timestamp 0
transform 1 0 7230 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8707_
timestamp 0
transform -1 0 6550 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8708_
timestamp 0
transform 1 0 6630 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8709_
timestamp 0
transform 1 0 6770 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8710_
timestamp 0
transform 1 0 6910 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8711_
timestamp 0
transform 1 0 7050 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8712_
timestamp 0
transform -1 0 6690 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8713_
timestamp 0
transform 1 0 7170 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8714_
timestamp 0
transform -1 0 6570 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8715_
timestamp 0
transform 1 0 7390 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8716_
timestamp 0
transform -1 0 7270 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8717_
timestamp 0
transform 1 0 6410 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8718_
timestamp 0
transform 1 0 6030 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8719_
timestamp 0
transform -1 0 6470 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8720_
timestamp 0
transform 1 0 6570 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8721_
timestamp 0
transform 1 0 5510 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8722_
timestamp 0
transform 1 0 5690 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8723_
timestamp 0
transform -1 0 5390 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8724_
timestamp 0
transform 1 0 5410 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8725_
timestamp 0
transform 1 0 6490 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8726_
timestamp 0
transform -1 0 6450 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8727_
timestamp 0
transform -1 0 6670 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8728_
timestamp 0
transform -1 0 6730 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8729_
timestamp 0
transform -1 0 6570 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8730_
timestamp 0
transform 1 0 5950 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8731_
timestamp 0
transform -1 0 6090 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8732_
timestamp 0
transform -1 0 6170 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8733_
timestamp 0
transform -1 0 5910 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8734_
timestamp 0
transform -1 0 5550 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8735_
timestamp 0
transform 1 0 5810 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8736_
timestamp 0
transform 1 0 6010 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8737_
timestamp 0
transform 1 0 5890 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8738_
timestamp 0
transform 1 0 5570 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8739_
timestamp 0
transform -1 0 5430 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8740_
timestamp 0
transform 1 0 5390 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__8741_
timestamp 0
transform -1 0 4830 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__8742_
timestamp 0
transform 1 0 5750 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8743_
timestamp 0
transform 1 0 6150 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8744_
timestamp 0
transform -1 0 6310 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8745_
timestamp 0
transform -1 0 5290 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8746_
timestamp 0
transform 1 0 5250 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8747_
timestamp 0
transform -1 0 4910 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8748_
timestamp 0
transform 1 0 5370 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8749_
timestamp 0
transform 1 0 5010 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8750_
timestamp 0
transform -1 0 5110 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__8751_
timestamp 0
transform 1 0 5230 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__8752_
timestamp 0
transform -1 0 4970 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__8753_
timestamp 0
transform 1 0 4290 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__8754_
timestamp 0
transform -1 0 5150 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8755_
timestamp 0
transform -1 0 4690 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__8756_
timestamp 0
transform 1 0 4070 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8757_
timestamp 0
transform 1 0 3910 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8758_
timestamp 0
transform -1 0 4050 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8759_
timestamp 0
transform -1 0 2950 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8760_
timestamp 0
transform 1 0 1030 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8761_
timestamp 0
transform -1 0 1750 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8762_
timestamp 0
transform 1 0 890 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__8763_
timestamp 0
transform 1 0 4270 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8764_
timestamp 0
transform -1 0 5230 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8765_
timestamp 0
transform -1 0 3990 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8766_
timestamp 0
transform -1 0 4150 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8767_
timestamp 0
transform -1 0 4970 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8768_
timestamp 0
transform -1 0 5090 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8769_
timestamp 0
transform 1 0 4930 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8770_
timestamp 0
transform 1 0 5210 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8771_
timestamp 0
transform -1 0 3430 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8772_
timestamp 0
transform -1 0 3550 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8773_
timestamp 0
transform -1 0 4770 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8774_
timestamp 0
transform -1 0 4890 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8775_
timestamp 0
transform 1 0 5350 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8776_
timestamp 0
transform -1 0 3790 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8777_
timestamp 0
transform 1 0 3790 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8778_
timestamp 0
transform -1 0 2770 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8779_
timestamp 0
transform -1 0 2790 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8780_
timestamp 0
transform -1 0 3950 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8781_
timestamp 0
transform 1 0 3790 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8782_
timestamp 0
transform -1 0 5230 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8783_
timestamp 0
transform 1 0 5070 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8784_
timestamp 0
transform 1 0 3270 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8785_
timestamp 0
transform 1 0 3130 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8786_
timestamp 0
transform 1 0 3130 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8787_
timestamp 0
transform 1 0 2970 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8788_
timestamp 0
transform -1 0 1690 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8789_
timestamp 0
transform 1 0 1130 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8790_
timestamp 0
transform -1 0 1470 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8791_
timestamp 0
transform 1 0 1290 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__8792_
timestamp 0
transform 1 0 5630 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8793_
timestamp 0
transform -1 0 4410 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8794_
timestamp 0
transform -1 0 4790 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8795_
timestamp 0
transform 1 0 3670 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__8796_
timestamp 0
transform -1 0 3830 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8797_
timestamp 0
transform 1 0 3670 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8798_
timestamp 0
transform 1 0 5250 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8799_
timestamp 0
transform 1 0 5110 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__8800_
timestamp 0
transform 1 0 3430 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8801_
timestamp 0
transform -1 0 3570 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__8802_
timestamp 0
transform -1 0 2490 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__8803_
timestamp 0
transform 1 0 2190 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__8804_
timestamp 0
transform -1 0 1710 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8805_
timestamp 0
transform 1 0 1550 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__8806_
timestamp 0
transform 1 0 4170 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8807_
timestamp 0
transform -1 0 4590 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8808_
timestamp 0
transform -1 0 4030 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8809_
timestamp 0
transform 1 0 3870 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8810_
timestamp 0
transform 1 0 5630 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8811_
timestamp 0
transform 1 0 5490 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__8812_
timestamp 0
transform 1 0 5570 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8813_
timestamp 0
transform 1 0 5410 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__8814_
timestamp 0
transform -1 0 4630 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8815_
timestamp 0
transform -1 0 4750 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__8816_
timestamp 0
transform -1 0 5310 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8817_
timestamp 0
transform 1 0 5130 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__8818_
timestamp 0
transform -1 0 5530 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__8819_
timestamp 0
transform 1 0 5510 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8820_
timestamp 0
transform 1 0 5430 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8821_
timestamp 0
transform -1 0 6030 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8822_
timestamp 0
transform 1 0 5650 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__8823_
timestamp 0
transform 1 0 5590 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__8824_
timestamp 0
transform -1 0 5730 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8825_
timestamp 0
transform 1 0 5310 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8826_
timestamp 0
transform -1 0 6430 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8827_
timestamp 0
transform 1 0 6250 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__8828_
timestamp 0
transform 1 0 6550 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8829_
timestamp 0
transform -1 0 6690 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8830_
timestamp 0
transform 1 0 6910 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8831_
timestamp 0
transform -1 0 7050 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__8832_
timestamp 0
transform 1 0 4730 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8833_
timestamp 0
transform -1 0 4910 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__8834_
timestamp 0
transform 1 0 5490 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8835_
timestamp 0
transform 1 0 5650 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__8836_
timestamp 0
transform -1 0 5350 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8837_
timestamp 0
transform -1 0 5470 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__8838_
timestamp 0
transform 1 0 5970 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8839_
timestamp 0
transform -1 0 5830 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__8920_
timestamp 0
transform 1 0 270 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__8921_
timestamp 0
transform -1 0 2810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__8922_
timestamp 0
transform -1 0 2930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__8923_
timestamp 0
transform -1 0 4190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__8924_
timestamp 0
transform -1 0 4050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__8925_
timestamp 0
transform 1 0 4970 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__8926_
timestamp 0
transform -1 0 4290 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__8927_
timestamp 0
transform 1 0 4170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__8928_
timestamp 0
transform 1 0 4530 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__8929_
timestamp 0
transform -1 0 4610 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__8930_
timestamp 0
transform 1 0 4470 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__8931_
timestamp 0
transform 1 0 4170 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__8932_
timestamp 0
transform 1 0 3990 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__8933_
timestamp 0
transform 1 0 3990 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__8934_
timestamp 0
transform 1 0 3730 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__8935_
timestamp 0
transform 1 0 3630 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__8936_
timestamp 0
transform 1 0 4310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__8937_
timestamp 0
transform 1 0 4470 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__8938_
timestamp 0
transform 1 0 4890 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__8939_
timestamp 0
transform -1 0 4630 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__8940_
timestamp 0
transform -1 0 4930 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__8941_
timestamp 0
transform -1 0 4790 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__8942_
timestamp 0
transform 1 0 3090 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__8943_
timestamp 0
transform 1 0 4630 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__8944_
timestamp 0
transform 1 0 5170 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__8945_
timestamp 0
transform 1 0 5590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__8946_
timestamp 0
transform 1 0 5450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__8947_
timestamp 0
transform 1 0 6230 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__8948_
timestamp 0
transform -1 0 6030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__8949_
timestamp 0
transform 1 0 5670 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__8950_
timestamp 0
transform -1 0 5370 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__8951_
timestamp 0
transform -1 0 4030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__8952_
timestamp 0
transform 1 0 4750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__8953_
timestamp 0
transform -1 0 5070 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__8954_
timestamp 0
transform -1 0 5890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__8955_
timestamp 0
transform 1 0 5570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__8956_
timestamp 0
transform 1 0 4970 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__8957_
timestamp 0
transform -1 0 4930 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__8958_
timestamp 0
transform -1 0 4970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__8959_
timestamp 0
transform -1 0 5110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__8960_
timestamp 0
transform 1 0 4690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__8961_
timestamp 0
transform 1 0 5070 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__8962_
timestamp 0
transform 1 0 3570 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__8963_
timestamp 0
transform -1 0 4810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__8964_
timestamp 0
transform 1 0 4510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__8965_
timestamp 0
transform -1 0 5830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__8966_
timestamp 0
transform 1 0 5750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__8967_
timestamp 0
transform -1 0 5530 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__8968_
timestamp 0
transform 1 0 5210 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__8969_
timestamp 0
transform -1 0 3990 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__8970_
timestamp 0
transform -1 0 4850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__8971_
timestamp 0
transform 1 0 5950 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__8972_
timestamp 0
transform -1 0 4410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__8973_
timestamp 0
transform 1 0 4610 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__8974_
timestamp 0
transform 1 0 4210 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__8975_
timestamp 0
transform -1 0 4490 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__8976_
timestamp 0
transform 1 0 4150 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__8977_
timestamp 0
transform -1 0 4350 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__8978_
timestamp 0
transform -1 0 3930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__8979_
timestamp 0
transform -1 0 2390 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__8980_
timestamp 0
transform -1 0 50 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__8981_
timestamp 0
transform -1 0 290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__8982_
timestamp 0
transform 1 0 1450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__8983_
timestamp 0
transform -1 0 1230 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__8984_
timestamp 0
transform -1 0 1370 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__8985_
timestamp 0
transform -1 0 1070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__8986_
timestamp 0
transform -1 0 910 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__8987_
timestamp 0
transform -1 0 1050 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__8988_
timestamp 0
transform -1 0 1190 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__8989_
timestamp 0
transform 1 0 910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__8990_
timestamp 0
transform -1 0 650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__8991_
timestamp 0
transform -1 0 790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__8992_
timestamp 0
transform -1 0 1590 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__8993_
timestamp 0
transform 1 0 1430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__8994_
timestamp 0
transform -1 0 1410 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__8995_
timestamp 0
transform 1 0 1050 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__8996_
timestamp 0
transform 1 0 1230 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__8997_
timestamp 0
transform -1 0 2510 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__8998_
timestamp 0
transform -1 0 2250 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__8999_
timestamp 0
transform -1 0 2630 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9000_
timestamp 0
transform -1 0 450 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9001_
timestamp 0
transform 1 0 3550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9002_
timestamp 0
transform 1 0 3430 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9003_
timestamp 0
transform 1 0 2710 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9004_
timestamp 0
transform -1 0 3550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9005_
timestamp 0
transform 1 0 4510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9006_
timestamp 0
transform 1 0 4570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9007_
timestamp 0
transform -1 0 3590 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9008_
timestamp 0
transform -1 0 450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9009_
timestamp 0
transform -1 0 570 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9010_
timestamp 0
transform 1 0 390 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9011_
timestamp 0
transform 1 0 30 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9012_
timestamp 0
transform -1 0 190 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9013_
timestamp 0
transform 1 0 310 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9014_
timestamp 0
transform -1 0 610 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9015_
timestamp 0
transform -1 0 770 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9016_
timestamp 0
transform -1 0 470 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9017_
timestamp 0
transform 1 0 450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9018_
timestamp 0
transform -1 0 1310 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9019_
timestamp 0
transform -1 0 150 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9020_
timestamp 0
transform -1 0 1070 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9021_
timestamp 0
transform -1 0 810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9022_
timestamp 0
transform -1 0 950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9023_
timestamp 0
transform -1 0 1670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9024_
timestamp 0
transform -1 0 1250 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9025_
timestamp 0
transform -1 0 1390 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9026_
timestamp 0
transform 1 0 1050 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9027_
timestamp 0
transform 1 0 910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9028_
timestamp 0
transform 1 0 1510 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9029_
timestamp 0
transform -1 0 1510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9030_
timestamp 0
transform -1 0 1190 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9031_
timestamp 0
transform 1 0 1690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9032_
timestamp 0
transform 1 0 1650 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9033_
timestamp 0
transform 1 0 1470 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9034_
timestamp 0
transform 1 0 1530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9035_
timestamp 0
transform 1 0 1530 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9036_
timestamp 0
transform 1 0 730 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9037_
timestamp 0
transform 1 0 730 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9038_
timestamp 0
transform -1 0 770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9039_
timestamp 0
transform -1 0 770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9040_
timestamp 0
transform -1 0 1030 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9041_
timestamp 0
transform 1 0 730 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9042_
timestamp 0
transform -1 0 910 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9043_
timestamp 0
transform -1 0 1690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9044_
timestamp 0
transform -1 0 1570 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9045_
timestamp 0
transform 1 0 1830 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9046_
timestamp 0
transform 1 0 1690 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9047_
timestamp 0
transform 1 0 1950 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9048_
timestamp 0
transform 1 0 2650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9049_
timestamp 0
transform 1 0 2810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9050_
timestamp 0
transform 1 0 2950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9051_
timestamp 0
transform 1 0 4190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9052_
timestamp 0
transform 1 0 7510 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9053_
timestamp 0
transform -1 0 6930 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9054_
timestamp 0
transform 1 0 7130 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9055_
timestamp 0
transform -1 0 3970 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9056_
timestamp 0
transform -1 0 2110 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9057_
timestamp 0
transform -1 0 450 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9058_
timestamp 0
transform 1 0 590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9059_
timestamp 0
transform -1 0 610 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9060_
timestamp 0
transform -1 0 310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9061_
timestamp 0
transform 1 0 430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9062_
timestamp 0
transform 1 0 570 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9063_
timestamp 0
transform 1 0 1970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9064_
timestamp 0
transform 1 0 2110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9065_
timestamp 0
transform 1 0 2090 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9066_
timestamp 0
transform 1 0 1670 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9067_
timestamp 0
transform 1 0 1950 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9068_
timestamp 0
transform 1 0 2410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9069_
timestamp 0
transform 1 0 2250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9070_
timestamp 0
transform 1 0 3270 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9071_
timestamp 0
transform 1 0 3530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9072_
timestamp 0
transform 1 0 3690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9073_
timestamp 0
transform 1 0 3810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9074_
timestamp 0
transform -1 0 3390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9075_
timestamp 0
transform 1 0 3910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9076_
timestamp 0
transform 1 0 4010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9077_
timestamp 0
transform 1 0 4370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9078_
timestamp 0
transform -1 0 4070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9079_
timestamp 0
transform 1 0 4850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9080_
timestamp 0
transform 1 0 4470 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9081_
timestamp 0
transform 1 0 3110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9082_
timestamp 0
transform 1 0 3970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9083_
timestamp 0
transform -1 0 2930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9084_
timestamp 0
transform 1 0 1830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9085_
timestamp 0
transform 1 0 550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9086_
timestamp 0
transform -1 0 330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9087_
timestamp 0
transform -1 0 670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9088_
timestamp 0
transform -1 0 930 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9089_
timestamp 0
transform 1 0 910 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9090_
timestamp 0
transform -1 0 1650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9091_
timestamp 0
transform 1 0 1530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9092_
timestamp 0
transform 1 0 1630 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9093_
timestamp 0
transform 1 0 1550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9094_
timestamp 0
transform 1 0 2630 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9095_
timestamp 0
transform -1 0 2670 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9096_
timestamp 0
transform -1 0 2790 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9097_
timestamp 0
transform -1 0 2790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9098_
timestamp 0
transform 1 0 3170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9099_
timestamp 0
transform 1 0 3030 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9100_
timestamp 0
transform 1 0 3490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9101_
timestamp 0
transform 1 0 3610 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9102_
timestamp 0
transform 1 0 4070 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9103_
timestamp 0
transform 1 0 4230 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9104_
timestamp 0
transform -1 0 4590 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9105_
timestamp 0
transform 1 0 3330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9106_
timestamp 0
transform 1 0 3550 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9107_
timestamp 0
transform -1 0 210 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9108_
timestamp 0
transform -1 0 390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9109_
timestamp 0
transform 1 0 490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9110_
timestamp 0
transform 1 0 630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9111_
timestamp 0
transform -1 0 790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9112_
timestamp 0
transform -1 0 950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9113_
timestamp 0
transform -1 0 1090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9114_
timestamp 0
transform 1 0 3330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9115_
timestamp 0
transform 1 0 3210 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9116_
timestamp 0
transform 1 0 3630 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9117_
timestamp 0
transform -1 0 2950 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9118_
timestamp 0
transform 1 0 3070 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9119_
timestamp 0
transform 1 0 3930 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9120_
timestamp 0
transform -1 0 3610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9121_
timestamp 0
transform -1 0 3470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9122_
timestamp 0
transform 1 0 3710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9123_
timestamp 0
transform 1 0 4350 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9124_
timestamp 0
transform 1 0 4910 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9125_
timestamp 0
transform 1 0 5070 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9126_
timestamp 0
transform -1 0 5830 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9127_
timestamp 0
transform -1 0 4290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9128_
timestamp 0
transform 1 0 2830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9129_
timestamp 0
transform 1 0 2930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9130_
timestamp 0
transform -1 0 450 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9131_
timestamp 0
transform 1 0 550 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9132_
timestamp 0
transform 1 0 990 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9133_
timestamp 0
transform -1 0 1070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9134_
timestamp 0
transform -1 0 1330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9135_
timestamp 0
transform 1 0 2630 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9136_
timestamp 0
transform -1 0 3110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9137_
timestamp 0
transform -1 0 2710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9138_
timestamp 0
transform -1 0 2810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9139_
timestamp 0
transform 1 0 3370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9140_
timestamp 0
transform 1 0 3230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9141_
timestamp 0
transform -1 0 3530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9142_
timestamp 0
transform -1 0 3650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9143_
timestamp 0
transform 1 0 4410 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9144_
timestamp 0
transform 1 0 4570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9145_
timestamp 0
transform 1 0 4710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9146_
timestamp 0
transform -1 0 4710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9147_
timestamp 0
transform -1 0 6330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9148_
timestamp 0
transform 1 0 4510 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9149_
timestamp 0
transform 1 0 3090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9150_
timestamp 0
transform 1 0 670 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9151_
timestamp 0
transform -1 0 630 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9152_
timestamp 0
transform -1 0 850 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9153_
timestamp 0
transform 1 0 4090 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9154_
timestamp 0
transform -1 0 3330 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9155_
timestamp 0
transform 1 0 2770 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9156_
timestamp 0
transform -1 0 3550 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9157_
timestamp 0
transform 1 0 4910 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9158_
timestamp 0
transform 1 0 3650 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9159_
timestamp 0
transform -1 0 3430 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9160_
timestamp 0
transform 1 0 3790 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9161_
timestamp 0
transform 1 0 5030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9162_
timestamp 0
transform 1 0 3770 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9163_
timestamp 0
transform 1 0 4090 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9164_
timestamp 0
transform -1 0 4770 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9165_
timestamp 0
transform 1 0 4670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9166_
timestamp 0
transform 1 0 5150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9167_
timestamp 0
transform 1 0 5290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9168_
timestamp 0
transform -1 0 6170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9169_
timestamp 0
transform 1 0 5030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9170_
timestamp 0
transform -1 0 4790 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9171_
timestamp 0
transform 1 0 4210 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9172_
timestamp 0
transform -1 0 4070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9173_
timestamp 0
transform -1 0 3770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9174_
timestamp 0
transform -1 0 3910 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9175_
timestamp 0
transform -1 0 4650 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9176_
timestamp 0
transform -1 0 4190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9177_
timestamp 0
transform -1 0 2970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9178_
timestamp 0
transform 1 0 270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9179_
timestamp 0
transform -1 0 410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9180_
timestamp 0
transform 1 0 670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9181_
timestamp 0
transform -1 0 1490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9182_
timestamp 0
transform -1 0 3230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9183_
timestamp 0
transform -1 0 3370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9184_
timestamp 0
transform 1 0 3950 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9185_
timestamp 0
transform 1 0 3890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9186_
timestamp 0
transform 1 0 4010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9187_
timestamp 0
transform 1 0 3470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9188_
timestamp 0
transform 1 0 3750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9189_
timestamp 0
transform -1 0 3630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9190_
timestamp 0
transform -1 0 4150 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9191_
timestamp 0
transform 1 0 4250 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9192_
timestamp 0
transform 1 0 4510 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9193_
timestamp 0
transform 1 0 4870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9194_
timestamp 0
transform 1 0 4370 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9195_
timestamp 0
transform 1 0 4310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9196_
timestamp 0
transform 1 0 4770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9197_
timestamp 0
transform 1 0 4630 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9198_
timestamp 0
transform -1 0 4890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9199_
timestamp 0
transform -1 0 5050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9200_
timestamp 0
transform -1 0 3730 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9201_
timestamp 0
transform -1 0 4030 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9202_
timestamp 0
transform -1 0 3890 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9203_
timestamp 0
transform -1 0 2370 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9204_
timestamp 0
transform -1 0 3210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9205_
timestamp 0
transform 1 0 1150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9206_
timestamp 0
transform -1 0 2790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9207_
timestamp 0
transform 1 0 2870 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9208_
timestamp 0
transform 1 0 2630 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9209_
timestamp 0
transform -1 0 2750 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9210_
timestamp 0
transform 1 0 2470 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9211_
timestamp 0
transform 1 0 2910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9212_
timestamp 0
transform 1 0 3010 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9213_
timestamp 0
transform 1 0 3050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9214_
timestamp 0
transform 1 0 4190 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9215_
timestamp 0
transform 1 0 4490 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9216_
timestamp 0
transform 1 0 4470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9217_
timestamp 0
transform 1 0 4610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9218_
timestamp 0
transform -1 0 4890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9219_
timestamp 0
transform -1 0 4310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9220_
timestamp 0
transform 1 0 4430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9221_
timestamp 0
transform 1 0 5070 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9222_
timestamp 0
transform 1 0 4710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9223_
timestamp 0
transform -1 0 4590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9224_
timestamp 0
transform -1 0 4090 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9225_
timestamp 0
transform 1 0 4350 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9226_
timestamp 0
transform -1 0 3650 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9227_
timestamp 0
transform 1 0 3330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9228_
timestamp 0
transform 1 0 3530 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9229_
timestamp 0
transform 1 0 1310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9230_
timestamp 0
transform 1 0 3390 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9231_
timestamp 0
transform 1 0 3130 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9232_
timestamp 0
transform 1 0 3310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9233_
timestamp 0
transform 1 0 3450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9234_
timestamp 0
transform 1 0 3750 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9235_
timestamp 0
transform -1 0 3270 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9236_
timestamp 0
transform 1 0 3910 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9237_
timestamp 0
transform 1 0 4030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9238_
timestamp 0
transform 1 0 4450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9239_
timestamp 0
transform 1 0 4590 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9240_
timestamp 0
transform 1 0 4730 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9241_
timestamp 0
transform -1 0 5170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9242_
timestamp 0
transform -1 0 2270 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9243_
timestamp 0
transform 1 0 890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9244_
timestamp 0
transform 1 0 3410 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9245_
timestamp 0
transform 1 0 3650 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9246_
timestamp 0
transform 1 0 3510 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9247_
timestamp 0
transform -1 0 3710 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9248_
timestamp 0
transform -1 0 3290 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9249_
timestamp 0
transform 1 0 3810 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9250_
timestamp 0
transform 1 0 3730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9251_
timestamp 0
transform 1 0 4090 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9252_
timestamp 0
transform 1 0 3810 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9253_
timestamp 0
transform -1 0 3970 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9254_
timestamp 0
transform 1 0 3950 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9255_
timestamp 0
transform -1 0 4110 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9256_
timestamp 0
transform 1 0 3590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9257_
timestamp 0
transform -1 0 3890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9258_
timestamp 0
transform -1 0 4330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9259_
timestamp 0
transform 1 0 4390 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9260_
timestamp 0
transform 1 0 4230 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9261_
timestamp 0
transform 1 0 4170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9262_
timestamp 0
transform 1 0 4530 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9263_
timestamp 0
transform 1 0 4690 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9264_
timestamp 0
transform 1 0 4830 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9265_
timestamp 0
transform -1 0 4790 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9266_
timestamp 0
transform 1 0 6210 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9267_
timestamp 0
transform -1 0 4210 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9268_
timestamp 0
transform 1 0 30 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9269_
timestamp 0
transform 1 0 270 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9270_
timestamp 0
transform -1 0 290 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9271_
timestamp 0
transform -1 0 50 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9272_
timestamp 0
transform -1 0 3570 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9273_
timestamp 0
transform 1 0 3810 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9274_
timestamp 0
transform 1 0 3930 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9275_
timestamp 0
transform 1 0 4070 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9276_
timestamp 0
transform -1 0 4210 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9277_
timestamp 0
transform 1 0 4450 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9278_
timestamp 0
transform -1 0 4330 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9279_
timestamp 0
transform 1 0 4310 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9280_
timestamp 0
transform 1 0 4670 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9281_
timestamp 0
transform -1 0 6090 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9282_
timestamp 0
transform 1 0 3570 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9283_
timestamp 0
transform 1 0 2550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9284_
timestamp 0
transform 1 0 2890 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9285_
timestamp 0
transform 1 0 2470 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9286_
timestamp 0
transform 1 0 1970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9287_
timestamp 0
transform 1 0 1690 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9288_
timestamp 0
transform -1 0 550 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9289_
timestamp 0
transform -1 0 1550 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9290_
timestamp 0
transform 1 0 1830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9291_
timestamp 0
transform -1 0 4250 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9292_
timestamp 0
transform -1 0 4390 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9293_
timestamp 0
transform -1 0 2370 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9294_
timestamp 0
transform -1 0 2510 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9295_
timestamp 0
transform -1 0 2370 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9296_
timestamp 0
transform -1 0 1930 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9297_
timestamp 0
transform -1 0 1930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9298_
timestamp 0
transform 1 0 1810 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9299_
timestamp 0
transform 1 0 2530 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9300_
timestamp 0
transform 1 0 2770 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9301_
timestamp 0
transform 1 0 2650 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9302_
timestamp 0
transform 1 0 1990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9303_
timestamp 0
transform 1 0 2310 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9304_
timestamp 0
transform 1 0 3190 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9305_
timestamp 0
transform -1 0 3850 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9306_
timestamp 0
transform -1 0 2210 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9307_
timestamp 0
transform 1 0 3250 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9308_
timestamp 0
transform 1 0 3110 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9309_
timestamp 0
transform 1 0 1430 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9310_
timestamp 0
transform 1 0 1270 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9311_
timestamp 0
transform -1 0 1810 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9312_
timestamp 0
transform 1 0 1850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9313_
timestamp 0
transform -1 0 2970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9314_
timestamp 0
transform -1 0 3090 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9315_
timestamp 0
transform 1 0 1270 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9316_
timestamp 0
transform -1 0 2310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9317_
timestamp 0
transform -1 0 2430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9318_
timestamp 0
transform -1 0 1570 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9319_
timestamp 0
transform 1 0 1390 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9320_
timestamp 0
transform 1 0 1710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9321_
timestamp 0
transform 1 0 1950 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9322_
timestamp 0
transform -1 0 2190 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9323_
timestamp 0
transform 1 0 2130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9324_
timestamp 0
transform -1 0 2210 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9325_
timestamp 0
transform 1 0 2210 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9326_
timestamp 0
transform 1 0 2370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9327_
timestamp 0
transform 1 0 2350 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9328_
timestamp 0
transform 1 0 2490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9329_
timestamp 0
transform -1 0 2630 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9330_
timestamp 0
transform 1 0 2750 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9331_
timestamp 0
transform 1 0 3030 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9332_
timestamp 0
transform 1 0 3690 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9333_
timestamp 0
transform 1 0 4050 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9334_
timestamp 0
transform 1 0 2490 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9335_
timestamp 0
transform -1 0 2170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9336_
timestamp 0
transform 1 0 2110 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9337_
timestamp 0
transform -1 0 1990 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9338_
timestamp 0
transform 1 0 2370 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9339_
timestamp 0
transform 1 0 1850 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9340_
timestamp 0
transform 1 0 1790 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9341_
timestamp 0
transform -1 0 1810 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9342_
timestamp 0
transform -1 0 1690 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9343_
timestamp 0
transform 1 0 1690 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9344_
timestamp 0
transform 1 0 1990 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9345_
timestamp 0
transform 1 0 2230 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9346_
timestamp 0
transform 1 0 2030 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9347_
timestamp 0
transform -1 0 2030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9348_
timestamp 0
transform 1 0 2270 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9349_
timestamp 0
transform 1 0 2730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9350_
timestamp 0
transform 1 0 2430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9351_
timestamp 0
transform 1 0 2830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9352_
timestamp 0
transform 1 0 3490 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9353_
timestamp 0
transform -1 0 3370 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9354_
timestamp 0
transform 1 0 3870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9355_
timestamp 0
transform 1 0 3890 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9356_
timestamp 0
transform -1 0 2610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9357_
timestamp 0
transform -1 0 2530 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9358_
timestamp 0
transform -1 0 2290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9359_
timestamp 0
transform 1 0 2130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9360_
timestamp 0
transform -1 0 1090 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9361_
timestamp 0
transform -1 0 1270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9362_
timestamp 0
transform 1 0 2050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9363_
timestamp 0
transform -1 0 1950 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9364_
timestamp 0
transform -1 0 2070 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9365_
timestamp 0
transform 1 0 1370 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9366_
timestamp 0
transform -1 0 2110 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9367_
timestamp 0
transform 1 0 1930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9368_
timestamp 0
transform 1 0 1790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9369_
timestamp 0
transform 1 0 2230 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9370_
timestamp 0
transform 1 0 2530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9371_
timestamp 0
transform 1 0 2090 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9372_
timestamp 0
transform 1 0 2630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9373_
timestamp 0
transform 1 0 3310 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9374_
timestamp 0
transform -1 0 3190 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9375_
timestamp 0
transform 1 0 3450 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9376_
timestamp 0
transform -1 0 5470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9377_
timestamp 0
transform -1 0 2410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9378_
timestamp 0
transform -1 0 170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9379_
timestamp 0
transform -1 0 830 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9380_
timestamp 0
transform -1 0 1430 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9381_
timestamp 0
transform -1 0 1550 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9382_
timestamp 0
transform -1 0 1310 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9383_
timestamp 0
transform -1 0 1430 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9384_
timestamp 0
transform 1 0 1850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9385_
timestamp 0
transform -1 0 1770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9386_
timestamp 0
transform -1 0 1710 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9387_
timestamp 0
transform -1 0 1730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9388_
timestamp 0
transform -1 0 1570 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9389_
timestamp 0
transform -1 0 1450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9390_
timestamp 0
transform 1 0 1570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9391_
timestamp 0
transform 1 0 1970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9392_
timestamp 0
transform -1 0 1750 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9393_
timestamp 0
transform 1 0 2010 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9394_
timestamp 0
transform -1 0 2450 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9395_
timestamp 0
transform 1 0 2690 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9396_
timestamp 0
transform 1 0 2550 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9397_
timestamp 0
transform 1 0 2690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9398_
timestamp 0
transform -1 0 5650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9399_
timestamp 0
transform 1 0 4210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9400_
timestamp 0
transform 1 0 2550 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9401_
timestamp 0
transform -1 0 1810 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9402_
timestamp 0
transform -1 0 550 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9403_
timestamp 0
transform -1 0 990 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9404_
timestamp 0
transform 1 0 1290 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9405_
timestamp 0
transform 1 0 1130 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9406_
timestamp 0
transform 1 0 1570 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9407_
timestamp 0
transform 1 0 1910 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9408_
timestamp 0
transform -1 0 1550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9409_
timestamp 0
transform 1 0 1650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9410_
timestamp 0
transform 1 0 1570 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9411_
timestamp 0
transform -1 0 1690 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9412_
timestamp 0
transform -1 0 1850 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9413_
timestamp 0
transform -1 0 2170 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9414_
timestamp 0
transform 1 0 1990 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9415_
timestamp 0
transform -1 0 2270 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9416_
timestamp 0
transform -1 0 3030 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9417_
timestamp 0
transform 1 0 3130 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9418_
timestamp 0
transform 1 0 3290 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9419_
timestamp 0
transform -1 0 3830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9420_
timestamp 0
transform -1 0 5390 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9421_
timestamp 0
transform -1 0 1450 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9422_
timestamp 0
transform -1 0 670 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9423_
timestamp 0
transform -1 0 630 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9424_
timestamp 0
transform -1 0 1030 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9425_
timestamp 0
transform 1 0 1010 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9426_
timestamp 0
transform -1 0 1370 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9427_
timestamp 0
transform 1 0 890 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9428_
timestamp 0
transform -1 0 1170 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9429_
timestamp 0
transform -1 0 1310 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9430_
timestamp 0
transform 1 0 1430 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9431_
timestamp 0
transform 1 0 1550 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9432_
timestamp 0
transform 1 0 1710 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9433_
timestamp 0
transform -1 0 1890 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9434_
timestamp 0
transform 1 0 2270 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9435_
timestamp 0
transform -1 0 2430 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9436_
timestamp 0
transform 1 0 2390 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9437_
timestamp 0
transform 1 0 2530 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9438_
timestamp 0
transform 1 0 2710 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9439_
timestamp 0
transform -1 0 2150 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9440_
timestamp 0
transform -1 0 2030 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9441_
timestamp 0
transform -1 0 1870 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9442_
timestamp 0
transform -1 0 1730 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9443_
timestamp 0
transform 1 0 2870 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9444_
timestamp 0
transform 1 0 3670 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9445_
timestamp 0
transform -1 0 3710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9446_
timestamp 0
transform -1 0 5230 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9447_
timestamp 0
transform -1 0 3730 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9448_
timestamp 0
transform 1 0 2650 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9449_
timestamp 0
transform 1 0 770 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9450_
timestamp 0
transform -1 0 410 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9451_
timestamp 0
transform 1 0 450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9452_
timestamp 0
transform -1 0 750 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9453_
timestamp 0
transform -1 0 150 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9454_
timestamp 0
transform -1 0 50 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9455_
timestamp 0
transform -1 0 1010 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9456_
timestamp 0
transform -1 0 610 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9457_
timestamp 0
transform 1 0 450 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9458_
timestamp 0
transform 1 0 290 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9459_
timestamp 0
transform -1 0 730 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9460_
timestamp 0
transform 1 0 830 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9461_
timestamp 0
transform -1 0 1170 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9462_
timestamp 0
transform 1 0 2770 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9463_
timestamp 0
transform 1 0 3030 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9464_
timestamp 0
transform 1 0 2930 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9465_
timestamp 0
transform 1 0 3150 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9466_
timestamp 0
transform -1 0 3330 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9467_
timestamp 0
transform -1 0 1290 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9468_
timestamp 0
transform -1 0 1610 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9469_
timestamp 0
transform -1 0 1450 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__9470_
timestamp 0
transform -1 0 710 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9471_
timestamp 0
transform -1 0 650 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9472_
timestamp 0
transform -1 0 1190 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9473_
timestamp 0
transform -1 0 890 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9474_
timestamp 0
transform 1 0 890 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9475_
timestamp 0
transform 1 0 750 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9476_
timestamp 0
transform -1 0 510 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9477_
timestamp 0
transform 1 0 610 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9478_
timestamp 0
transform 1 0 790 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9479_
timestamp 0
transform 1 0 330 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9480_
timestamp 0
transform 1 0 1010 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9481_
timestamp 0
transform 1 0 1130 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9482_
timestamp 0
transform 1 0 2230 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9483_
timestamp 0
transform 1 0 2510 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9484_
timestamp 0
transform 1 0 2070 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9485_
timestamp 0
transform 1 0 2370 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9486_
timestamp 0
transform -1 0 3170 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9487_
timestamp 0
transform 1 0 3010 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9488_
timestamp 0
transform -1 0 2190 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9489_
timestamp 0
transform 1 0 2290 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9490_
timestamp 0
transform -1 0 490 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9491_
timestamp 0
transform -1 0 310 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9492_
timestamp 0
transform 1 0 470 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9493_
timestamp 0
transform -1 0 430 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9494_
timestamp 0
transform 1 0 550 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9495_
timestamp 0
transform 1 0 530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9496_
timestamp 0
transform -1 0 410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9497_
timestamp 0
transform -1 0 690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9498_
timestamp 0
transform 1 0 1290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9499_
timestamp 0
transform 1 0 2390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9500_
timestamp 0
transform 1 0 2530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9501_
timestamp 0
transform 1 0 2630 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9502_
timestamp 0
transform 1 0 5110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9503_
timestamp 0
transform 1 0 930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9504_
timestamp 0
transform 1 0 930 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9505_
timestamp 0
transform 1 0 1290 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9506_
timestamp 0
transform -1 0 1230 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9507_
timestamp 0
transform -1 0 1090 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9508_
timestamp 0
transform -1 0 330 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9509_
timestamp 0
transform 1 0 290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9510_
timestamp 0
transform -1 0 190 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9511_
timestamp 0
transform -1 0 50 0 1 250
box -6 -8 26 248
use FILL  FILL_1__9512_
timestamp 0
transform 1 0 330 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9513_
timestamp 0
transform -1 0 50 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9514_
timestamp 0
transform -1 0 50 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9515_
timestamp 0
transform 1 0 170 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9516_
timestamp 0
transform 1 0 170 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9517_
timestamp 0
transform 1 0 150 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9518_
timestamp 0
transform -1 0 50 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__9519_
timestamp 0
transform -1 0 50 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9520_
timestamp 0
transform 1 0 190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__9521_
timestamp 0
transform 1 0 150 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__9522_
timestamp 0
transform -1 0 4950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__9523_
timestamp 0
transform -1 0 3210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9524_
timestamp 0
transform 1 0 30 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9525_
timestamp 0
transform 1 0 150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__9526_
timestamp 0
transform 1 0 2610 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9527_
timestamp 0
transform -1 0 2750 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9528_
timestamp 0
transform 1 0 3010 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9529_
timestamp 0
transform -1 0 2890 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__9530_
timestamp 0
transform 1 0 2830 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9531_
timestamp 0
transform 1 0 2970 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9532_
timestamp 0
transform 1 0 3130 0 1 730
box -6 -8 26 248
use FILL  FILL_1__9533_
timestamp 0
transform 1 0 750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9534_
timestamp 0
transform 1 0 1410 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9535_
timestamp 0
transform 1 0 1570 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9536_
timestamp 0
transform 1 0 1270 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9537_
timestamp 0
transform -1 0 1590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9538_
timestamp 0
transform 1 0 1690 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9539_
timestamp 0
transform 1 0 3610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9540_
timestamp 0
transform 1 0 3230 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9541_
timestamp 0
transform 1 0 2070 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9542_
timestamp 0
transform -1 0 1490 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9543_
timestamp 0
transform 1 0 1250 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9544_
timestamp 0
transform -1 0 1170 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9545_
timestamp 0
transform 1 0 970 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9546_
timestamp 0
transform 1 0 810 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9547_
timestamp 0
transform -1 0 850 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9548_
timestamp 0
transform 1 0 850 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9549_
timestamp 0
transform -1 0 390 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9550_
timestamp 0
transform -1 0 710 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9551_
timestamp 0
transform -1 0 530 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9552_
timestamp 0
transform -1 0 1450 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9553_
timestamp 0
transform -1 0 1310 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9554_
timestamp 0
transform -1 0 1570 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9555_
timestamp 0
transform 1 0 1670 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9556_
timestamp 0
transform 1 0 630 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9557_
timestamp 0
transform 1 0 1010 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9558_
timestamp 0
transform 1 0 150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9559_
timestamp 0
transform 1 0 30 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9560_
timestamp 0
transform -1 0 190 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9561_
timestamp 0
transform -1 0 210 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9562_
timestamp 0
transform -1 0 50 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9563_
timestamp 0
transform -1 0 50 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9564_
timestamp 0
transform -1 0 50 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9565_
timestamp 0
transform 1 0 250 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9566_
timestamp 0
transform -1 0 150 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9567_
timestamp 0
transform -1 0 570 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9568_
timestamp 0
transform -1 0 410 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9569_
timestamp 0
transform -1 0 2090 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9570_
timestamp 0
transform -1 0 170 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9571_
timestamp 0
transform 1 0 290 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9572_
timestamp 0
transform -1 0 910 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9573_
timestamp 0
transform -1 0 50 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9574_
timestamp 0
transform 1 0 450 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9575_
timestamp 0
transform -1 0 590 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9576_
timestamp 0
transform -1 0 630 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9577_
timestamp 0
transform 1 0 630 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9578_
timestamp 0
transform 1 0 770 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9579_
timestamp 0
transform -1 0 710 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9580_
timestamp 0
transform -1 0 590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9581_
timestamp 0
transform -1 0 410 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9582_
timestamp 0
transform 1 0 550 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9583_
timestamp 0
transform -1 0 1970 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9584_
timestamp 0
transform 1 0 4330 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9585_
timestamp 0
transform 1 0 3070 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9586_
timestamp 0
transform 1 0 970 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9587_
timestamp 0
transform -1 0 1150 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9588_
timestamp 0
transform 1 0 1090 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9589_
timestamp 0
transform 1 0 3170 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9590_
timestamp 0
transform 1 0 3330 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9591_
timestamp 0
transform 1 0 3450 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9592_
timestamp 0
transform 1 0 690 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9593_
timestamp 0
transform 1 0 3850 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9594_
timestamp 0
transform -1 0 3730 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9595_
timestamp 0
transform 1 0 3750 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9596_
timestamp 0
transform -1 0 3690 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9597_
timestamp 0
transform -1 0 2410 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9598_
timestamp 0
transform -1 0 1490 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9599_
timestamp 0
transform -1 0 1150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9600_
timestamp 0
transform 1 0 1370 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9601_
timestamp 0
transform 1 0 1510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9602_
timestamp 0
transform 1 0 2870 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9603_
timestamp 0
transform -1 0 2750 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9604_
timestamp 0
transform -1 0 3030 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9605_
timestamp 0
transform 1 0 3270 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9606_
timestamp 0
transform 1 0 3870 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9607_
timestamp 0
transform -1 0 3770 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9608_
timestamp 0
transform -1 0 4670 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9609_
timestamp 0
transform -1 0 4810 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9610_
timestamp 0
transform -1 0 4470 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9611_
timestamp 0
transform -1 0 3590 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9612_
timestamp 0
transform -1 0 3850 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9613_
timestamp 0
transform -1 0 3150 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9614_
timestamp 0
transform 1 0 3390 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9615_
timestamp 0
transform 1 0 3970 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9616_
timestamp 0
transform 1 0 310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9617_
timestamp 0
transform 1 0 350 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9618_
timestamp 0
transform 1 0 310 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9619_
timestamp 0
transform 1 0 490 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9620_
timestamp 0
transform -1 0 450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9621_
timestamp 0
transform -1 0 2450 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9622_
timestamp 0
transform 1 0 2450 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9623_
timestamp 0
transform -1 0 2770 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9624_
timestamp 0
transform 1 0 2990 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9625_
timestamp 0
transform 1 0 4250 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9626_
timestamp 0
transform -1 0 4150 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9627_
timestamp 0
transform -1 0 4530 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9628_
timestamp 0
transform 1 0 4370 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9629_
timestamp 0
transform -1 0 4610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9630_
timestamp 0
transform 1 0 4010 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9631_
timestamp 0
transform -1 0 2290 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9632_
timestamp 0
transform 1 0 1390 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9633_
timestamp 0
transform 1 0 1510 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9634_
timestamp 0
transform -1 0 1670 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9635_
timestamp 0
transform -1 0 2050 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9636_
timestamp 0
transform 1 0 2210 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9637_
timestamp 0
transform -1 0 2170 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9638_
timestamp 0
transform 1 0 2330 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9639_
timestamp 0
transform 1 0 4130 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9640_
timestamp 0
transform 1 0 4130 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9641_
timestamp 0
transform -1 0 4290 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9642_
timestamp 0
transform 1 0 3910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9643_
timestamp 0
transform -1 0 1350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9644_
timestamp 0
transform 1 0 1630 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9645_
timestamp 0
transform 1 0 1950 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9646_
timestamp 0
transform 1 0 2810 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9647_
timestamp 0
transform 1 0 1950 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9648_
timestamp 0
transform 1 0 2670 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9649_
timestamp 0
transform -1 0 2630 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9650_
timestamp 0
transform -1 0 2890 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9651_
timestamp 0
transform 1 0 3110 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9652_
timestamp 0
transform -1 0 3450 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9653_
timestamp 0
transform -1 0 3290 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9654_
timestamp 0
transform -1 0 3310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9655_
timestamp 0
transform -1 0 3270 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9656_
timestamp 0
transform -1 0 3430 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9657_
timestamp 0
transform 1 0 3530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9658_
timestamp 0
transform -1 0 2950 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9659_
timestamp 0
transform 1 0 2110 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9660_
timestamp 0
transform -1 0 1990 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9661_
timestamp 0
transform -1 0 2390 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9662_
timestamp 0
transform -1 0 2850 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9663_
timestamp 0
transform 1 0 2990 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9664_
timestamp 0
transform -1 0 3150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9665_
timestamp 0
transform -1 0 3630 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9666_
timestamp 0
transform -1 0 2570 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9667_
timestamp 0
transform 1 0 2390 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9668_
timestamp 0
transform 1 0 2570 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9669_
timestamp 0
transform -1 0 2710 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9670_
timestamp 0
transform 1 0 2670 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9671_
timestamp 0
transform -1 0 2810 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9672_
timestamp 0
transform 1 0 2650 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9673_
timestamp 0
transform 1 0 2910 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9674_
timestamp 0
transform 1 0 3170 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9675_
timestamp 0
transform 1 0 3330 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9676_
timestamp 0
transform 1 0 3470 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9677_
timestamp 0
transform -1 0 4170 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9678_
timestamp 0
transform -1 0 3050 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9679_
timestamp 0
transform 1 0 3990 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9680_
timestamp 0
transform -1 0 3010 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9681_
timestamp 0
transform -1 0 3610 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9682_
timestamp 0
transform -1 0 2870 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9683_
timestamp 0
transform -1 0 190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9684_
timestamp 0
transform -1 0 290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9685_
timestamp 0
transform -1 0 50 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9686_
timestamp 0
transform -1 0 50 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9687_
timestamp 0
transform -1 0 210 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9688_
timestamp 0
transform -1 0 450 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9689_
timestamp 0
transform 1 0 690 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9690_
timestamp 0
transform -1 0 870 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9691_
timestamp 0
transform -1 0 50 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9692_
timestamp 0
transform -1 0 450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9693_
timestamp 0
transform -1 0 310 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9694_
timestamp 0
transform 1 0 4350 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9695_
timestamp 0
transform -1 0 50 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9696_
timestamp 0
transform -1 0 50 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9697_
timestamp 0
transform -1 0 170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9698_
timestamp 0
transform -1 0 290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9699_
timestamp 0
transform -1 0 3670 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9700_
timestamp 0
transform 1 0 1410 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9701_
timestamp 0
transform 1 0 1250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9702_
timestamp 0
transform 1 0 1350 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9703_
timestamp 0
transform -1 0 1770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9704_
timestamp 0
transform 1 0 1150 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9705_
timestamp 0
transform 1 0 990 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9706_
timestamp 0
transform -1 0 690 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9707_
timestamp 0
transform 1 0 390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9708_
timestamp 0
transform -1 0 1830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9709_
timestamp 0
transform -1 0 1690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9710_
timestamp 0
transform -1 0 910 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9711_
timestamp 0
transform -1 0 1050 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9712_
timestamp 0
transform -1 0 2890 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9713_
timestamp 0
transform -1 0 2930 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9714_
timestamp 0
transform -1 0 290 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9715_
timestamp 0
transform -1 0 290 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9716_
timestamp 0
transform -1 0 2350 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9717_
timestamp 0
transform 1 0 2010 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9718_
timestamp 0
transform -1 0 1890 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9719_
timestamp 0
transform -1 0 3370 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9720_
timestamp 0
transform 1 0 3590 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9721_
timestamp 0
transform 1 0 3450 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9722_
timestamp 0
transform 1 0 2330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9723_
timestamp 0
transform 1 0 2190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9724_
timestamp 0
transform -1 0 3030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9725_
timestamp 0
transform -1 0 3170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9726_
timestamp 0
transform 1 0 2990 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9727_
timestamp 0
transform -1 0 3410 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9728_
timestamp 0
transform -1 0 2110 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9729_
timestamp 0
transform -1 0 2450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9730_
timestamp 0
transform 1 0 2190 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9731_
timestamp 0
transform 1 0 2050 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9732_
timestamp 0
transform -1 0 2830 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9733_
timestamp 0
transform -1 0 3230 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9734_
timestamp 0
transform -1 0 2490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9735_
timestamp 0
transform 1 0 2610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9736_
timestamp 0
transform -1 0 830 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9737_
timestamp 0
transform -1 0 970 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9738_
timestamp 0
transform -1 0 2270 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9739_
timestamp 0
transform -1 0 2510 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9740_
timestamp 0
transform 1 0 1250 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9741_
timestamp 0
transform 1 0 1090 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9742_
timestamp 0
transform -1 0 1830 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9743_
timestamp 0
transform 1 0 1650 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9744_
timestamp 0
transform -1 0 1830 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9745_
timestamp 0
transform 1 0 1270 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9746_
timestamp 0
transform 1 0 2090 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9747_
timestamp 0
transform -1 0 2270 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9748_
timestamp 0
transform -1 0 2310 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9749_
timestamp 0
transform 1 0 2150 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9750_
timestamp 0
transform 1 0 2590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9751_
timestamp 0
transform 1 0 2430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9752_
timestamp 0
transform -1 0 2570 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9753_
timestamp 0
transform -1 0 2690 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9754_
timestamp 0
transform 1 0 3110 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9755_
timestamp 0
transform 1 0 2950 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9756_
timestamp 0
transform 1 0 1310 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9757_
timestamp 0
transform -1 0 1710 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9758_
timestamp 0
transform -1 0 1030 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9759_
timestamp 0
transform -1 0 1190 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9760_
timestamp 0
transform 1 0 1810 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9761_
timestamp 0
transform 1 0 1670 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9762_
timestamp 0
transform 1 0 1130 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9763_
timestamp 0
transform -1 0 990 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9844_
timestamp 0
transform 1 0 9470 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9845_
timestamp 0
transform 1 0 9810 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9846_
timestamp 0
transform 1 0 11250 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9847_
timestamp 0
transform 1 0 9930 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9848_
timestamp 0
transform 1 0 11670 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__9849_
timestamp 0
transform 1 0 11850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9850_
timestamp 0
transform -1 0 10790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9851_
timestamp 0
transform -1 0 10990 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9852_
timestamp 0
transform 1 0 10510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9853_
timestamp 0
transform 1 0 10630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9854_
timestamp 0
transform -1 0 10670 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9855_
timestamp 0
transform -1 0 10850 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9856_
timestamp 0
transform -1 0 9790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9857_
timestamp 0
transform 1 0 9850 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9858_
timestamp 0
transform -1 0 9050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9859_
timestamp 0
transform 1 0 11670 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__9860_
timestamp 0
transform -1 0 11810 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__9861_
timestamp 0
transform -1 0 11550 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__9862_
timestamp 0
transform -1 0 10450 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__9863_
timestamp 0
transform 1 0 9850 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9864_
timestamp 0
transform -1 0 10390 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__9865_
timestamp 0
transform -1 0 10230 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__9866_
timestamp 0
transform 1 0 9410 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9867_
timestamp 0
transform -1 0 9270 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__9868_
timestamp 0
transform -1 0 14150 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9869_
timestamp 0
transform -1 0 12590 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9870_
timestamp 0
transform -1 0 12590 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9871_
timestamp 0
transform -1 0 13630 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9872_
timestamp 0
transform -1 0 12870 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9873_
timestamp 0
transform 1 0 12710 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9874_
timestamp 0
transform -1 0 12430 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9875_
timestamp 0
transform -1 0 12190 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9876_
timestamp 0
transform -1 0 12170 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9877_
timestamp 0
transform -1 0 13210 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__9878_
timestamp 0
transform -1 0 12910 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__9879_
timestamp 0
transform -1 0 13070 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__9880_
timestamp 0
transform -1 0 12990 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__9881_
timestamp 0
transform -1 0 12890 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9882_
timestamp 0
transform 1 0 12730 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__9883_
timestamp 0
transform -1 0 12750 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__9884_
timestamp 0
transform 1 0 12330 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9885_
timestamp 0
transform 1 0 12590 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__9886_
timestamp 0
transform 1 0 13570 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__9887_
timestamp 0
transform -1 0 12230 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9888_
timestamp 0
transform -1 0 12170 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9889_
timestamp 0
transform 1 0 12310 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__9890_
timestamp 0
transform -1 0 11230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9891_
timestamp 0
transform -1 0 11370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9892_
timestamp 0
transform -1 0 11090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9893_
timestamp 0
transform -1 0 10890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9894_
timestamp 0
transform -1 0 10770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9895_
timestamp 0
transform 1 0 11870 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9896_
timestamp 0
transform -1 0 11590 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9897_
timestamp 0
transform -1 0 11710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9898_
timestamp 0
transform 1 0 11270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9899_
timestamp 0
transform -1 0 11450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9900_
timestamp 0
transform 1 0 10430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9901_
timestamp 0
transform -1 0 10310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9902_
timestamp 0
transform -1 0 12510 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9903_
timestamp 0
transform 1 0 12930 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9904_
timestamp 0
transform 1 0 15010 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9905_
timestamp 0
transform 1 0 15510 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9906_
timestamp 0
transform 1 0 15010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9907_
timestamp 0
transform -1 0 14750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9908_
timestamp 0
transform -1 0 14890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__9909_
timestamp 0
transform -1 0 13350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9910_
timestamp 0
transform -1 0 14150 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9911_
timestamp 0
transform 1 0 13990 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9912_
timestamp 0
transform -1 0 13970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9913_
timestamp 0
transform -1 0 13390 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9914_
timestamp 0
transform -1 0 13110 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9915_
timestamp 0
transform -1 0 13250 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9916_
timestamp 0
transform -1 0 12570 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9917_
timestamp 0
transform 1 0 13790 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9918_
timestamp 0
transform 1 0 13650 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9919_
timestamp 0
transform 1 0 13470 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9920_
timestamp 0
transform -1 0 13490 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9921_
timestamp 0
transform 1 0 12550 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9922_
timestamp 0
transform 1 0 13030 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9923_
timestamp 0
transform -1 0 12850 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9924_
timestamp 0
transform 1 0 12630 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9925_
timestamp 0
transform -1 0 12330 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__9926_
timestamp 0
transform -1 0 12370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9927_
timestamp 0
transform 1 0 12690 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9928_
timestamp 0
transform 1 0 12690 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9929_
timestamp 0
transform -1 0 10930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9930_
timestamp 0
transform -1 0 12210 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9931_
timestamp 0
transform -1 0 13910 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9932_
timestamp 0
transform 1 0 14310 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9933_
timestamp 0
transform 1 0 13690 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9934_
timestamp 0
transform -1 0 14410 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9935_
timestamp 0
transform -1 0 11590 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9936_
timestamp 0
transform -1 0 12790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9937_
timestamp 0
transform 1 0 13050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9938_
timestamp 0
transform 1 0 12610 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9939_
timestamp 0
transform -1 0 13930 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9940_
timestamp 0
transform -1 0 12910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9941_
timestamp 0
transform 1 0 13190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9942_
timestamp 0
transform 1 0 13790 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__9943_
timestamp 0
transform 1 0 14830 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9944_
timestamp 0
transform 1 0 15790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__9945_
timestamp 0
transform -1 0 15930 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9946_
timestamp 0
transform 1 0 15770 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__9947_
timestamp 0
transform -1 0 13750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__9948_
timestamp 0
transform 1 0 14450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9949_
timestamp 0
transform 1 0 14310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9950_
timestamp 0
transform -1 0 14150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9951_
timestamp 0
transform -1 0 13590 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9952_
timestamp 0
transform 1 0 13810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9953_
timestamp 0
transform 1 0 13670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__9954_
timestamp 0
transform -1 0 13690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9955_
timestamp 0
transform -1 0 13090 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9956_
timestamp 0
transform -1 0 13230 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9957_
timestamp 0
transform -1 0 13530 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9958_
timestamp 0
transform -1 0 13370 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9959_
timestamp 0
transform 1 0 13210 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9960_
timestamp 0
transform 1 0 14470 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9961_
timestamp 0
transform 1 0 13870 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9962_
timestamp 0
transform -1 0 14650 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9963_
timestamp 0
transform 1 0 14310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9964_
timestamp 0
transform 1 0 14130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9965_
timestamp 0
transform 1 0 14470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9966_
timestamp 0
transform 1 0 14630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__9967_
timestamp 0
transform 1 0 13810 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9968_
timestamp 0
transform 1 0 13670 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9969_
timestamp 0
transform -1 0 13610 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9970_
timestamp 0
transform 1 0 13530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9971_
timestamp 0
transform -1 0 13450 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9972_
timestamp 0
transform 1 0 13150 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9973_
timestamp 0
transform -1 0 13310 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9974_
timestamp 0
transform 1 0 13290 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9975_
timestamp 0
transform 1 0 12310 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9976_
timestamp 0
transform 1 0 7710 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__9977_
timestamp 0
transform -1 0 8210 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__9978_
timestamp 0
transform 1 0 7670 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__9979_
timestamp 0
transform 1 0 12850 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__9980_
timestamp 0
transform 1 0 13710 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9981_
timestamp 0
transform -1 0 15350 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__9982_
timestamp 0
transform 1 0 15170 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9983_
timestamp 0
transform 1 0 14210 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9984_
timestamp 0
transform -1 0 13910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__9985_
timestamp 0
transform 1 0 14050 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9986_
timestamp 0
transform -1 0 14570 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__9987_
timestamp 0
transform -1 0 14190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9988_
timestamp 0
transform 1 0 14150 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9989_
timestamp 0
transform -1 0 14090 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9990_
timestamp 0
transform 1 0 13370 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9991_
timestamp 0
transform -1 0 13970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__9992_
timestamp 0
transform -1 0 13870 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9993_
timestamp 0
transform 1 0 13990 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__9994_
timestamp 0
transform 1 0 14590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9995_
timestamp 0
transform -1 0 14150 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9996_
timestamp 0
transform 1 0 14010 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9997_
timestamp 0
transform -1 0 13910 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9998_
timestamp 0
transform -1 0 14310 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__9999_
timestamp 0
transform -1 0 13770 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10000_
timestamp 0
transform 1 0 13290 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10001_
timestamp 0
transform -1 0 13610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10002_
timestamp 0
transform -1 0 13470 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10003_
timestamp 0
transform -1 0 13230 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10004_
timestamp 0
transform 1 0 13730 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10005_
timestamp 0
transform 1 0 14430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10006_
timestamp 0
transform -1 0 14150 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10007_
timestamp 0
transform -1 0 14610 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10008_
timestamp 0
transform 1 0 14310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10009_
timestamp 0
transform 1 0 16190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10010_
timestamp 0
transform 1 0 16430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10011_
timestamp 0
transform 1 0 16290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10012_
timestamp 0
transform -1 0 15230 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10013_
timestamp 0
transform -1 0 15710 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10014_
timestamp 0
transform -1 0 14730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10015_
timestamp 0
transform 1 0 14450 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10016_
timestamp 0
transform 1 0 14150 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10017_
timestamp 0
transform -1 0 15510 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10018_
timestamp 0
transform 1 0 14810 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10019_
timestamp 0
transform -1 0 14310 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10020_
timestamp 0
transform -1 0 14710 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10021_
timestamp 0
transform 1 0 14390 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10022_
timestamp 0
transform -1 0 14710 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10023_
timestamp 0
transform 1 0 14850 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10024_
timestamp 0
transform -1 0 14390 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10025_
timestamp 0
transform -1 0 14250 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10026_
timestamp 0
transform -1 0 14010 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10027_
timestamp 0
transform -1 0 13850 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10028_
timestamp 0
transform 1 0 13570 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10029_
timestamp 0
transform 1 0 14470 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10030_
timestamp 0
transform 1 0 14950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10031_
timestamp 0
transform 1 0 16790 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10032_
timestamp 0
transform -1 0 15170 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__10033_
timestamp 0
transform 1 0 16870 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10034_
timestamp 0
transform -1 0 16030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10035_
timestamp 0
transform -1 0 16170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10036_
timestamp 0
transform -1 0 14690 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10037_
timestamp 0
transform -1 0 14830 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10038_
timestamp 0
transform 1 0 15210 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10039_
timestamp 0
transform -1 0 14930 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10040_
timestamp 0
transform 1 0 15070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10041_
timestamp 0
transform 1 0 15090 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10042_
timestamp 0
transform 1 0 14950 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10043_
timestamp 0
transform -1 0 15010 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10044_
timestamp 0
transform -1 0 14630 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10045_
timestamp 0
transform -1 0 14490 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10046_
timestamp 0
transform 1 0 14750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10047_
timestamp 0
transform -1 0 14650 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10048_
timestamp 0
transform -1 0 14810 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10049_
timestamp 0
transform -1 0 14670 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10050_
timestamp 0
transform 1 0 13970 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10051_
timestamp 0
transform 1 0 14950 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10052_
timestamp 0
transform 1 0 15550 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10053_
timestamp 0
transform 1 0 14530 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10054_
timestamp 0
transform 1 0 16370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10055_
timestamp 0
transform -1 0 16310 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10056_
timestamp 0
transform 1 0 15990 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10057_
timestamp 0
transform -1 0 15790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10058_
timestamp 0
transform -1 0 15790 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10059_
timestamp 0
transform -1 0 15390 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10060_
timestamp 0
transform 1 0 15310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10061_
timestamp 0
transform 1 0 15690 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10062_
timestamp 0
transform -1 0 15570 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10063_
timestamp 0
transform -1 0 15430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10064_
timestamp 0
transform -1 0 15290 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10065_
timestamp 0
transform 1 0 15310 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10066_
timestamp 0
transform 1 0 15250 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10067_
timestamp 0
transform -1 0 14870 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__10068_
timestamp 0
transform 1 0 14970 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10069_
timestamp 0
transform -1 0 14850 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10070_
timestamp 0
transform 1 0 13010 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10071_
timestamp 0
transform 1 0 14430 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10072_
timestamp 0
transform -1 0 15590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10073_
timestamp 0
transform 1 0 15230 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10074_
timestamp 0
transform -1 0 16170 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10075_
timestamp 0
transform -1 0 15950 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10076_
timestamp 0
transform -1 0 16090 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10077_
timestamp 0
transform 1 0 15670 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10078_
timestamp 0
transform 1 0 15950 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10079_
timestamp 0
transform 1 0 15510 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10080_
timestamp 0
transform 1 0 15830 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10081_
timestamp 0
transform -1 0 15710 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10082_
timestamp 0
transform 1 0 16050 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10083_
timestamp 0
transform -1 0 16010 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10084_
timestamp 0
transform 1 0 16110 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10085_
timestamp 0
transform -1 0 15630 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10086_
timestamp 0
transform 1 0 15130 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10087_
timestamp 0
transform -1 0 15050 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10088_
timestamp 0
transform 1 0 14890 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10089_
timestamp 0
transform -1 0 15130 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10090_
timestamp 0
transform -1 0 15290 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10091_
timestamp 0
transform -1 0 15130 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10092_
timestamp 0
transform 1 0 14530 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10093_
timestamp 0
transform -1 0 13190 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10094_
timestamp 0
transform 1 0 15830 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10095_
timestamp 0
transform 1 0 14750 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10096_
timestamp 0
transform 1 0 15430 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10097_
timestamp 0
transform 1 0 15170 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10098_
timestamp 0
transform 1 0 15590 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10099_
timestamp 0
transform -1 0 15770 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10100_
timestamp 0
transform 1 0 15890 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10101_
timestamp 0
transform 1 0 15790 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10102_
timestamp 0
transform 1 0 16490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10103_
timestamp 0
transform 1 0 16490 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10104_
timestamp 0
transform 1 0 16630 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10105_
timestamp 0
transform 1 0 16210 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10106_
timestamp 0
transform -1 0 16290 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10107_
timestamp 0
transform -1 0 16090 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10108_
timestamp 0
transform 1 0 16210 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10109_
timestamp 0
transform 1 0 16150 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10110_
timestamp 0
transform -1 0 16010 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10111_
timestamp 0
transform -1 0 16130 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10112_
timestamp 0
transform 1 0 16250 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10113_
timestamp 0
transform 1 0 15950 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10114_
timestamp 0
transform 1 0 15870 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10115_
timestamp 0
transform -1 0 15510 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10116_
timestamp 0
transform 1 0 15370 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10117_
timestamp 0
transform 1 0 15550 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10118_
timestamp 0
transform -1 0 15430 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10119_
timestamp 0
transform 1 0 13470 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10120_
timestamp 0
transform 1 0 13670 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10121_
timestamp 0
transform -1 0 14710 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10122_
timestamp 0
transform 1 0 13510 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10123_
timestamp 0
transform 1 0 13890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__10124_
timestamp 0
transform 1 0 15990 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10125_
timestamp 0
transform 1 0 15710 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10126_
timestamp 0
transform 1 0 15850 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10127_
timestamp 0
transform 1 0 16490 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10128_
timestamp 0
transform 1 0 16370 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10129_
timestamp 0
transform 1 0 16450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10130_
timestamp 0
transform -1 0 16790 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10131_
timestamp 0
transform -1 0 16530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10132_
timestamp 0
transform -1 0 16930 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10133_
timestamp 0
transform 1 0 16770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10134_
timestamp 0
transform 1 0 16610 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10135_
timestamp 0
transform 1 0 16910 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10136_
timestamp 0
transform -1 0 16650 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10137_
timestamp 0
transform -1 0 16850 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10138_
timestamp 0
transform 1 0 16610 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10139_
timestamp 0
transform -1 0 16450 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10140_
timestamp 0
transform -1 0 16150 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10141_
timestamp 0
transform -1 0 16290 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10142_
timestamp 0
transform 1 0 14030 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10143_
timestamp 0
transform -1 0 15910 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10144_
timestamp 0
transform -1 0 16030 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10145_
timestamp 0
transform 1 0 15730 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10146_
timestamp 0
transform 1 0 15990 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10147_
timestamp 0
transform 1 0 16150 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10148_
timestamp 0
transform 1 0 16570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10149_
timestamp 0
transform -1 0 16450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10150_
timestamp 0
transform -1 0 16470 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__10151_
timestamp 0
transform 1 0 16430 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10152_
timestamp 0
transform 1 0 17030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10153_
timestamp 0
transform 1 0 16610 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10154_
timestamp 0
transform 1 0 16970 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10155_
timestamp 0
transform 1 0 16930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10156_
timestamp 0
transform 1 0 16770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10157_
timestamp 0
transform 1 0 17050 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10158_
timestamp 0
transform 1 0 16230 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__10159_
timestamp 0
transform 1 0 16670 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10160_
timestamp 0
transform 1 0 16810 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10161_
timestamp 0
transform -1 0 16710 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10162_
timestamp 0
transform -1 0 16330 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10163_
timestamp 0
transform -1 0 16290 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10164_
timestamp 0
transform -1 0 16190 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10165_
timestamp 0
transform 1 0 13310 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10166_
timestamp 0
transform 1 0 16810 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10167_
timestamp 0
transform 1 0 16350 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10168_
timestamp 0
transform -1 0 17050 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10169_
timestamp 0
transform 1 0 15710 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__10170_
timestamp 0
transform -1 0 16890 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10171_
timestamp 0
transform -1 0 16930 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10172_
timestamp 0
transform 1 0 16730 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10173_
timestamp 0
transform -1 0 16110 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__10174_
timestamp 0
transform 1 0 17010 0 1 250
box -6 -8 26 248
use FILL  FILL_1__10175_
timestamp 0
transform -1 0 17090 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__10176_
timestamp 0
transform -1 0 17050 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10177_
timestamp 0
transform 1 0 16950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10178_
timestamp 0
transform -1 0 16830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10179_
timestamp 0
transform 1 0 17030 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10180_
timestamp 0
transform -1 0 17050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10181_
timestamp 0
transform 1 0 16990 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10182_
timestamp 0
transform 1 0 16450 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10183_
timestamp 0
transform -1 0 16910 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10184_
timestamp 0
transform -1 0 17010 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10185_
timestamp 0
transform -1 0 16770 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10186_
timestamp 0
transform 1 0 16590 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10187_
timestamp 0
transform -1 0 16450 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10188_
timestamp 0
transform -1 0 16310 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10189_
timestamp 0
transform 1 0 14470 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10190_
timestamp 0
transform -1 0 12110 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10191_
timestamp 0
transform -1 0 16890 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10192_
timestamp 0
transform 1 0 17050 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10193_
timestamp 0
transform 1 0 16810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10194_
timestamp 0
transform -1 0 16930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10195_
timestamp 0
transform 1 0 17050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10196_
timestamp 0
transform 1 0 16730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10197_
timestamp 0
transform 1 0 15290 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__10198_
timestamp 0
transform -1 0 16870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10199_
timestamp 0
transform 1 0 16970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10200_
timestamp 0
transform 1 0 17090 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10201_
timestamp 0
transform -1 0 16870 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10202_
timestamp 0
transform 1 0 16730 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10203_
timestamp 0
transform -1 0 16710 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10204_
timestamp 0
transform -1 0 16570 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10205_
timestamp 0
transform 1 0 12450 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10206_
timestamp 0
transform -1 0 11570 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10207_
timestamp 0
transform 1 0 14290 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10208_
timestamp 0
transform 1 0 14530 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10209_
timestamp 0
transform 1 0 14390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10210_
timestamp 0
transform 1 0 14150 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10211_
timestamp 0
transform -1 0 12790 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10212_
timestamp 0
transform -1 0 12530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10213_
timestamp 0
transform -1 0 13050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10214_
timestamp 0
transform -1 0 14030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10215_
timestamp 0
transform 1 0 15750 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10216_
timestamp 0
transform 1 0 15650 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10217_
timestamp 0
transform 1 0 15490 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10218_
timestamp 0
transform 1 0 15330 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10219_
timestamp 0
transform 1 0 15370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10220_
timestamp 0
transform 1 0 15370 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10221_
timestamp 0
transform 1 0 14930 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10222_
timestamp 0
transform 1 0 12970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10223_
timestamp 0
transform -1 0 15250 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10224_
timestamp 0
transform 1 0 15650 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10225_
timestamp 0
transform 1 0 15350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10226_
timestamp 0
transform -1 0 15110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10227_
timestamp 0
transform 1 0 13230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10228_
timestamp 0
transform -1 0 11950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10229_
timestamp 0
transform 1 0 10810 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10230_
timestamp 0
transform 1 0 13110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10231_
timestamp 0
transform -1 0 14870 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10232_
timestamp 0
transform 1 0 14690 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10233_
timestamp 0
transform -1 0 14190 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10234_
timestamp 0
transform -1 0 14310 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10235_
timestamp 0
transform 1 0 14930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10236_
timestamp 0
transform -1 0 15530 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10237_
timestamp 0
transform -1 0 15810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10238_
timestamp 0
transform -1 0 15950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10239_
timestamp 0
transform 1 0 15930 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10240_
timestamp 0
transform -1 0 15650 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10241_
timestamp 0
transform 1 0 15610 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10242_
timestamp 0
transform -1 0 15730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10243_
timestamp 0
transform -1 0 15810 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10244_
timestamp 0
transform -1 0 15650 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10245_
timestamp 0
transform -1 0 14270 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10246_
timestamp 0
transform -1 0 15550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10247_
timestamp 0
transform 1 0 15090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10248_
timestamp 0
transform 1 0 14570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10249_
timestamp 0
transform -1 0 12770 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10250_
timestamp 0
transform -1 0 12370 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10251_
timestamp 0
transform -1 0 12930 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10252_
timestamp 0
transform 1 0 12450 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10253_
timestamp 0
transform 1 0 12670 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10254_
timestamp 0
transform 1 0 12810 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10255_
timestamp 0
transform 1 0 12950 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10256_
timestamp 0
transform -1 0 10970 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10257_
timestamp 0
transform -1 0 11070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10258_
timestamp 0
transform 1 0 12590 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10259_
timestamp 0
transform 1 0 14530 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10260_
timestamp 0
transform 1 0 16310 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10261_
timestamp 0
transform 1 0 16170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10262_
timestamp 0
transform -1 0 16110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10263_
timestamp 0
transform 1 0 16210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10264_
timestamp 0
transform -1 0 14730 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10265_
timestamp 0
transform -1 0 14950 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10266_
timestamp 0
transform 1 0 14810 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10267_
timestamp 0
transform -1 0 15250 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10268_
timestamp 0
transform -1 0 14530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10269_
timestamp 0
transform 1 0 14390 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10270_
timestamp 0
transform 1 0 15070 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10271_
timestamp 0
transform -1 0 14670 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10272_
timestamp 0
transform -1 0 13430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10273_
timestamp 0
transform 1 0 13170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10274_
timestamp 0
transform -1 0 13290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10275_
timestamp 0
transform 1 0 13030 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10276_
timestamp 0
transform -1 0 12230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10277_
timestamp 0
transform 1 0 12210 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10278_
timestamp 0
transform -1 0 12090 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10279_
timestamp 0
transform -1 0 11430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10280_
timestamp 0
transform 1 0 12870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10281_
timestamp 0
transform -1 0 12870 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10282_
timestamp 0
transform 1 0 16670 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10283_
timestamp 0
transform 1 0 16530 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10284_
timestamp 0
transform 1 0 16050 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10285_
timestamp 0
transform 1 0 15730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10286_
timestamp 0
transform 1 0 14810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10287_
timestamp 0
transform -1 0 14970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10288_
timestamp 0
transform 1 0 14830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10289_
timestamp 0
transform 1 0 14770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10290_
timestamp 0
transform -1 0 14390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10291_
timestamp 0
transform -1 0 14110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10292_
timestamp 0
transform -1 0 14650 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10293_
timestamp 0
transform -1 0 13470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10294_
timestamp 0
transform -1 0 12790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10295_
timestamp 0
transform 1 0 13590 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10296_
timestamp 0
transform -1 0 12650 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10297_
timestamp 0
transform -1 0 12610 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10298_
timestamp 0
transform -1 0 12750 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10299_
timestamp 0
transform -1 0 12470 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10300_
timestamp 0
transform 1 0 11990 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10301_
timestamp 0
transform 1 0 12890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10302_
timestamp 0
transform -1 0 16950 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10303_
timestamp 0
transform 1 0 16770 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10304_
timestamp 0
transform 1 0 16370 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10305_
timestamp 0
transform 1 0 16230 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10306_
timestamp 0
transform 1 0 15470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10307_
timestamp 0
transform 1 0 15330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10308_
timestamp 0
transform -1 0 15350 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10309_
timestamp 0
transform 1 0 14790 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10310_
timestamp 0
transform -1 0 14830 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10311_
timestamp 0
transform -1 0 14510 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10312_
timestamp 0
transform 1 0 14950 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10313_
timestamp 0
transform 1 0 15390 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10314_
timestamp 0
transform -1 0 14370 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10315_
timestamp 0
transform -1 0 14670 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10316_
timestamp 0
transform 1 0 15070 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10317_
timestamp 0
transform -1 0 13810 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10318_
timestamp 0
transform -1 0 13510 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10319_
timestamp 0
transform -1 0 13230 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10320_
timestamp 0
transform -1 0 13370 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10321_
timestamp 0
transform -1 0 13110 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10322_
timestamp 0
transform 1 0 12410 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10323_
timestamp 0
transform 1 0 12210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10324_
timestamp 0
transform 1 0 13770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10325_
timestamp 0
transform 1 0 15810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10326_
timestamp 0
transform -1 0 16030 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10327_
timestamp 0
transform 1 0 16130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10328_
timestamp 0
transform 1 0 15830 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10329_
timestamp 0
transform -1 0 15970 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10330_
timestamp 0
transform -1 0 16110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10331_
timestamp 0
transform -1 0 15970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10332_
timestamp 0
transform 1 0 14930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10333_
timestamp 0
transform 1 0 15070 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10334_
timestamp 0
transform 1 0 15670 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10335_
timestamp 0
transform 1 0 15550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10336_
timestamp 0
transform -1 0 15130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10337_
timestamp 0
transform -1 0 14630 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10338_
timestamp 0
transform 1 0 15250 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10339_
timestamp 0
transform -1 0 13930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10340_
timestamp 0
transform 1 0 13650 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10341_
timestamp 0
transform -1 0 13510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10342_
timestamp 0
transform -1 0 13370 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10343_
timestamp 0
transform 1 0 12310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10344_
timestamp 0
transform 1 0 11350 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10345_
timestamp 0
transform -1 0 15690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10346_
timestamp 0
transform 1 0 16290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10347_
timestamp 0
transform 1 0 16490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10348_
timestamp 0
transform 1 0 16350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10349_
timestamp 0
transform 1 0 15150 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10350_
timestamp 0
transform -1 0 15470 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10351_
timestamp 0
transform 1 0 15590 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10352_
timestamp 0
transform 1 0 15310 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10353_
timestamp 0
transform 1 0 15010 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10354_
timestamp 0
transform 1 0 14750 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10355_
timestamp 0
transform -1 0 14890 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10356_
timestamp 0
transform -1 0 14490 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10357_
timestamp 0
transform 1 0 13930 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10358_
timestamp 0
transform 1 0 14210 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10359_
timestamp 0
transform 1 0 14070 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10360_
timestamp 0
transform -1 0 14210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10361_
timestamp 0
transform -1 0 14230 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10362_
timestamp 0
transform -1 0 14630 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10363_
timestamp 0
transform -1 0 13650 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10364_
timestamp 0
transform 1 0 14050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10365_
timestamp 0
transform 1 0 14450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10366_
timestamp 0
transform 1 0 14310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10367_
timestamp 0
transform -1 0 14370 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10368_
timestamp 0
transform -1 0 13850 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10369_
timestamp 0
transform 1 0 12910 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10370_
timestamp 0
transform 1 0 11470 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10371_
timestamp 0
transform 1 0 12810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10372_
timestamp 0
transform -1 0 14010 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10373_
timestamp 0
transform 1 0 15230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10374_
timestamp 0
transform 1 0 16330 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10375_
timestamp 0
transform 1 0 16450 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10376_
timestamp 0
transform 1 0 16210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10377_
timestamp 0
transform -1 0 14850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10378_
timestamp 0
transform -1 0 15150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10379_
timestamp 0
transform 1 0 15450 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10380_
timestamp 0
transform -1 0 15010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10381_
timestamp 0
transform -1 0 14710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10382_
timestamp 0
transform 1 0 15490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10383_
timestamp 0
transform 1 0 15490 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__10384_
timestamp 0
transform -1 0 15630 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__10385_
timestamp 0
transform 1 0 15210 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__10386_
timestamp 0
transform 1 0 13430 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10387_
timestamp 0
transform -1 0 13310 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10388_
timestamp 0
transform -1 0 13210 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10389_
timestamp 0
transform -1 0 13050 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10390_
timestamp 0
transform 1 0 12910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10391_
timestamp 0
transform 1 0 14550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10392_
timestamp 0
transform -1 0 14290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10393_
timestamp 0
transform 1 0 14410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10394_
timestamp 0
transform 1 0 16130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__10395_
timestamp 0
transform -1 0 15370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10396_
timestamp 0
transform -1 0 16230 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10397_
timestamp 0
transform 1 0 16270 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10398_
timestamp 0
transform 1 0 16590 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__10399_
timestamp 0
transform -1 0 16550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__10400_
timestamp 0
transform 1 0 15650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10401_
timestamp 0
transform -1 0 16270 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__10402_
timestamp 0
transform 1 0 16390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__10403_
timestamp 0
transform -1 0 16710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__10404_
timestamp 0
transform 1 0 16190 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__10405_
timestamp 0
transform -1 0 16070 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__10406_
timestamp 0
transform -1 0 14130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10407_
timestamp 0
transform -1 0 14130 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10408_
timestamp 0
transform -1 0 15350 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__10409_
timestamp 0
transform -1 0 13730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10410_
timestamp 0
transform 1 0 13670 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10411_
timestamp 0
transform 1 0 12770 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10412_
timestamp 0
transform -1 0 13870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10413_
timestamp 0
transform -1 0 13990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10414_
timestamp 0
transform 1 0 16970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10415_
timestamp 0
transform 1 0 16910 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__10416_
timestamp 0
transform -1 0 16870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__10417_
timestamp 0
transform 1 0 16990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__10418_
timestamp 0
transform 1 0 15410 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__10419_
timestamp 0
transform 1 0 16930 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__10420_
timestamp 0
transform 1 0 16930 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__10421_
timestamp 0
transform 1 0 16690 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__10422_
timestamp 0
transform -1 0 16090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10423_
timestamp 0
transform -1 0 13330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10424_
timestamp 0
transform -1 0 13190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10425_
timestamp 0
transform -1 0 13030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10426_
timestamp 0
transform 1 0 13070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10427_
timestamp 0
transform 1 0 16810 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__10428_
timestamp 0
transform -1 0 15950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10429_
timestamp 0
transform -1 0 16330 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__10430_
timestamp 0
transform -1 0 16450 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__10431_
timestamp 0
transform 1 0 15790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10432_
timestamp 0
transform -1 0 16330 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__10433_
timestamp 0
transform 1 0 16390 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__10434_
timestamp 0
transform 1 0 16570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10435_
timestamp 0
transform -1 0 16910 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10436_
timestamp 0
transform 1 0 16850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10437_
timestamp 0
transform -1 0 16750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10438_
timestamp 0
transform -1 0 16670 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10439_
timestamp 0
transform 1 0 17030 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10440_
timestamp 0
transform -1 0 17050 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__10441_
timestamp 0
transform -1 0 16910 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10442_
timestamp 0
transform 1 0 16510 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10443_
timestamp 0
transform 1 0 15970 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10444_
timestamp 0
transform -1 0 15850 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10445_
timestamp 0
transform -1 0 15730 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10446_
timestamp 0
transform 1 0 13170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__10447_
timestamp 0
transform 1 0 12090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10448_
timestamp 0
transform 1 0 16410 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10449_
timestamp 0
transform 1 0 16110 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__10450_
timestamp 0
transform 1 0 16690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10451_
timestamp 0
transform 1 0 16630 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10452_
timestamp 0
transform 1 0 16590 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10453_
timestamp 0
transform 1 0 16490 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10454_
timestamp 0
transform -1 0 13210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10455_
timestamp 0
transform -1 0 13070 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10456_
timestamp 0
transform -1 0 12490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10457_
timestamp 0
transform 1 0 11170 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10458_
timestamp 0
transform -1 0 9410 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10459_
timestamp 0
transform -1 0 9310 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10460_
timestamp 0
transform 1 0 9690 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10461_
timestamp 0
transform 1 0 9550 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10462_
timestamp 0
transform 1 0 9730 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10463_
timestamp 0
transform 1 0 9970 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10464_
timestamp 0
transform 1 0 9830 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10465_
timestamp 0
transform 1 0 9270 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10466_
timestamp 0
transform -1 0 9130 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10467_
timestamp 0
transform 1 0 10590 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10468_
timestamp 0
transform -1 0 9970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10469_
timestamp 0
transform -1 0 9850 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10470_
timestamp 0
transform 1 0 9950 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10471_
timestamp 0
transform -1 0 9830 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10472_
timestamp 0
transform -1 0 8910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10473_
timestamp 0
transform -1 0 8650 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10474_
timestamp 0
transform -1 0 8770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10475_
timestamp 0
transform -1 0 8630 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10476_
timestamp 0
transform -1 0 8790 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10477_
timestamp 0
transform -1 0 8870 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10478_
timestamp 0
transform -1 0 9010 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10479_
timestamp 0
transform 1 0 8890 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10480_
timestamp 0
transform 1 0 8790 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10481_
timestamp 0
transform 1 0 8910 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10482_
timestamp 0
transform -1 0 11110 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10483_
timestamp 0
transform -1 0 10250 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10484_
timestamp 0
transform -1 0 10390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10485_
timestamp 0
transform 1 0 9350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10486_
timestamp 0
transform -1 0 9230 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10487_
timestamp 0
transform 1 0 9070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10488_
timestamp 0
transform -1 0 8990 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10489_
timestamp 0
transform -1 0 8730 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10490_
timestamp 0
transform -1 0 8870 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10491_
timestamp 0
transform 1 0 9750 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10492_
timestamp 0
transform 1 0 9570 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10493_
timestamp 0
transform -1 0 9510 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10494_
timestamp 0
transform 1 0 9870 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10495_
timestamp 0
transform 1 0 10010 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10496_
timestamp 0
transform 1 0 10250 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10497_
timestamp 0
transform 1 0 11310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10498_
timestamp 0
transform -1 0 11190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10499_
timestamp 0
transform 1 0 11010 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10500_
timestamp 0
transform -1 0 11050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10501_
timestamp 0
transform 1 0 10490 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10502_
timestamp 0
transform 1 0 10370 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10503_
timestamp 0
transform -1 0 9630 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10504_
timestamp 0
transform -1 0 9490 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10505_
timestamp 0
transform -1 0 9190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10506_
timestamp 0
transform 1 0 9310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10507_
timestamp 0
transform 1 0 9610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10508_
timestamp 0
transform 1 0 10990 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__10509_
timestamp 0
transform -1 0 10590 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10510_
timestamp 0
transform -1 0 10890 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10511_
timestamp 0
transform 1 0 10710 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10512_
timestamp 0
transform 1 0 10110 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10513_
timestamp 0
transform 1 0 10490 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10514_
timestamp 0
transform -1 0 10390 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10515_
timestamp 0
transform 1 0 10450 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__10516_
timestamp 0
transform 1 0 10110 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10517_
timestamp 0
transform 1 0 10710 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__10518_
timestamp 0
transform 1 0 10970 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__10519_
timestamp 0
transform -1 0 10870 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__10520_
timestamp 0
transform -1 0 10830 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__10521_
timestamp 0
transform -1 0 11190 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10522_
timestamp 0
transform -1 0 12910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10523_
timestamp 0
transform 1 0 13130 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10524_
timestamp 0
transform -1 0 13010 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10525_
timestamp 0
transform -1 0 12870 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10526_
timestamp 0
transform -1 0 10950 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10527_
timestamp 0
transform -1 0 11090 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10528_
timestamp 0
transform -1 0 10830 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10529_
timestamp 0
transform -1 0 10570 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10530_
timestamp 0
transform 1 0 10970 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__10531_
timestamp 0
transform 1 0 10850 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__10532_
timestamp 0
transform 1 0 10710 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__10533_
timestamp 0
transform 1 0 10550 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__10534_
timestamp 0
transform -1 0 9470 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10535_
timestamp 0
transform 1 0 10590 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__10536_
timestamp 0
transform -1 0 10710 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__10537_
timestamp 0
transform 1 0 10650 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10538_
timestamp 0
transform 1 0 10350 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__10539_
timestamp 0
transform -1 0 10550 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__10540_
timestamp 0
transform -1 0 11450 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10541_
timestamp 0
transform 1 0 10910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10542_
timestamp 0
transform -1 0 10510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10543_
timestamp 0
transform -1 0 10790 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10544_
timestamp 0
transform -1 0 10650 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10545_
timestamp 0
transform 1 0 10850 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10546_
timestamp 0
transform 1 0 10970 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10547_
timestamp 0
transform 1 0 10450 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10548_
timestamp 0
transform -1 0 10130 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__10549_
timestamp 0
transform -1 0 9870 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__10550_
timestamp 0
transform -1 0 10010 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__10551_
timestamp 0
transform 1 0 9710 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10552_
timestamp 0
transform -1 0 9590 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10553_
timestamp 0
transform -1 0 9270 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10554_
timestamp 0
transform -1 0 9830 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10555_
timestamp 0
transform 1 0 10250 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10556_
timestamp 0
transform 1 0 10710 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10557_
timestamp 0
transform -1 0 10590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10558_
timestamp 0
transform -1 0 10450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10559_
timestamp 0
transform -1 0 10190 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10560_
timestamp 0
transform -1 0 10130 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10561_
timestamp 0
transform 1 0 10290 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10562_
timestamp 0
transform -1 0 10270 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10563_
timestamp 0
transform -1 0 9530 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10564_
timestamp 0
transform -1 0 9690 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10565_
timestamp 0
transform 1 0 9350 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10566_
timestamp 0
transform 1 0 11130 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__10567_
timestamp 0
transform -1 0 11330 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10568_
timestamp 0
transform 1 0 11430 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10569_
timestamp 0
transform -1 0 11430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10570_
timestamp 0
transform -1 0 11130 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10571_
timestamp 0
transform 1 0 11550 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10572_
timestamp 0
transform -1 0 11230 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10573_
timestamp 0
transform 1 0 10090 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10574_
timestamp 0
transform 1 0 9970 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10575_
timestamp 0
transform 1 0 10090 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10576_
timestamp 0
transform -1 0 10430 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10577_
timestamp 0
transform -1 0 10270 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10578_
timestamp 0
transform 1 0 11410 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__10579_
timestamp 0
transform 1 0 11530 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__10580_
timestamp 0
transform 1 0 11650 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__10581_
timestamp 0
transform -1 0 11290 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__10582_
timestamp 0
transform 1 0 11370 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__10583_
timestamp 0
transform 1 0 11510 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10584_
timestamp 0
transform 1 0 11650 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10585_
timestamp 0
transform -1 0 11630 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10586_
timestamp 0
transform -1 0 11370 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__10587_
timestamp 0
transform 1 0 11650 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__10588_
timestamp 0
transform -1 0 11510 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__10589_
timestamp 0
transform -1 0 11810 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__10590_
timestamp 0
transform -1 0 11350 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10591_
timestamp 0
transform -1 0 11490 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10592_
timestamp 0
transform -1 0 11250 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10593_
timestamp 0
transform 1 0 11350 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10594_
timestamp 0
transform -1 0 11870 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10595_
timestamp 0
transform -1 0 12050 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10596_
timestamp 0
transform 1 0 11890 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__10597_
timestamp 0
transform -1 0 11990 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__10598_
timestamp 0
transform 1 0 12470 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__10599_
timestamp 0
transform -1 0 12330 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__10600_
timestamp 0
transform -1 0 12190 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__10601_
timestamp 0
transform -1 0 11950 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__10602_
timestamp 0
transform -1 0 12230 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__10603_
timestamp 0
transform -1 0 12090 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__10604_
timestamp 0
transform 1 0 10450 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10605_
timestamp 0
transform -1 0 11270 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10606_
timestamp 0
transform 1 0 10590 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10607_
timestamp 0
transform 1 0 15210 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10608_
timestamp 0
transform -1 0 16590 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10609_
timestamp 0
transform -1 0 16110 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10610_
timestamp 0
transform 1 0 16730 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__10611_
timestamp 0
transform 1 0 11570 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10612_
timestamp 0
transform 1 0 10730 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10613_
timestamp 0
transform 1 0 11270 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10614_
timestamp 0
transform -1 0 11450 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10615_
timestamp 0
transform -1 0 11190 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10616_
timestamp 0
transform 1 0 10870 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10617_
timestamp 0
transform -1 0 11050 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10618_
timestamp 0
transform -1 0 10630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10619_
timestamp 0
transform -1 0 12770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10620_
timestamp 0
transform 1 0 12590 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10621_
timestamp 0
transform 1 0 11970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__10622_
timestamp 0
transform 1 0 11930 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__10623_
timestamp 0
transform 1 0 10130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10624_
timestamp 0
transform 1 0 13590 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10625_
timestamp 0
transform 1 0 13430 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10626_
timestamp 0
transform -1 0 13730 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10627_
timestamp 0
transform -1 0 13850 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__10628_
timestamp 0
transform 1 0 12410 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10629_
timestamp 0
transform 1 0 12070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10630_
timestamp 0
transform -1 0 12270 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10631_
timestamp 0
transform 1 0 11870 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10632_
timestamp 0
transform 1 0 12450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10633_
timestamp 0
transform -1 0 12610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10634_
timestamp 0
transform -1 0 13410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10635_
timestamp 0
transform 1 0 13510 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10636_
timestamp 0
transform 1 0 16290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10637_
timestamp 0
transform -1 0 16430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__10638_
timestamp 0
transform 1 0 15210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10639_
timestamp 0
transform -1 0 15870 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__10640_
timestamp 0
transform -1 0 11850 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10641_
timestamp 0
transform -1 0 12110 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10642_
timestamp 0
transform 1 0 11930 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10643_
timestamp 0
transform -1 0 11990 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10644_
timestamp 0
transform 1 0 12370 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10645_
timestamp 0
transform 1 0 12230 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10646_
timestamp 0
transform -1 0 12410 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10647_
timestamp 0
transform 1 0 11990 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10648_
timestamp 0
transform -1 0 12950 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10649_
timestamp 0
transform 1 0 12770 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10650_
timestamp 0
transform 1 0 15370 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10651_
timestamp 0
transform 1 0 15210 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10652_
timestamp 0
transform -1 0 15070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10653_
timestamp 0
transform -1 0 15190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10654_
timestamp 0
transform -1 0 11710 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10655_
timestamp 0
transform -1 0 11710 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10656_
timestamp 0
transform 1 0 12210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10657_
timestamp 0
transform 1 0 12070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10658_
timestamp 0
transform -1 0 11870 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10659_
timestamp 0
transform -1 0 12190 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__10660_
timestamp 0
transform -1 0 13370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10661_
timestamp 0
transform -1 0 13410 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10662_
timestamp 0
transform 1 0 11770 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10663_
timestamp 0
transform -1 0 11910 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10664_
timestamp 0
transform 1 0 11690 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10665_
timestamp 0
transform -1 0 11830 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10666_
timestamp 0
transform -1 0 9730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10667_
timestamp 0
transform -1 0 11570 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10668_
timestamp 0
transform 1 0 11150 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10669_
timestamp 0
transform -1 0 10130 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10670_
timestamp 0
transform -1 0 10950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10671_
timestamp 0
transform 1 0 10790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10672_
timestamp 0
transform -1 0 10650 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10673_
timestamp 0
transform -1 0 10770 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__10674_
timestamp 0
transform -1 0 10230 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10675_
timestamp 0
transform -1 0 10350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__10676_
timestamp 0
transform 1 0 11050 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10677_
timestamp 0
transform 1 0 10910 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__10678_
timestamp 0
transform 1 0 11130 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10679_
timestamp 0
transform 1 0 11270 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10680_
timestamp 0
transform -1 0 9670 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10681_
timestamp 0
transform -1 0 9730 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10682_
timestamp 0
transform -1 0 10070 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__10683_
timestamp 0
transform -1 0 10110 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__10684_
timestamp 0
transform 1 0 9370 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10685_
timestamp 0
transform 1 0 9210 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10686_
timestamp 0
transform -1 0 8590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10687_
timestamp 0
transform -1 0 8710 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__10768_
timestamp 0
transform -1 0 5670 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__10769_
timestamp 0
transform -1 0 4850 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__10770_
timestamp 0
transform -1 0 4750 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__10771_
timestamp 0
transform -1 0 5530 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__10772_
timestamp 0
transform 1 0 5630 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__10773_
timestamp 0
transform -1 0 4370 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__10774_
timestamp 0
transform 1 0 5550 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__10775_
timestamp 0
transform 1 0 5570 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__10776_
timestamp 0
transform -1 0 2690 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__10777_
timestamp 0
transform 1 0 5430 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__10778_
timestamp 0
transform 1 0 5930 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__10779_
timestamp 0
transform 1 0 5770 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__10780_
timestamp 0
transform -1 0 4550 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__10781_
timestamp 0
transform -1 0 5810 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__10782_
timestamp 0
transform 1 0 5450 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__10783_
timestamp 0
transform 1 0 5110 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__10784_
timestamp 0
transform 1 0 5330 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__10785_
timestamp 0
transform 1 0 5490 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__10786_
timestamp 0
transform -1 0 6750 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__10787_
timestamp 0
transform -1 0 5610 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__10788_
timestamp 0
transform -1 0 6110 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__10789_
timestamp 0
transform 1 0 6250 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__10790_
timestamp 0
transform 1 0 6470 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__10791_
timestamp 0
transform 1 0 6630 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__10792_
timestamp 0
transform -1 0 5910 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10793_
timestamp 0
transform -1 0 5310 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__10794_
timestamp 0
transform 1 0 5450 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__10795_
timestamp 0
transform 1 0 5830 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10796_
timestamp 0
transform 1 0 6150 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__10797_
timestamp 0
transform 1 0 6010 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__10798_
timestamp 0
transform 1 0 5590 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__10799_
timestamp 0
transform 1 0 5130 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__10800_
timestamp 0
transform 1 0 6310 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__10801_
timestamp 0
transform -1 0 5630 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__10802_
timestamp 0
transform -1 0 5630 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__10803_
timestamp 0
transform 1 0 5750 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__10804_
timestamp 0
transform -1 0 5350 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__10805_
timestamp 0
transform 1 0 5750 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__10806_
timestamp 0
transform 1 0 5890 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__10807_
timestamp 0
transform 1 0 5910 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__10808_
timestamp 0
transform 1 0 5090 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__10809_
timestamp 0
transform 1 0 6190 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__10810_
timestamp 0
transform 1 0 1090 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__10811_
timestamp 0
transform 1 0 1930 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__10812_
timestamp 0
transform 1 0 1230 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__10813_
timestamp 0
transform 1 0 1550 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__10814_
timestamp 0
transform 1 0 1550 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__10815_
timestamp 0
transform -1 0 1410 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__10816_
timestamp 0
transform 1 0 1670 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__10817_
timestamp 0
transform 1 0 2770 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__10818_
timestamp 0
transform -1 0 2290 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__10819_
timestamp 0
transform 1 0 2730 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__10820_
timestamp 0
transform -1 0 2030 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__10821_
timestamp 0
transform -1 0 2150 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__10822_
timestamp 0
transform -1 0 1850 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__10823_
timestamp 0
transform 1 0 2130 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__10824_
timestamp 0
transform -1 0 2790 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__10825_
timestamp 0
transform -1 0 2970 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__10826_
timestamp 0
transform -1 0 5050 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__10827_
timestamp 0
transform -1 0 4990 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10828_
timestamp 0
transform -1 0 650 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__10829_
timestamp 0
transform -1 0 450 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__10830_
timestamp 0
transform -1 0 1270 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__10831_
timestamp 0
transform 1 0 1490 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__10832_
timestamp 0
transform 1 0 1350 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__10833_
timestamp 0
transform -1 0 50 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__10834_
timestamp 0
transform 1 0 2250 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10835_
timestamp 0
transform 1 0 2110 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10836_
timestamp 0
transform 1 0 1870 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__10837_
timestamp 0
transform 1 0 2950 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__10838_
timestamp 0
transform 1 0 3370 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__10839_
timestamp 0
transform 1 0 3050 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__10840_
timestamp 0
transform -1 0 1890 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__10841_
timestamp 0
transform 1 0 3010 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10842_
timestamp 0
transform 1 0 2630 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__10843_
timestamp 0
transform -1 0 2790 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__10844_
timestamp 0
transform -1 0 3230 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__10845_
timestamp 0
transform -1 0 4730 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__10846_
timestamp 0
transform 1 0 4830 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__10847_
timestamp 0
transform -1 0 4570 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__10848_
timestamp 0
transform -1 0 3170 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10849_
timestamp 0
transform -1 0 1450 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__10850_
timestamp 0
transform -1 0 1330 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__10851_
timestamp 0
transform -1 0 4430 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__10852_
timestamp 0
transform -1 0 4910 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__10853_
timestamp 0
transform 1 0 1810 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__10854_
timestamp 0
transform -1 0 4490 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__10855_
timestamp 0
transform 1 0 3870 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10856_
timestamp 0
transform 1 0 2650 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10857_
timestamp 0
transform 1 0 3090 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10858_
timestamp 0
transform 1 0 3390 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10859_
timestamp 0
transform -1 0 2970 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__10860_
timestamp 0
transform 1 0 3570 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__10861_
timestamp 0
transform 1 0 3490 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__10862_
timestamp 0
transform 1 0 2870 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__10863_
timestamp 0
transform 1 0 3290 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10864_
timestamp 0
transform 1 0 3430 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10865_
timestamp 0
transform 1 0 3570 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10866_
timestamp 0
transform 1 0 4410 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10867_
timestamp 0
transform 1 0 730 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__10868_
timestamp 0
transform 1 0 1730 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10869_
timestamp 0
transform 1 0 1990 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10870_
timestamp 0
transform 1 0 1830 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10871_
timestamp 0
transform -1 0 2410 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10872_
timestamp 0
transform -1 0 2050 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10873_
timestamp 0
transform -1 0 2190 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10874_
timestamp 0
transform -1 0 2270 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10875_
timestamp 0
transform -1 0 2650 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__10876_
timestamp 0
transform 1 0 2430 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__10877_
timestamp 0
transform 1 0 2190 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__10878_
timestamp 0
transform -1 0 3030 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10879_
timestamp 0
transform -1 0 1930 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__10880_
timestamp 0
transform -1 0 2070 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__10881_
timestamp 0
transform -1 0 2110 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__10882_
timestamp 0
transform -1 0 2290 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__10883_
timestamp 0
transform 1 0 3870 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10884_
timestamp 0
transform -1 0 2330 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10885_
timestamp 0
transform -1 0 2510 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10886_
timestamp 0
transform 1 0 2430 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10887_
timestamp 0
transform -1 0 3130 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10888_
timestamp 0
transform 1 0 3610 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10889_
timestamp 0
transform 1 0 3270 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10890_
timestamp 0
transform 1 0 3450 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10891_
timestamp 0
transform -1 0 4490 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10892_
timestamp 0
transform 1 0 4290 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10893_
timestamp 0
transform -1 0 4450 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10894_
timestamp 0
transform 1 0 4150 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10895_
timestamp 0
transform 1 0 4550 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10896_
timestamp 0
transform 1 0 4510 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10897_
timestamp 0
transform 1 0 4830 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10898_
timestamp 0
transform -1 0 4690 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10899_
timestamp 0
transform -1 0 4610 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__10900_
timestamp 0
transform -1 0 8350 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__10901_
timestamp 0
transform -1 0 7850 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__10902_
timestamp 0
transform -1 0 7970 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__10903_
timestamp 0
transform 1 0 5490 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__10904_
timestamp 0
transform 1 0 4690 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10905_
timestamp 0
transform -1 0 2470 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__10906_
timestamp 0
transform -1 0 2630 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10907_
timestamp 0
transform -1 0 3790 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10908_
timestamp 0
transform -1 0 3590 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10909_
timestamp 0
transform 1 0 3710 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10910_
timestamp 0
transform 1 0 3930 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10911_
timestamp 0
transform 1 0 4630 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10912_
timestamp 0
transform 1 0 4770 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10913_
timestamp 0
transform -1 0 4250 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10914_
timestamp 0
transform 1 0 4010 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10915_
timestamp 0
transform -1 0 4110 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10916_
timestamp 0
transform 1 0 4910 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10917_
timestamp 0
transform 1 0 5050 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10918_
timestamp 0
transform 1 0 5530 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10919_
timestamp 0
transform -1 0 5090 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10920_
timestamp 0
transform 1 0 4830 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10921_
timestamp 0
transform 1 0 4970 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10922_
timestamp 0
transform -1 0 5230 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10923_
timestamp 0
transform 1 0 5210 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__10924_
timestamp 0
transform -1 0 1030 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__10925_
timestamp 0
transform 1 0 5330 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10926_
timestamp 0
transform 1 0 5470 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10927_
timestamp 0
transform 1 0 5630 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10928_
timestamp 0
transform 1 0 5610 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__10929_
timestamp 0
transform 1 0 5370 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10930_
timestamp 0
transform 1 0 5350 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__10931_
timestamp 0
transform 1 0 3650 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__10932_
timestamp 0
transform -1 0 4350 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10933_
timestamp 0
transform 1 0 1250 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__10934_
timestamp 0
transform 1 0 1610 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__10935_
timestamp 0
transform 1 0 1470 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__10936_
timestamp 0
transform 1 0 1750 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__10937_
timestamp 0
transform 1 0 1470 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__10938_
timestamp 0
transform 1 0 1210 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__10939_
timestamp 0
transform -1 0 3830 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__10940_
timestamp 0
transform -1 0 2050 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__10941_
timestamp 0
transform 1 0 1830 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__10942_
timestamp 0
transform 1 0 3370 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__10943_
timestamp 0
transform 1 0 3650 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__10944_
timestamp 0
transform 1 0 3510 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__10945_
timestamp 0
transform -1 0 3790 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__10946_
timestamp 0
transform 1 0 4050 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__10947_
timestamp 0
transform 1 0 3910 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__10948_
timestamp 0
transform -1 0 4530 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__10949_
timestamp 0
transform -1 0 4650 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__10950_
timestamp 0
transform -1 0 5070 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__10951_
timestamp 0
transform -1 0 5210 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__10952_
timestamp 0
transform -1 0 5390 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__10953_
timestamp 0
transform -1 0 4770 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__10954_
timestamp 0
transform -1 0 4530 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__10955_
timestamp 0
transform -1 0 1770 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__10956_
timestamp 0
transform -1 0 1450 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__10957_
timestamp 0
transform -1 0 1570 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__10958_
timestamp 0
transform 1 0 1690 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__10959_
timestamp 0
transform 1 0 1610 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__10960_
timestamp 0
transform 1 0 3290 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__10961_
timestamp 0
transform 1 0 2390 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__10962_
timestamp 0
transform 1 0 2750 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__10963_
timestamp 0
transform 1 0 3650 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__10964_
timestamp 0
transform 1 0 3950 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__10965_
timestamp 0
transform -1 0 3390 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__10966_
timestamp 0
transform 1 0 3510 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__10967_
timestamp 0
transform 1 0 4410 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__10968_
timestamp 0
transform 1 0 3750 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__10969_
timestamp 0
transform -1 0 3630 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__10970_
timestamp 0
transform 1 0 3870 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__10971_
timestamp 0
transform -1 0 4750 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__10972_
timestamp 0
transform 1 0 4890 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__10973_
timestamp 0
transform 1 0 5050 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__10974_
timestamp 0
transform -1 0 5770 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__10975_
timestamp 0
transform -1 0 5010 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__10976_
timestamp 0
transform -1 0 4130 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__10977_
timestamp 0
transform 1 0 3790 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__10978_
timestamp 0
transform 1 0 1130 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__10979_
timestamp 0
transform 1 0 1270 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__10980_
timestamp 0
transform -1 0 1350 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__10981_
timestamp 0
transform 1 0 2530 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__10982_
timestamp 0
transform 1 0 2450 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__10983_
timestamp 0
transform 1 0 3810 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__10984_
timestamp 0
transform 1 0 2870 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__10985_
timestamp 0
transform -1 0 3130 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__10986_
timestamp 0
transform 1 0 3210 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__10987_
timestamp 0
transform 1 0 4090 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__10988_
timestamp 0
transform 1 0 4230 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__10989_
timestamp 0
transform 1 0 4850 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__10990_
timestamp 0
transform 1 0 5070 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__10991_
timestamp 0
transform 1 0 5130 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__10992_
timestamp 0
transform 1 0 5290 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__10993_
timestamp 0
transform 1 0 5430 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__10994_
timestamp 0
transform 1 0 5430 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__10995_
timestamp 0
transform -1 0 5950 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__10996_
timestamp 0
transform 1 0 1950 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__10997_
timestamp 0
transform -1 0 3190 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__10998_
timestamp 0
transform -1 0 1270 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__10999_
timestamp 0
transform -1 0 2950 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11000_
timestamp 0
transform -1 0 2230 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11001_
timestamp 0
transform 1 0 2490 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11002_
timestamp 0
transform 1 0 2650 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11003_
timestamp 0
transform -1 0 3670 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11004_
timestamp 0
transform 1 0 3190 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11005_
timestamp 0
transform 1 0 2890 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11006_
timestamp 0
transform 1 0 2750 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11007_
timestamp 0
transform 1 0 3310 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11008_
timestamp 0
transform 1 0 3430 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11009_
timestamp 0
transform 1 0 3890 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11010_
timestamp 0
transform 1 0 4250 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11011_
timestamp 0
transform -1 0 4390 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11012_
timestamp 0
transform -1 0 4590 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11013_
timestamp 0
transform -1 0 4650 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11014_
timestamp 0
transform 1 0 5190 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11015_
timestamp 0
transform 1 0 5330 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11016_
timestamp 0
transform -1 0 5790 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11017_
timestamp 0
transform 1 0 5730 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11018_
timestamp 0
transform 1 0 3050 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11019_
timestamp 0
transform 1 0 4850 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11020_
timestamp 0
transform -1 0 4930 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11021_
timestamp 0
transform 1 0 4490 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11022_
timestamp 0
transform -1 0 4770 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11023_
timestamp 0
transform -1 0 3770 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11024_
timestamp 0
transform -1 0 1290 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11025_
timestamp 0
transform -1 0 3050 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11026_
timestamp 0
transform -1 0 2110 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11027_
timestamp 0
transform -1 0 2150 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11028_
timestamp 0
transform -1 0 2050 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11029_
timestamp 0
transform -1 0 1430 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11030_
timestamp 0
transform -1 0 1570 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11031_
timestamp 0
transform 1 0 1690 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11032_
timestamp 0
transform -1 0 2350 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11033_
timestamp 0
transform 1 0 1790 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11034_
timestamp 0
transform 1 0 1390 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11035_
timestamp 0
transform 1 0 1910 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11036_
timestamp 0
transform 1 0 2190 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11037_
timestamp 0
transform 1 0 2050 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11038_
timestamp 0
transform 1 0 4010 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11039_
timestamp 0
transform 1 0 4250 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11040_
timestamp 0
transform -1 0 4150 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11041_
timestamp 0
transform -1 0 4570 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11042_
timestamp 0
transform 1 0 4710 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11043_
timestamp 0
transform 1 0 5230 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11044_
timestamp 0
transform 1 0 5390 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11045_
timestamp 0
transform 1 0 5190 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11046_
timestamp 0
transform -1 0 5350 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11047_
timestamp 0
transform -1 0 5670 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11048_
timestamp 0
transform -1 0 4150 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11049_
timestamp 0
transform 1 0 4430 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11050_
timestamp 0
transform -1 0 4310 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11051_
timestamp 0
transform -1 0 2790 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11052_
timestamp 0
transform 1 0 2190 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11053_
timestamp 0
transform -1 0 1590 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11054_
timestamp 0
transform 1 0 2330 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11055_
timestamp 0
transform -1 0 1970 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11056_
timestamp 0
transform 1 0 2350 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11057_
timestamp 0
transform 1 0 2610 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11058_
timestamp 0
transform -1 0 2630 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11059_
timestamp 0
transform 1 0 2470 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11060_
timestamp 0
transform -1 0 2470 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11061_
timestamp 0
transform 1 0 2890 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11062_
timestamp 0
transform -1 0 3890 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11063_
timestamp 0
transform 1 0 4910 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11064_
timestamp 0
transform 1 0 5030 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11065_
timestamp 0
transform 1 0 5170 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11066_
timestamp 0
transform -1 0 5510 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11067_
timestamp 0
transform -1 0 3330 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11068_
timestamp 0
transform 1 0 3590 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11069_
timestamp 0
transform -1 0 3470 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11070_
timestamp 0
transform 1 0 3590 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11071_
timestamp 0
transform -1 0 3750 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11072_
timestamp 0
transform -1 0 4030 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11073_
timestamp 0
transform 1 0 3950 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11074_
timestamp 0
transform 1 0 3250 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11075_
timestamp 0
transform 1 0 1730 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11076_
timestamp 0
transform 1 0 2950 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11077_
timestamp 0
transform -1 0 2310 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11078_
timestamp 0
transform 1 0 3110 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11079_
timestamp 0
transform 1 0 2610 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11080_
timestamp 0
transform 1 0 2830 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11081_
timestamp 0
transform 1 0 3510 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11082_
timestamp 0
transform 1 0 3050 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11083_
timestamp 0
transform 1 0 2970 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11084_
timestamp 0
transform 1 0 3210 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11085_
timestamp 0
transform 1 0 4030 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11086_
timestamp 0
transform 1 0 4450 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11087_
timestamp 0
transform 1 0 4610 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11088_
timestamp 0
transform 1 0 4750 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11089_
timestamp 0
transform -1 0 5470 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11090_
timestamp 0
transform -1 0 3790 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11091_
timestamp 0
transform 1 0 2130 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11092_
timestamp 0
transform 1 0 2730 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11093_
timestamp 0
transform 1 0 2650 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11094_
timestamp 0
transform 1 0 2790 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11095_
timestamp 0
transform -1 0 2990 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11096_
timestamp 0
transform -1 0 3530 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11097_
timestamp 0
transform 1 0 3650 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11098_
timestamp 0
transform -1 0 3950 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11099_
timestamp 0
transform 1 0 3550 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11100_
timestamp 0
transform 1 0 3090 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11101_
timestamp 0
transform -1 0 3430 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11102_
timestamp 0
transform 1 0 3790 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11103_
timestamp 0
transform -1 0 4370 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11104_
timestamp 0
transform 1 0 3370 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11105_
timestamp 0
transform 1 0 4090 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11106_
timestamp 0
transform 1 0 4310 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11107_
timestamp 0
transform 1 0 4370 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11108_
timestamp 0
transform 1 0 4490 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11109_
timestamp 0
transform 1 0 4170 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11110_
timestamp 0
transform 1 0 4210 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11111_
timestamp 0
transform 1 0 4910 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11112_
timestamp 0
transform 1 0 5090 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11113_
timestamp 0
transform -1 0 5730 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__11114_
timestamp 0
transform -1 0 6090 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11115_
timestamp 0
transform 1 0 4650 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11116_
timestamp 0
transform -1 0 2610 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11117_
timestamp 0
transform -1 0 2450 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11118_
timestamp 0
transform -1 0 1990 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11119_
timestamp 0
transform -1 0 2490 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11120_
timestamp 0
transform -1 0 3030 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11121_
timestamp 0
transform 1 0 3130 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11122_
timestamp 0
transform 1 0 3270 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11123_
timestamp 0
transform 1 0 3250 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11124_
timestamp 0
transform 1 0 4450 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11125_
timestamp 0
transform 1 0 4550 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11126_
timestamp 0
transform -1 0 4790 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11127_
timestamp 0
transform 1 0 4790 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11128_
timestamp 0
transform 1 0 4950 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11129_
timestamp 0
transform -1 0 5950 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11130_
timestamp 0
transform 1 0 1990 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11131_
timestamp 0
transform -1 0 3450 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11132_
timestamp 0
transform 1 0 3510 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11133_
timestamp 0
transform -1 0 3390 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11134_
timestamp 0
transform 1 0 2330 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11135_
timestamp 0
transform -1 0 4090 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11136_
timestamp 0
transform 1 0 3710 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11137_
timestamp 0
transform -1 0 4270 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__11138_
timestamp 0
transform -1 0 2210 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11139_
timestamp 0
transform 1 0 1130 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11140_
timestamp 0
transform 1 0 990 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11141_
timestamp 0
transform -1 0 4090 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11142_
timestamp 0
transform -1 0 4230 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11143_
timestamp 0
transform 1 0 730 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11144_
timestamp 0
transform 1 0 150 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11145_
timestamp 0
transform -1 0 1470 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11146_
timestamp 0
transform -1 0 1370 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11147_
timestamp 0
transform 1 0 890 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11148_
timestamp 0
transform -1 0 1150 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11149_
timestamp 0
transform 1 0 1010 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11150_
timestamp 0
transform 1 0 1750 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11151_
timestamp 0
transform -1 0 1650 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11152_
timestamp 0
transform 1 0 1610 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11153_
timestamp 0
transform -1 0 2550 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11154_
timestamp 0
transform -1 0 1930 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__11155_
timestamp 0
transform 1 0 3370 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11156_
timestamp 0
transform 1 0 3230 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11157_
timestamp 0
transform 1 0 3530 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11158_
timestamp 0
transform -1 0 3670 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11159_
timestamp 0
transform 1 0 1690 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11160_
timestamp 0
transform 1 0 450 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11161_
timestamp 0
transform 1 0 870 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11162_
timestamp 0
transform -1 0 750 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11163_
timestamp 0
transform -1 0 50 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11164_
timestamp 0
transform 1 0 1830 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11165_
timestamp 0
transform 1 0 1670 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11166_
timestamp 0
transform 1 0 310 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11167_
timestamp 0
transform 1 0 150 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__11168_
timestamp 0
transform 1 0 310 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11169_
timestamp 0
transform 1 0 1230 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11170_
timestamp 0
transform 1 0 550 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11171_
timestamp 0
transform -1 0 750 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11172_
timestamp 0
transform -1 0 1610 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11173_
timestamp 0
transform 1 0 1650 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11174_
timestamp 0
transform 1 0 1850 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11175_
timestamp 0
transform -1 0 1510 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11176_
timestamp 0
transform 1 0 1950 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11177_
timestamp 0
transform 1 0 1950 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11178_
timestamp 0
transform -1 0 1830 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11179_
timestamp 0
transform 1 0 2090 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11180_
timestamp 0
transform 1 0 2390 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11181_
timestamp 0
transform -1 0 2150 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11182_
timestamp 0
transform -1 0 1710 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11183_
timestamp 0
transform 1 0 1170 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11184_
timestamp 0
transform 1 0 1530 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11185_
timestamp 0
transform 1 0 1390 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11186_
timestamp 0
transform 1 0 590 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11187_
timestamp 0
transform -1 0 470 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11188_
timestamp 0
transform 1 0 1850 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11189_
timestamp 0
transform 1 0 1290 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11190_
timestamp 0
transform -1 0 1190 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11191_
timestamp 0
transform 1 0 890 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11192_
timestamp 0
transform 1 0 790 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11193_
timestamp 0
transform 1 0 890 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11194_
timestamp 0
transform -1 0 1310 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11195_
timestamp 0
transform -1 0 1050 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11196_
timestamp 0
transform -1 0 930 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11197_
timestamp 0
transform 1 0 1050 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11198_
timestamp 0
transform 1 0 1070 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11199_
timestamp 0
transform 1 0 1150 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11200_
timestamp 0
transform 1 0 1410 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11201_
timestamp 0
transform -1 0 1290 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11202_
timestamp 0
transform 1 0 1550 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11203_
timestamp 0
transform 1 0 1970 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11204_
timestamp 0
transform -1 0 930 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11205_
timestamp 0
transform -1 0 330 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11206_
timestamp 0
transform 1 0 1990 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11207_
timestamp 0
transform 1 0 1890 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11208_
timestamp 0
transform -1 0 610 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11209_
timestamp 0
transform 1 0 170 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11210_
timestamp 0
transform -1 0 1570 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11211_
timestamp 0
transform -1 0 1330 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11212_
timestamp 0
transform 1 0 1430 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11213_
timestamp 0
transform -1 0 50 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11214_
timestamp 0
transform -1 0 770 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11215_
timestamp 0
transform 1 0 310 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11216_
timestamp 0
transform 1 0 330 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11217_
timestamp 0
transform 1 0 570 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11218_
timestamp 0
transform -1 0 190 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11219_
timestamp 0
transform -1 0 450 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11220_
timestamp 0
transform -1 0 50 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11221_
timestamp 0
transform 1 0 170 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11222_
timestamp 0
transform -1 0 50 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11223_
timestamp 0
transform 1 0 410 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11224_
timestamp 0
transform -1 0 2350 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11225_
timestamp 0
transform -1 0 290 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11226_
timestamp 0
transform -1 0 2570 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11227_
timestamp 0
transform -1 0 2690 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11228_
timestamp 0
transform -1 0 310 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11229_
timestamp 0
transform -1 0 310 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11230_
timestamp 0
transform 1 0 30 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11231_
timestamp 0
transform -1 0 170 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__11232_
timestamp 0
transform 1 0 330 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11233_
timestamp 0
transform -1 0 490 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11234_
timestamp 0
transform 1 0 150 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11235_
timestamp 0
transform -1 0 190 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__11236_
timestamp 0
transform -1 0 50 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11237_
timestamp 0
transform -1 0 50 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11238_
timestamp 0
transform -1 0 50 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__11239_
timestamp 0
transform 1 0 310 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__11240_
timestamp 0
transform 1 0 190 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11241_
timestamp 0
transform -1 0 50 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11242_
timestamp 0
transform -1 0 50 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11243_
timestamp 0
transform 1 0 330 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11244_
timestamp 0
transform -1 0 210 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11245_
timestamp 0
transform -1 0 490 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11246_
timestamp 0
transform -1 0 1150 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11247_
timestamp 0
transform -1 0 210 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11248_
timestamp 0
transform -1 0 50 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11249_
timestamp 0
transform -1 0 50 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__11250_
timestamp 0
transform 1 0 1090 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11251_
timestamp 0
transform -1 0 790 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11252_
timestamp 0
transform -1 0 50 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11253_
timestamp 0
transform -1 0 170 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11254_
timestamp 0
transform 1 0 470 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__11255_
timestamp 0
transform -1 0 310 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__11256_
timestamp 0
transform -1 0 210 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11257_
timestamp 0
transform 1 0 610 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11258_
timestamp 0
transform -1 0 550 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11259_
timestamp 0
transform 1 0 450 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11260_
timestamp 0
transform -1 0 350 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11261_
timestamp 0
transform -1 0 210 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11262_
timestamp 0
transform 1 0 490 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11263_
timestamp 0
transform -1 0 170 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11264_
timestamp 0
transform -1 0 50 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11265_
timestamp 0
transform 1 0 150 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11266_
timestamp 0
transform 1 0 310 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11267_
timestamp 0
transform -1 0 50 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11268_
timestamp 0
transform -1 0 1510 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11269_
timestamp 0
transform 1 0 150 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__11270_
timestamp 0
transform -1 0 950 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__11271_
timestamp 0
transform 1 0 550 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11272_
timestamp 0
transform 1 0 470 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__11273_
timestamp 0
transform 1 0 430 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__11274_
timestamp 0
transform 1 0 690 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11275_
timestamp 0
transform -1 0 590 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11276_
timestamp 0
transform -1 0 710 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11277_
timestamp 0
transform -1 0 450 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11278_
timestamp 0
transform -1 0 590 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11279_
timestamp 0
transform 1 0 570 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11280_
timestamp 0
transform -1 0 710 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11281_
timestamp 0
transform 1 0 190 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11282_
timestamp 0
transform -1 0 150 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11283_
timestamp 0
transform -1 0 310 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11284_
timestamp 0
transform 1 0 430 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11285_
timestamp 0
transform -1 0 590 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11286_
timestamp 0
transform 1 0 710 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11287_
timestamp 0
transform 1 0 30 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11288_
timestamp 0
transform 1 0 290 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11289_
timestamp 0
transform 1 0 270 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11290_
timestamp 0
transform 1 0 430 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11291_
timestamp 0
transform 1 0 850 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11292_
timestamp 0
transform 1 0 990 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11293_
timestamp 0
transform -1 0 1230 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11294_
timestamp 0
transform -1 0 1350 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11295_
timestamp 0
transform -1 0 1230 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11296_
timestamp 0
transform -1 0 610 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11297_
timestamp 0
transform 1 0 830 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11298_
timestamp 0
transform -1 0 1190 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11299_
timestamp 0
transform -1 0 990 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11300_
timestamp 0
transform 1 0 290 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11301_
timestamp 0
transform 1 0 890 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11302_
timestamp 0
transform 1 0 730 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__11303_
timestamp 0
transform 1 0 570 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__11304_
timestamp 0
transform -1 0 710 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__11305_
timestamp 0
transform -1 0 770 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11306_
timestamp 0
transform 1 0 810 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__11307_
timestamp 0
transform -1 0 590 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__11308_
timestamp 0
transform -1 0 990 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__11309_
timestamp 0
transform 1 0 730 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11310_
timestamp 0
transform 1 0 150 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11311_
timestamp 0
transform -1 0 50 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11312_
timestamp 0
transform 1 0 450 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11313_
timestamp 0
transform 1 0 550 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11314_
timestamp 0
transform -1 0 830 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11315_
timestamp 0
transform 1 0 690 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11316_
timestamp 0
transform 1 0 810 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11317_
timestamp 0
transform 1 0 930 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11318_
timestamp 0
transform -1 0 870 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11319_
timestamp 0
transform 1 0 830 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__11320_
timestamp 0
transform -1 0 50 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__11321_
timestamp 0
transform -1 0 50 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11322_
timestamp 0
transform -1 0 1110 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11323_
timestamp 0
transform 1 0 1230 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__11324_
timestamp 0
transform 1 0 950 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11325_
timestamp 0
transform -1 0 990 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__11326_
timestamp 0
transform 1 0 1050 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11327_
timestamp 0
transform -1 0 1310 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__11328_
timestamp 0
transform -1 0 1130 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__11329_
timestamp 0
transform 1 0 1130 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__11330_
timestamp 0
transform -1 0 730 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11331_
timestamp 0
transform -1 0 730 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11332_
timestamp 0
transform 1 0 1270 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11333_
timestamp 0
transform -1 0 330 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11334_
timestamp 0
transform -1 0 550 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11335_
timestamp 0
transform 1 0 870 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11336_
timestamp 0
transform -1 0 470 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11337_
timestamp 0
transform -1 0 590 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11338_
timestamp 0
transform 1 0 670 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11339_
timestamp 0
transform 1 0 1370 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__11340_
timestamp 0
transform 1 0 1450 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__11341_
timestamp 0
transform 1 0 1330 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11342_
timestamp 0
transform -1 0 1210 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11343_
timestamp 0
transform -1 0 1130 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11344_
timestamp 0
transform -1 0 990 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11345_
timestamp 0
transform -1 0 1010 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11346_
timestamp 0
transform 1 0 1130 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11347_
timestamp 0
transform -1 0 870 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11348_
timestamp 0
transform 1 0 990 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11349_
timestamp 0
transform -1 0 730 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11350_
timestamp 0
transform -1 0 1850 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11351_
timestamp 0
transform -1 0 1090 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11352_
timestamp 0
transform 1 0 1190 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11353_
timestamp 0
transform -1 0 870 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11354_
timestamp 0
transform 1 0 1110 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11355_
timestamp 0
transform 1 0 1330 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11356_
timestamp 0
transform 1 0 810 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11357_
timestamp 0
transform 1 0 1070 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__11358_
timestamp 0
transform 1 0 1210 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11359_
timestamp 0
transform 1 0 1370 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11360_
timestamp 0
transform -1 0 1530 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11361_
timestamp 0
transform 1 0 1490 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__11362_
timestamp 0
transform -1 0 1610 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__11363_
timestamp 0
transform 1 0 1650 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__11364_
timestamp 0
transform -1 0 1650 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__11365_
timestamp 0
transform 1 0 1750 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__11366_
timestamp 0
transform -1 0 1510 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11367_
timestamp 0
transform 1 0 1610 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11368_
timestamp 0
transform -1 0 1490 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11369_
timestamp 0
transform 1 0 1750 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11370_
timestamp 0
transform -1 0 1670 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11371_
timestamp 0
transform -1 0 1590 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11372_
timestamp 0
transform -1 0 1450 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11373_
timestamp 0
transform 1 0 1550 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11374_
timestamp 0
transform 1 0 1370 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11375_
timestamp 0
transform -1 0 2370 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11376_
timestamp 0
transform -1 0 2750 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11377_
timestamp 0
transform -1 0 2510 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__11378_
timestamp 0
transform 1 0 1850 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11379_
timestamp 0
transform -1 0 1710 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11380_
timestamp 0
transform -1 0 1710 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11381_
timestamp 0
transform -1 0 2410 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11382_
timestamp 0
transform 1 0 4230 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11383_
timestamp 0
transform 1 0 4390 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11384_
timestamp 0
transform -1 0 3970 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11385_
timestamp 0
transform 1 0 4490 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11386_
timestamp 0
transform 1 0 4750 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11387_
timestamp 0
transform 1 0 5970 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11388_
timestamp 0
transform 1 0 5410 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11389_
timestamp 0
transform -1 0 6110 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11390_
timestamp 0
transform 1 0 4710 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11391_
timestamp 0
transform -1 0 3590 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11392_
timestamp 0
transform -1 0 3690 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11393_
timestamp 0
transform 1 0 4610 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11394_
timestamp 0
transform 1 0 3790 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11395_
timestamp 0
transform 1 0 4730 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11396_
timestamp 0
transform -1 0 4890 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11397_
timestamp 0
transform 1 0 5170 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11398_
timestamp 0
transform 1 0 5030 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11399_
timestamp 0
transform 1 0 5310 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11400_
timestamp 0
transform 1 0 5450 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11401_
timestamp 0
transform 1 0 4950 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11402_
timestamp 0
transform 1 0 5810 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11403_
timestamp 0
transform 1 0 5930 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11404_
timestamp 0
transform -1 0 4630 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11405_
timestamp 0
transform 1 0 4810 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11406_
timestamp 0
transform -1 0 2790 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11407_
timestamp 0
transform 1 0 3270 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11408_
timestamp 0
transform 1 0 3090 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11409_
timestamp 0
transform -1 0 4110 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11410_
timestamp 0
transform 1 0 4210 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11411_
timestamp 0
transform -1 0 4390 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11412_
timestamp 0
transform 1 0 4390 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11413_
timestamp 0
transform 1 0 5210 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11414_
timestamp 0
transform -1 0 5110 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11415_
timestamp 0
transform -1 0 5370 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11416_
timestamp 0
transform -1 0 5510 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11417_
timestamp 0
transform -1 0 6690 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11418_
timestamp 0
transform 1 0 5310 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11419_
timestamp 0
transform -1 0 6290 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11420_
timestamp 0
transform 1 0 5190 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11421_
timestamp 0
transform -1 0 3610 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11422_
timestamp 0
transform -1 0 3730 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11423_
timestamp 0
transform 1 0 3410 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11424_
timestamp 0
transform 1 0 3610 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11425_
timestamp 0
transform 1 0 6650 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11426_
timestamp 0
transform -1 0 6550 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11427_
timestamp 0
transform 1 0 7170 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11428_
timestamp 0
transform 1 0 7050 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11429_
timestamp 0
transform -1 0 6390 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11430_
timestamp 0
transform 1 0 6510 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11431_
timestamp 0
transform 1 0 6790 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11432_
timestamp 0
transform 1 0 6110 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11433_
timestamp 0
transform 1 0 6510 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__11434_
timestamp 0
transform 1 0 3810 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11435_
timestamp 0
transform 1 0 3970 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11436_
timestamp 0
transform -1 0 4490 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11437_
timestamp 0
transform 1 0 6690 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11438_
timestamp 0
transform -1 0 6490 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11439_
timestamp 0
transform 1 0 6850 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11440_
timestamp 0
transform 1 0 6910 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11441_
timestamp 0
transform -1 0 6130 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11442_
timestamp 0
transform -1 0 5990 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11443_
timestamp 0
transform -1 0 5850 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11444_
timestamp 0
transform 1 0 6990 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11445_
timestamp 0
transform 1 0 6130 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__11446_
timestamp 0
transform -1 0 3930 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11447_
timestamp 0
transform -1 0 3930 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11448_
timestamp 0
transform 1 0 4010 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11449_
timestamp 0
transform 1 0 4150 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11450_
timestamp 0
transform 1 0 6370 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__11451_
timestamp 0
transform -1 0 6250 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__11452_
timestamp 0
transform 1 0 6610 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__11453_
timestamp 0
transform 1 0 6890 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__11454_
timestamp 0
transform 1 0 7310 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11455_
timestamp 0
transform 1 0 7270 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__11456_
timestamp 0
transform -1 0 7410 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__11457_
timestamp 0
transform 1 0 7150 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11458_
timestamp 0
transform -1 0 6410 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11459_
timestamp 0
transform -1 0 6370 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11460_
timestamp 0
transform -1 0 6470 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11461_
timestamp 0
transform -1 0 6750 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__11462_
timestamp 0
transform -1 0 6610 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11463_
timestamp 0
transform 1 0 6570 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11464_
timestamp 0
transform 1 0 3870 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11465_
timestamp 0
transform -1 0 4310 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11466_
timestamp 0
transform -1 0 4590 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11467_
timestamp 0
transform 1 0 4430 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11468_
timestamp 0
transform 1 0 4690 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11469_
timestamp 0
transform -1 0 5210 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11470_
timestamp 0
transform 1 0 5310 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11471_
timestamp 0
transform -1 0 5490 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11472_
timestamp 0
transform 1 0 6070 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11473_
timestamp 0
transform 1 0 7050 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11474_
timestamp 0
transform 1 0 6930 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11475_
timestamp 0
transform 1 0 6770 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11476_
timestamp 0
transform -1 0 6810 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11477_
timestamp 0
transform 1 0 5690 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11478_
timestamp 0
transform 1 0 6070 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11479_
timestamp 0
transform 1 0 5310 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11480_
timestamp 0
transform -1 0 3410 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11481_
timestamp 0
transform 1 0 3530 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11482_
timestamp 0
transform 1 0 3670 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11483_
timestamp 0
transform 1 0 5650 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11484_
timestamp 0
transform 1 0 5770 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11485_
timestamp 0
transform -1 0 5550 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11486_
timestamp 0
transform 1 0 5890 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11487_
timestamp 0
transform 1 0 6130 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11488_
timestamp 0
transform -1 0 6010 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11489_
timestamp 0
transform 1 0 5810 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11490_
timestamp 0
transform -1 0 5470 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11491_
timestamp 0
transform -1 0 2550 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11492_
timestamp 0
transform 1 0 2650 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11493_
timestamp 0
transform 1 0 3070 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11494_
timestamp 0
transform -1 0 3510 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11495_
timestamp 0
transform 1 0 3210 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11496_
timestamp 0
transform 1 0 3350 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11497_
timestamp 0
transform -1 0 6030 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11498_
timestamp 0
transform -1 0 5970 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11499_
timestamp 0
transform -1 0 6070 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11500_
timestamp 0
transform -1 0 6230 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11501_
timestamp 0
transform -1 0 5910 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11502_
timestamp 0
transform 1 0 5070 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11503_
timestamp 0
transform -1 0 4950 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11504_
timestamp 0
transform -1 0 5210 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11505_
timestamp 0
transform 1 0 5310 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11506_
timestamp 0
transform -1 0 4330 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11507_
timestamp 0
transform -1 0 3770 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11508_
timestamp 0
transform -1 0 3830 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11509_
timestamp 0
transform -1 0 3910 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11510_
timestamp 0
transform 1 0 4470 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11511_
timestamp 0
transform 1 0 4610 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11512_
timestamp 0
transform -1 0 4790 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11513_
timestamp 0
transform 1 0 5170 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11514_
timestamp 0
transform 1 0 4010 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11515_
timestamp 0
transform 1 0 4150 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11516_
timestamp 0
transform 1 0 4490 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11517_
timestamp 0
transform 1 0 4590 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11518_
timestamp 0
transform 1 0 3290 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11519_
timestamp 0
transform -1 0 3430 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11520_
timestamp 0
transform -1 0 3550 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11521_
timestamp 0
transform 1 0 3670 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11522_
timestamp 0
transform -1 0 4510 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11523_
timestamp 0
transform 1 0 4650 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11524_
timestamp 0
transform 1 0 4790 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11525_
timestamp 0
transform 1 0 5270 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11526_
timestamp 0
transform -1 0 4630 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11527_
timestamp 0
transform 1 0 5110 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11528_
timestamp 0
transform -1 0 4070 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11529_
timestamp 0
transform 1 0 2690 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11530_
timestamp 0
transform -1 0 3790 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11531_
timestamp 0
transform 1 0 2110 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11532_
timestamp 0
transform 1 0 2050 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11533_
timestamp 0
transform 1 0 2810 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11534_
timestamp 0
transform 1 0 2710 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11535_
timestamp 0
transform -1 0 2090 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11536_
timestamp 0
transform -1 0 3450 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11537_
timestamp 0
transform -1 0 2490 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11538_
timestamp 0
transform -1 0 2650 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11539_
timestamp 0
transform -1 0 2770 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11540_
timestamp 0
transform -1 0 2490 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11541_
timestamp 0
transform -1 0 2630 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11542_
timestamp 0
transform -1 0 3310 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11543_
timestamp 0
transform -1 0 2190 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11544_
timestamp 0
transform -1 0 2310 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11545_
timestamp 0
transform -1 0 2330 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11546_
timestamp 0
transform -1 0 2450 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11547_
timestamp 0
transform 1 0 1990 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11548_
timestamp 0
transform 1 0 2190 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11549_
timestamp 0
transform 1 0 2030 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11550_
timestamp 0
transform 1 0 2890 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__11551_
timestamp 0
transform 1 0 2730 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__11552_
timestamp 0
transform -1 0 3430 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11553_
timestamp 0
transform 1 0 3250 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11554_
timestamp 0
transform -1 0 3230 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11555_
timestamp 0
transform 1 0 3070 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11556_
timestamp 0
transform 1 0 2630 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11557_
timestamp 0
transform -1 0 2510 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11558_
timestamp 0
transform 1 0 2950 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__11559_
timestamp 0
transform 1 0 2810 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__11560_
timestamp 0
transform -1 0 4130 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11561_
timestamp 0
transform 1 0 3950 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11562_
timestamp 0
transform -1 0 3190 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11563_
timestamp 0
transform 1 0 3110 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__11564_
timestamp 0
transform -1 0 4270 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11565_
timestamp 0
transform 1 0 3710 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11566_
timestamp 0
transform -1 0 4130 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11567_
timestamp 0
transform 1 0 3550 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__11568_
timestamp 0
transform -1 0 3290 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11569_
timestamp 0
transform -1 0 3450 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__11570_
timestamp 0
transform 1 0 4190 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11571_
timestamp 0
transform 1 0 4330 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11572_
timestamp 0
transform 1 0 3310 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11573_
timestamp 0
transform -1 0 3450 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__11574_
timestamp 0
transform 1 0 5010 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11575_
timestamp 0
transform 1 0 4850 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11576_
timestamp 0
transform 1 0 4390 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11577_
timestamp 0
transform 1 0 4230 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__11578_
timestamp 0
transform -1 0 4290 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11579_
timestamp 0
transform -1 0 4150 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11580_
timestamp 0
transform 1 0 3350 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11581_
timestamp 0
transform -1 0 3530 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__11582_
timestamp 0
transform 1 0 5110 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11583_
timestamp 0
transform 1 0 4970 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11584_
timestamp 0
transform -1 0 3650 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11585_
timestamp 0
transform 1 0 3770 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__11586_
timestamp 0
transform -1 0 3610 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11587_
timestamp 0
transform 1 0 3310 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11588_
timestamp 0
transform -1 0 3290 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11589_
timestamp 0
transform -1 0 3130 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11590_
timestamp 0
transform 1 0 6250 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11591_
timestamp 0
transform 1 0 2930 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__11592_
timestamp 0
transform -1 0 3810 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11593_
timestamp 0
transform 1 0 4190 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11594_
timestamp 0
transform 1 0 3850 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11595_
timestamp 0
transform -1 0 4030 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11596_
timestamp 0
transform -1 0 4830 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11597_
timestamp 0
transform 1 0 4670 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11598_
timestamp 0
transform 1 0 4550 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11599_
timestamp 0
transform 1 0 4390 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__11600_
timestamp 0
transform -1 0 6830 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__11601_
timestamp 0
transform 1 0 6650 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__11602_
timestamp 0
transform -1 0 5890 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__11603_
timestamp 0
transform -1 0 6010 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__11604_
timestamp 0
transform 1 0 3950 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11605_
timestamp 0
transform -1 0 4130 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11606_
timestamp 0
transform 1 0 4790 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11607_
timestamp 0
transform 1 0 4650 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__11608_
timestamp 0
transform -1 0 3730 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11609_
timestamp 0
transform -1 0 3870 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11610_
timestamp 0
transform -1 0 4130 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11611_
timestamp 0
transform -1 0 4250 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11692_
timestamp 0
transform 1 0 9890 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__11693_
timestamp 0
transform 1 0 11330 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11694_
timestamp 0
transform -1 0 12630 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__11695_
timestamp 0
transform 1 0 13270 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__11696_
timestamp 0
transform 1 0 11510 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__11697_
timestamp 0
transform -1 0 11430 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11698_
timestamp 0
transform -1 0 11770 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11699_
timestamp 0
transform -1 0 11090 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__11700_
timestamp 0
transform -1 0 11850 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__11701_
timestamp 0
transform -1 0 11590 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11702_
timestamp 0
transform -1 0 10810 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11703_
timestamp 0
transform -1 0 10930 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__11704_
timestamp 0
transform -1 0 11230 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11705_
timestamp 0
transform -1 0 11890 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__11706_
timestamp 0
transform 1 0 12050 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__11707_
timestamp 0
transform 1 0 11490 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11708_
timestamp 0
transform -1 0 11910 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11709_
timestamp 0
transform -1 0 11630 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11710_
timestamp 0
transform 1 0 9610 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11711_
timestamp 0
transform 1 0 10790 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11712_
timestamp 0
transform -1 0 10930 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11713_
timestamp 0
transform 1 0 11070 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11714_
timestamp 0
transform 1 0 11410 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__11715_
timestamp 0
transform 1 0 11210 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11716_
timestamp 0
transform -1 0 13790 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11717_
timestamp 0
transform -1 0 13490 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11718_
timestamp 0
transform -1 0 13650 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11719_
timestamp 0
transform -1 0 13550 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11720_
timestamp 0
transform -1 0 13130 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11721_
timestamp 0
transform 1 0 12970 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11722_
timestamp 0
transform -1 0 12930 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11723_
timestamp 0
transform -1 0 12430 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11724_
timestamp 0
transform 1 0 12850 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11725_
timestamp 0
transform -1 0 13370 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11726_
timestamp 0
transform 1 0 13170 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11727_
timestamp 0
transform 1 0 13330 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11728_
timestamp 0
transform 1 0 12450 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11729_
timestamp 0
transform 1 0 12830 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11730_
timestamp 0
transform 1 0 12690 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11731_
timestamp 0
transform -1 0 12770 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11732_
timestamp 0
transform 1 0 12570 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11733_
timestamp 0
transform 1 0 12730 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11734_
timestamp 0
transform -1 0 13210 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11735_
timestamp 0
transform -1 0 13030 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11736_
timestamp 0
transform -1 0 13050 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11737_
timestamp 0
transform -1 0 13410 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11738_
timestamp 0
transform -1 0 12350 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11739_
timestamp 0
transform -1 0 12490 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11740_
timestamp 0
transform -1 0 12630 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11741_
timestamp 0
transform 1 0 12970 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__11742_
timestamp 0
transform -1 0 12930 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11743_
timestamp 0
transform -1 0 14570 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11744_
timestamp 0
transform 1 0 12890 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11745_
timestamp 0
transform -1 0 12970 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__11746_
timestamp 0
transform 1 0 12750 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11747_
timestamp 0
transform -1 0 12770 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11748_
timestamp 0
transform -1 0 12590 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11749_
timestamp 0
transform -1 0 14250 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11750_
timestamp 0
transform 1 0 12470 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__11751_
timestamp 0
transform 1 0 12750 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__11752_
timestamp 0
transform 1 0 16210 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11753_
timestamp 0
transform -1 0 16150 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__11754_
timestamp 0
transform -1 0 14770 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11755_
timestamp 0
transform 1 0 14990 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11756_
timestamp 0
transform 1 0 14850 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11757_
timestamp 0
transform -1 0 16310 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__11758_
timestamp 0
transform -1 0 15710 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__11759_
timestamp 0
transform 1 0 15810 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__11760_
timestamp 0
transform 1 0 14830 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__11761_
timestamp 0
transform 1 0 13210 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__11762_
timestamp 0
transform 1 0 13310 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__11763_
timestamp 0
transform 1 0 13070 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__11764_
timestamp 0
transform 1 0 13130 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__11765_
timestamp 0
transform 1 0 13370 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__11766_
timestamp 0
transform 1 0 13230 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__11767_
timestamp 0
transform -1 0 12910 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__11768_
timestamp 0
transform 1 0 12730 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__11769_
timestamp 0
transform 1 0 13130 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__11770_
timestamp 0
transform -1 0 12650 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11771_
timestamp 0
transform 1 0 12890 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11772_
timestamp 0
transform 1 0 14870 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__11773_
timestamp 0
transform -1 0 12450 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11774_
timestamp 0
transform -1 0 13290 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__11775_
timestamp 0
transform -1 0 13010 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__11776_
timestamp 0
transform 1 0 12590 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__11777_
timestamp 0
transform -1 0 12170 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__11778_
timestamp 0
transform -1 0 12430 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__11779_
timestamp 0
transform -1 0 13950 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__11780_
timestamp 0
transform -1 0 15230 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__11781_
timestamp 0
transform 1 0 15290 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__11782_
timestamp 0
transform -1 0 15070 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__11783_
timestamp 0
transform 1 0 12450 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__11784_
timestamp 0
transform -1 0 13170 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__11785_
timestamp 0
transform 1 0 13290 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__11786_
timestamp 0
transform -1 0 12870 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__11787_
timestamp 0
transform -1 0 13030 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__11788_
timestamp 0
transform 1 0 12830 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__11789_
timestamp 0
transform -1 0 13150 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__11790_
timestamp 0
transform -1 0 12310 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11791_
timestamp 0
transform -1 0 12010 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11792_
timestamp 0
transform 1 0 15610 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__11793_
timestamp 0
transform -1 0 15430 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__11794_
timestamp 0
transform -1 0 15570 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__11795_
timestamp 0
transform -1 0 15630 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__11796_
timestamp 0
transform -1 0 15150 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11797_
timestamp 0
transform 1 0 15270 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__11798_
timestamp 0
transform 1 0 15630 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__11799_
timestamp 0
transform -1 0 14810 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__11800_
timestamp 0
transform 1 0 15350 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__11801_
timestamp 0
transform -1 0 15510 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__11802_
timestamp 0
transform 1 0 13450 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__11803_
timestamp 0
transform -1 0 14910 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__11804_
timestamp 0
transform 1 0 15030 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__11805_
timestamp 0
transform -1 0 15190 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__11806_
timestamp 0
transform -1 0 15150 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__11807_
timestamp 0
transform -1 0 13410 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__11808_
timestamp 0
transform 1 0 15370 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__11809_
timestamp 0
transform -1 0 15490 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__11810_
timestamp 0
transform -1 0 15550 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__11811_
timestamp 0
transform 1 0 14630 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__11812_
timestamp 0
transform 1 0 13430 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__11813_
timestamp 0
transform -1 0 14550 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__11814_
timestamp 0
transform -1 0 14630 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__11815_
timestamp 0
transform 1 0 13270 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11816_
timestamp 0
transform -1 0 13010 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11817_
timestamp 0
transform -1 0 12370 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__11818_
timestamp 0
transform -1 0 13150 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11819_
timestamp 0
transform 1 0 12470 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__11820_
timestamp 0
transform -1 0 12650 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__11821_
timestamp 0
transform 1 0 12830 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__11822_
timestamp 0
transform -1 0 12690 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__11823_
timestamp 0
transform -1 0 12550 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__11824_
timestamp 0
transform 1 0 9350 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11825_
timestamp 0
transform -1 0 8730 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11826_
timestamp 0
transform -1 0 8850 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__11827_
timestamp 0
transform 1 0 12490 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11828_
timestamp 0
transform 1 0 12750 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11829_
timestamp 0
transform 1 0 15310 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__11830_
timestamp 0
transform 1 0 15150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__11831_
timestamp 0
transform 1 0 14690 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__11832_
timestamp 0
transform 1 0 14930 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__11833_
timestamp 0
transform -1 0 14790 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__11834_
timestamp 0
transform -1 0 14810 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11835_
timestamp 0
transform -1 0 13770 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__11836_
timestamp 0
transform 1 0 13610 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__11837_
timestamp 0
transform 1 0 13550 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11838_
timestamp 0
transform 1 0 13550 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__11839_
timestamp 0
transform -1 0 13450 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11840_
timestamp 0
transform -1 0 13030 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__11841_
timestamp 0
transform 1 0 13150 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__11842_
timestamp 0
transform -1 0 13150 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__11843_
timestamp 0
transform 1 0 13230 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__11844_
timestamp 0
transform 1 0 13230 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11845_
timestamp 0
transform -1 0 13150 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11846_
timestamp 0
transform -1 0 12990 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__11847_
timestamp 0
transform -1 0 13010 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11848_
timestamp 0
transform 1 0 15350 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11849_
timestamp 0
transform -1 0 12790 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11850_
timestamp 0
transform -1 0 12630 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11851_
timestamp 0
transform 1 0 13070 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11852_
timestamp 0
transform 1 0 12910 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11853_
timestamp 0
transform 1 0 13390 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__11854_
timestamp 0
transform -1 0 13410 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11855_
timestamp 0
transform 1 0 16150 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__11856_
timestamp 0
transform 1 0 13890 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__11857_
timestamp 0
transform -1 0 14730 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__11858_
timestamp 0
transform 1 0 14370 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__11859_
timestamp 0
transform 1 0 14490 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__11860_
timestamp 0
transform -1 0 15630 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__11861_
timestamp 0
transform 1 0 15630 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11862_
timestamp 0
transform 1 0 17010 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__11863_
timestamp 0
transform 1 0 16430 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__11864_
timestamp 0
transform 1 0 15970 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__11865_
timestamp 0
transform 1 0 15910 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11866_
timestamp 0
transform 1 0 15770 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11867_
timestamp 0
transform 1 0 17070 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__11868_
timestamp 0
transform 1 0 16690 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11869_
timestamp 0
transform 1 0 16770 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__11870_
timestamp 0
transform -1 0 15810 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11871_
timestamp 0
transform -1 0 15670 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11872_
timestamp 0
transform -1 0 14910 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11873_
timestamp 0
transform 1 0 14770 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11874_
timestamp 0
transform -1 0 13650 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11875_
timestamp 0
transform -1 0 13510 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11876_
timestamp 0
transform 1 0 13230 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11877_
timestamp 0
transform 1 0 15150 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11878_
timestamp 0
transform -1 0 17070 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11879_
timestamp 0
transform 1 0 14410 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__11880_
timestamp 0
transform 1 0 14670 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__11881_
timestamp 0
transform 1 0 14450 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__11882_
timestamp 0
transform -1 0 15510 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__11883_
timestamp 0
transform -1 0 15770 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__11884_
timestamp 0
transform -1 0 15790 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11885_
timestamp 0
transform -1 0 16090 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11886_
timestamp 0
transform -1 0 16810 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11887_
timestamp 0
transform 1 0 16850 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11888_
timestamp 0
transform 1 0 16950 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11889_
timestamp 0
transform 1 0 16730 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11890_
timestamp 0
transform 1 0 16730 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11891_
timestamp 0
transform 1 0 16790 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11892_
timestamp 0
transform -1 0 16890 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11893_
timestamp 0
transform -1 0 17010 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11894_
timestamp 0
transform 1 0 16990 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11895_
timestamp 0
transform 1 0 17050 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11896_
timestamp 0
transform -1 0 15470 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11897_
timestamp 0
transform -1 0 15330 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11898_
timestamp 0
transform 1 0 13990 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11899_
timestamp 0
transform 1 0 16310 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11900_
timestamp 0
transform -1 0 16930 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__11901_
timestamp 0
transform 1 0 16930 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__11902_
timestamp 0
transform -1 0 14690 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11903_
timestamp 0
transform 1 0 14950 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11904_
timestamp 0
transform 1 0 15350 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11905_
timestamp 0
transform 1 0 15490 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11906_
timestamp 0
transform 1 0 15570 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__11907_
timestamp 0
transform 1 0 16590 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11908_
timestamp 0
transform -1 0 16550 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__11909_
timestamp 0
transform 1 0 16490 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11910_
timestamp 0
transform -1 0 16350 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11911_
timestamp 0
transform -1 0 16350 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11912_
timestamp 0
transform 1 0 16470 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11913_
timestamp 0
transform 1 0 16790 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11914_
timestamp 0
transform 1 0 16670 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11915_
timestamp 0
transform -1 0 15170 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11916_
timestamp 0
transform -1 0 15030 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11917_
timestamp 0
transform -1 0 14710 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11918_
timestamp 0
transform 1 0 12550 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11919_
timestamp 0
transform 1 0 14410 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11920_
timestamp 0
transform -1 0 16410 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__11921_
timestamp 0
transform 1 0 16590 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11922_
timestamp 0
transform -1 0 15210 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11923_
timestamp 0
transform -1 0 15210 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__11924_
timestamp 0
transform 1 0 15270 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__11925_
timestamp 0
transform -1 0 16070 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11926_
timestamp 0
transform 1 0 16070 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11927_
timestamp 0
transform 1 0 16430 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11928_
timestamp 0
transform 1 0 16170 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11929_
timestamp 0
transform -1 0 16190 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11930_
timestamp 0
transform -1 0 15930 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11931_
timestamp 0
transform 1 0 16290 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11932_
timestamp 0
transform 1 0 15930 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11933_
timestamp 0
transform 1 0 16070 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11934_
timestamp 0
transform -1 0 16650 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11935_
timestamp 0
transform 1 0 16870 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11936_
timestamp 0
transform 1 0 16890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11937_
timestamp 0
transform 1 0 16550 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11938_
timestamp 0
transform -1 0 15770 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11939_
timestamp 0
transform -1 0 15630 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11940_
timestamp 0
transform 1 0 14530 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11941_
timestamp 0
transform 1 0 12850 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11942_
timestamp 0
transform -1 0 16050 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11943_
timestamp 0
transform 1 0 16990 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11944_
timestamp 0
transform 1 0 16730 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11945_
timestamp 0
transform -1 0 16610 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11946_
timestamp 0
transform 1 0 16430 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11947_
timestamp 0
transform -1 0 15990 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11948_
timestamp 0
transform -1 0 16290 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__11949_
timestamp 0
transform -1 0 16210 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11950_
timestamp 0
transform 1 0 14550 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__11951_
timestamp 0
transform -1 0 15330 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__11952_
timestamp 0
transform 1 0 15430 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__11953_
timestamp 0
transform 1 0 15870 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__11954_
timestamp 0
transform 1 0 15730 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11955_
timestamp 0
transform 1 0 16570 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11956_
timestamp 0
transform 1 0 16390 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__11957_
timestamp 0
transform 1 0 16310 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11958_
timestamp 0
transform 1 0 15870 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11959_
timestamp 0
transform -1 0 16190 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11960_
timestamp 0
transform -1 0 16450 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11961_
timestamp 0
transform -1 0 16050 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__11962_
timestamp 0
transform 1 0 15830 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11963_
timestamp 0
transform 1 0 15610 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11964_
timestamp 0
transform 1 0 15710 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11965_
timestamp 0
transform 1 0 15910 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11966_
timestamp 0
transform -1 0 15490 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11967_
timestamp 0
transform -1 0 13250 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__11968_
timestamp 0
transform 1 0 13790 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11969_
timestamp 0
transform -1 0 14350 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11970_
timestamp 0
transform 1 0 12970 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11971_
timestamp 0
transform 1 0 14070 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11972_
timestamp 0
transform 1 0 16110 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11973_
timestamp 0
transform 1 0 16190 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__11974_
timestamp 0
transform 1 0 16270 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11975_
timestamp 0
transform 1 0 15410 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11976_
timestamp 0
transform -1 0 15710 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__11977_
timestamp 0
transform -1 0 15730 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__11978_
timestamp 0
transform -1 0 15570 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__11979_
timestamp 0
transform 1 0 15990 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__11980_
timestamp 0
transform 1 0 15370 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11981_
timestamp 0
transform -1 0 15630 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11982_
timestamp 0
transform -1 0 15250 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11983_
timestamp 0
transform 1 0 15470 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11984_
timestamp 0
transform -1 0 15850 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__11985_
timestamp 0
transform 1 0 15510 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11986_
timestamp 0
transform 1 0 15250 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11987_
timestamp 0
transform 1 0 15250 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11988_
timestamp 0
transform -1 0 15130 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11989_
timestamp 0
transform 1 0 14950 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11990_
timestamp 0
transform 1 0 14170 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__11991_
timestamp 0
transform -1 0 15750 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11992_
timestamp 0
transform -1 0 15470 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11993_
timestamp 0
transform -1 0 15890 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11994_
timestamp 0
transform -1 0 15610 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11995_
timestamp 0
transform -1 0 15330 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11996_
timestamp 0
transform -1 0 15150 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__11997_
timestamp 0
transform -1 0 15030 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__11998_
timestamp 0
transform 1 0 14670 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__11999_
timestamp 0
transform -1 0 15530 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__12000_
timestamp 0
transform -1 0 15310 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__12001_
timestamp 0
transform -1 0 15450 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12002_
timestamp 0
transform -1 0 15170 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__12003_
timestamp 0
transform -1 0 15130 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__12004_
timestamp 0
transform -1 0 15110 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__12005_
timestamp 0
transform 1 0 14790 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__12006_
timestamp 0
transform 1 0 15010 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__12007_
timestamp 0
transform -1 0 15430 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__12008_
timestamp 0
transform 1 0 14690 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__12009_
timestamp 0
transform 1 0 14830 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__12010_
timestamp 0
transform -1 0 14810 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__12011_
timestamp 0
transform -1 0 14670 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__12012_
timestamp 0
transform -1 0 14510 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__12013_
timestamp 0
transform 1 0 13450 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__12014_
timestamp 0
transform 1 0 14650 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__12015_
timestamp 0
transform 1 0 15110 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12016_
timestamp 0
transform -1 0 14770 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__12017_
timestamp 0
transform -1 0 14870 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__12018_
timestamp 0
transform -1 0 14870 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__12019_
timestamp 0
transform 1 0 14570 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__12020_
timestamp 0
transform 1 0 14510 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__12021_
timestamp 0
transform -1 0 14450 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__12022_
timestamp 0
transform 1 0 14290 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__12023_
timestamp 0
transform -1 0 14290 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__12024_
timestamp 0
transform -1 0 14530 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__12025_
timestamp 0
transform -1 0 14170 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__12026_
timestamp 0
transform -1 0 14390 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__12027_
timestamp 0
transform -1 0 14350 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__12028_
timestamp 0
transform 1 0 14950 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__12029_
timestamp 0
transform -1 0 14990 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__12030_
timestamp 0
transform -1 0 14650 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__12031_
timestamp 0
transform -1 0 14490 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__12032_
timestamp 0
transform 1 0 14390 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__12033_
timestamp 0
transform -1 0 14710 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__12034_
timestamp 0
transform -1 0 14550 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__12035_
timestamp 0
transform 1 0 14250 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__12036_
timestamp 0
transform -1 0 14070 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__12037_
timestamp 0
transform 1 0 13890 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__12038_
timestamp 0
transform -1 0 13030 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__12039_
timestamp 0
transform -1 0 14230 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__12040_
timestamp 0
transform 1 0 14670 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12041_
timestamp 0
transform 1 0 14790 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12042_
timestamp 0
transform -1 0 14430 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12043_
timestamp 0
transform -1 0 14550 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12044_
timestamp 0
transform 1 0 14210 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12045_
timestamp 0
transform -1 0 14190 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__12046_
timestamp 0
transform -1 0 14050 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__12047_
timestamp 0
transform -1 0 13930 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__12048_
timestamp 0
transform 1 0 13810 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__12049_
timestamp 0
transform -1 0 13950 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__12050_
timestamp 0
transform -1 0 14130 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__12051_
timestamp 0
transform -1 0 13670 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__12052_
timestamp 0
transform -1 0 13530 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__12053_
timestamp 0
transform 1 0 13370 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__12054_
timestamp 0
transform 1 0 12850 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12055_
timestamp 0
transform -1 0 15830 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12056_
timestamp 0
transform 1 0 16030 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12057_
timestamp 0
transform 1 0 15930 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12058_
timestamp 0
transform -1 0 16030 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12059_
timestamp 0
transform -1 0 12570 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12060_
timestamp 0
transform 1 0 12850 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12061_
timestamp 0
transform -1 0 12610 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12062_
timestamp 0
transform 1 0 16150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12063_
timestamp 0
transform 1 0 16490 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12064_
timestamp 0
transform -1 0 16630 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12065_
timestamp 0
transform -1 0 17050 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12066_
timestamp 0
transform 1 0 17030 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12067_
timestamp 0
transform 1 0 16710 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12068_
timestamp 0
transform 1 0 16670 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12069_
timestamp 0
transform -1 0 16250 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12070_
timestamp 0
transform 1 0 12850 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12071_
timestamp 0
transform 1 0 17030 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12072_
timestamp 0
transform -1 0 16910 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12073_
timestamp 0
transform 1 0 17070 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12074_
timestamp 0
transform -1 0 16930 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12075_
timestamp 0
transform -1 0 13010 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12076_
timestamp 0
transform -1 0 12730 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12077_
timestamp 0
transform -1 0 12570 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12078_
timestamp 0
transform -1 0 13150 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12079_
timestamp 0
transform 1 0 15570 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__12080_
timestamp 0
transform 1 0 16990 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12081_
timestamp 0
transform 1 0 13790 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12082_
timestamp 0
transform 1 0 13650 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12083_
timestamp 0
transform -1 0 16730 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12084_
timestamp 0
transform 1 0 16570 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12085_
timestamp 0
transform -1 0 16090 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12086_
timestamp 0
transform -1 0 16210 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12087_
timestamp 0
transform -1 0 16710 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12088_
timestamp 0
transform 1 0 16470 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12089_
timestamp 0
transform 1 0 16750 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12090_
timestamp 0
transform 1 0 16970 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12091_
timestamp 0
transform 1 0 16790 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12092_
timestamp 0
transform 1 0 16550 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12093_
timestamp 0
transform -1 0 15430 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12094_
timestamp 0
transform 1 0 16710 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12095_
timestamp 0
transform -1 0 16570 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12096_
timestamp 0
transform 1 0 16370 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12097_
timestamp 0
transform -1 0 15150 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12098_
timestamp 0
transform -1 0 15170 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12099_
timestamp 0
transform 1 0 15270 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12100_
timestamp 0
transform -1 0 15030 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12101_
timestamp 0
transform 1 0 13790 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12102_
timestamp 0
transform -1 0 13670 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12103_
timestamp 0
transform -1 0 13510 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12104_
timestamp 0
transform -1 0 12710 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12105_
timestamp 0
transform -1 0 13170 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12106_
timestamp 0
transform 1 0 15270 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12107_
timestamp 0
transform -1 0 16830 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12108_
timestamp 0
transform -1 0 15550 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12109_
timestamp 0
transform -1 0 15690 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12110_
timestamp 0
transform 1 0 16570 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12111_
timestamp 0
transform 1 0 16150 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12112_
timestamp 0
transform -1 0 16330 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12113_
timestamp 0
transform 1 0 16890 0 1 250
box -6 -8 26 248
use FILL  FILL_1__12114_
timestamp 0
transform -1 0 16470 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12115_
timestamp 0
transform 1 0 16370 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12116_
timestamp 0
transform 1 0 16930 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12117_
timestamp 0
transform -1 0 16790 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12118_
timestamp 0
transform 1 0 16530 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12119_
timestamp 0
transform 1 0 16630 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12120_
timestamp 0
transform 1 0 16470 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12121_
timestamp 0
transform -1 0 16090 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12122_
timestamp 0
transform 1 0 16310 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12123_
timestamp 0
transform -1 0 15970 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12124_
timestamp 0
transform -1 0 15690 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12125_
timestamp 0
transform 1 0 15830 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12126_
timestamp 0
transform -1 0 15550 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12127_
timestamp 0
transform -1 0 13310 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12128_
timestamp 0
transform 1 0 16170 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12129_
timestamp 0
transform 1 0 17030 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12130_
timestamp 0
transform -1 0 15010 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__12131_
timestamp 0
transform 1 0 15370 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__12132_
timestamp 0
transform -1 0 16250 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12133_
timestamp 0
transform -1 0 16810 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12134_
timestamp 0
transform 1 0 16870 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12135_
timestamp 0
transform 1 0 17010 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12136_
timestamp 0
transform 1 0 16870 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12137_
timestamp 0
transform 1 0 16910 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12138_
timestamp 0
transform 1 0 17030 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12139_
timestamp 0
transform 1 0 17050 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12140_
timestamp 0
transform 1 0 16770 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12141_
timestamp 0
transform -1 0 16550 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12142_
timestamp 0
transform 1 0 16530 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12143_
timestamp 0
transform 1 0 16690 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12144_
timestamp 0
transform 1 0 16630 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12145_
timestamp 0
transform 1 0 16890 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12146_
timestamp 0
transform 1 0 16750 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12147_
timestamp 0
transform 1 0 16850 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12148_
timestamp 0
transform 1 0 14370 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12149_
timestamp 0
transform 1 0 16390 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12150_
timestamp 0
transform -1 0 14930 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12151_
timestamp 0
transform 1 0 15030 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12152_
timestamp 0
transform -1 0 15650 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12153_
timestamp 0
transform -1 0 15870 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12154_
timestamp 0
transform -1 0 16550 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12155_
timestamp 0
transform 1 0 16650 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12156_
timestamp 0
transform 1 0 17090 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12157_
timestamp 0
transform 1 0 16930 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12158_
timestamp 0
transform 1 0 16990 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12159_
timestamp 0
transform -1 0 16870 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12160_
timestamp 0
transform 1 0 16850 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12161_
timestamp 0
transform 1 0 16710 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12162_
timestamp 0
transform 1 0 16710 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12163_
timestamp 0
transform 1 0 16990 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12164_
timestamp 0
transform -1 0 16590 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12165_
timestamp 0
transform -1 0 16570 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12166_
timestamp 0
transform -1 0 16150 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12167_
timestamp 0
transform -1 0 15350 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12168_
timestamp 0
transform 1 0 15490 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12169_
timestamp 0
transform 1 0 15210 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12170_
timestamp 0
transform 1 0 13790 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12171_
timestamp 0
transform 1 0 13970 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12172_
timestamp 0
transform 1 0 15850 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12173_
timestamp 0
transform -1 0 16130 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12174_
timestamp 0
transform -1 0 15970 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12175_
timestamp 0
transform 1 0 16090 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12176_
timestamp 0
transform 1 0 16450 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12177_
timestamp 0
transform 1 0 16290 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12178_
timestamp 0
transform 1 0 16150 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12179_
timestamp 0
transform 1 0 16230 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12180_
timestamp 0
transform -1 0 16670 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12181_
timestamp 0
transform -1 0 16530 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12182_
timestamp 0
transform -1 0 16390 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12183_
timestamp 0
transform -1 0 16270 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12184_
timestamp 0
transform -1 0 16270 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12185_
timestamp 0
transform -1 0 16010 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12186_
timestamp 0
transform -1 0 16430 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12187_
timestamp 0
transform -1 0 15470 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12188_
timestamp 0
transform 1 0 15090 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12189_
timestamp 0
transform -1 0 14950 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12190_
timestamp 0
transform -1 0 14810 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12191_
timestamp 0
transform 1 0 14070 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12192_
timestamp 0
transform 1 0 12650 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12193_
timestamp 0
transform -1 0 15970 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12194_
timestamp 0
transform 1 0 16010 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12195_
timestamp 0
transform -1 0 16130 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12196_
timestamp 0
transform -1 0 16230 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12197_
timestamp 0
transform 1 0 15650 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12198_
timestamp 0
transform -1 0 16290 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12199_
timestamp 0
transform 1 0 15910 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12200_
timestamp 0
transform -1 0 16030 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12201_
timestamp 0
transform 1 0 15390 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12202_
timestamp 0
transform 1 0 15270 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12203_
timestamp 0
transform 1 0 15110 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12204_
timestamp 0
transform -1 0 15010 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12205_
timestamp 0
transform -1 0 16410 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12206_
timestamp 0
transform -1 0 16030 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12207_
timestamp 0
transform 1 0 15710 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12208_
timestamp 0
transform 1 0 15570 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12209_
timestamp 0
transform 1 0 15330 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12210_
timestamp 0
transform -1 0 15190 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12211_
timestamp 0
transform -1 0 16270 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12212_
timestamp 0
transform -1 0 15870 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12213_
timestamp 0
transform -1 0 16110 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12214_
timestamp 0
transform -1 0 15730 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12215_
timestamp 0
transform -1 0 15050 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12216_
timestamp 0
transform -1 0 14910 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12217_
timestamp 0
transform 1 0 13130 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12218_
timestamp 0
transform 1 0 12990 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12219_
timestamp 0
transform 1 0 13970 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12220_
timestamp 0
transform -1 0 14790 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12221_
timestamp 0
transform 1 0 16150 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12222_
timestamp 0
transform 1 0 15810 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12223_
timestamp 0
transform -1 0 15770 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12224_
timestamp 0
transform -1 0 15970 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12225_
timestamp 0
transform 1 0 15470 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12226_
timestamp 0
transform 1 0 15810 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12227_
timestamp 0
transform -1 0 15810 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12228_
timestamp 0
transform -1 0 15590 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12229_
timestamp 0
transform -1 0 15430 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12230_
timestamp 0
transform -1 0 15890 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12231_
timestamp 0
transform -1 0 15710 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12232_
timestamp 0
transform -1 0 15730 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12233_
timestamp 0
transform 1 0 15530 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12234_
timestamp 0
transform -1 0 14510 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12235_
timestamp 0
transform 1 0 14650 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12236_
timestamp 0
transform -1 0 14390 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12237_
timestamp 0
transform -1 0 14250 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12238_
timestamp 0
transform 1 0 14070 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__12239_
timestamp 0
transform 1 0 14830 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12240_
timestamp 0
transform -1 0 14730 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12241_
timestamp 0
transform -1 0 14570 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12242_
timestamp 0
transform -1 0 14430 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12243_
timestamp 0
transform 1 0 16010 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12244_
timestamp 0
transform -1 0 16110 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12245_
timestamp 0
transform -1 0 15970 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12246_
timestamp 0
transform -1 0 15210 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12247_
timestamp 0
transform -1 0 14830 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12248_
timestamp 0
transform -1 0 15330 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12249_
timestamp 0
transform -1 0 15090 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12250_
timestamp 0
transform -1 0 14530 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12251_
timestamp 0
transform -1 0 15230 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12252_
timestamp 0
transform 1 0 14950 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12253_
timestamp 0
transform -1 0 14670 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12254_
timestamp 0
transform -1 0 14150 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12255_
timestamp 0
transform -1 0 13750 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12256_
timestamp 0
transform -1 0 14290 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12257_
timestamp 0
transform -1 0 13870 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12258_
timestamp 0
transform 1 0 13550 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12259_
timestamp 0
transform -1 0 13490 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12260_
timestamp 0
transform -1 0 14010 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12261_
timestamp 0
transform -1 0 14090 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12262_
timestamp 0
transform 1 0 15810 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12263_
timestamp 0
transform 1 0 14890 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12264_
timestamp 0
transform -1 0 15090 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12265_
timestamp 0
transform 1 0 14930 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12266_
timestamp 0
transform -1 0 14810 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12267_
timestamp 0
transform -1 0 14530 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12268_
timestamp 0
transform 1 0 14670 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12269_
timestamp 0
transform 1 0 14630 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12270_
timestamp 0
transform 1 0 14270 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12271_
timestamp 0
transform -1 0 13990 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12272_
timestamp 0
transform 1 0 14110 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12273_
timestamp 0
transform -1 0 13850 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12274_
timestamp 0
transform 1 0 13390 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12275_
timestamp 0
transform -1 0 14210 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12276_
timestamp 0
transform 1 0 14310 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12277_
timestamp 0
transform -1 0 14430 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12278_
timestamp 0
transform 1 0 14610 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12279_
timestamp 0
transform -1 0 14470 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12280_
timestamp 0
transform 1 0 15670 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12281_
timestamp 0
transform -1 0 15590 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12282_
timestamp 0
transform 1 0 15370 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12283_
timestamp 0
transform -1 0 14770 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12284_
timestamp 0
transform 1 0 14490 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12285_
timestamp 0
transform -1 0 14590 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12286_
timestamp 0
transform 1 0 14410 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12287_
timestamp 0
transform -1 0 14250 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12288_
timestamp 0
transform 1 0 14370 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12289_
timestamp 0
transform -1 0 14090 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12290_
timestamp 0
transform 1 0 14270 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12291_
timestamp 0
transform -1 0 13810 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12292_
timestamp 0
transform 1 0 13950 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12293_
timestamp 0
transform -1 0 13690 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12294_
timestamp 0
transform 1 0 13490 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12295_
timestamp 0
transform -1 0 13130 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12296_
timestamp 0
transform -1 0 14410 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12297_
timestamp 0
transform -1 0 14150 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12298_
timestamp 0
transform 1 0 14270 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12299_
timestamp 0
transform 1 0 14150 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12300_
timestamp 0
transform 1 0 14270 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12301_
timestamp 0
transform -1 0 14150 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12302_
timestamp 0
transform -1 0 14010 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12303_
timestamp 0
transform -1 0 13850 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12304_
timestamp 0
transform -1 0 13710 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12305_
timestamp 0
transform -1 0 11890 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12306_
timestamp 0
transform 1 0 10690 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12307_
timestamp 0
transform 1 0 10830 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12308_
timestamp 0
transform -1 0 10950 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12309_
timestamp 0
transform 1 0 11070 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12310_
timestamp 0
transform 1 0 11190 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12311_
timestamp 0
transform 1 0 11510 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12312_
timestamp 0
transform 1 0 11270 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12313_
timestamp 0
transform -1 0 11270 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12314_
timestamp 0
transform -1 0 10950 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12315_
timestamp 0
transform 1 0 10730 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12316_
timestamp 0
transform -1 0 10610 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12317_
timestamp 0
transform -1 0 10050 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12318_
timestamp 0
transform -1 0 10330 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12319_
timestamp 0
transform -1 0 10190 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12320_
timestamp 0
transform 1 0 10250 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12321_
timestamp 0
transform -1 0 10210 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12322_
timestamp 0
transform -1 0 10110 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12323_
timestamp 0
transform -1 0 10090 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12324_
timestamp 0
transform -1 0 10870 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12325_
timestamp 0
transform -1 0 10730 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12326_
timestamp 0
transform -1 0 10990 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12327_
timestamp 0
transform 1 0 11090 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12328_
timestamp 0
transform 1 0 10450 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12329_
timestamp 0
transform 1 0 10550 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12330_
timestamp 0
transform -1 0 12470 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12331_
timestamp 0
transform -1 0 11530 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12332_
timestamp 0
transform -1 0 11670 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12333_
timestamp 0
transform 1 0 11230 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12334_
timestamp 0
transform -1 0 11090 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12335_
timestamp 0
transform 1 0 10950 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12336_
timestamp 0
transform -1 0 10850 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12337_
timestamp 0
transform -1 0 10350 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12338_
timestamp 0
transform -1 0 10410 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12339_
timestamp 0
transform 1 0 10250 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12340_
timestamp 0
transform 1 0 10090 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12341_
timestamp 0
transform 1 0 11150 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12342_
timestamp 0
transform -1 0 10650 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12343_
timestamp 0
transform 1 0 11010 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12344_
timestamp 0
transform 1 0 11650 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12345_
timestamp 0
transform 1 0 12610 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12346_
timestamp 0
transform -1 0 12330 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12347_
timestamp 0
transform 1 0 11930 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12348_
timestamp 0
transform -1 0 12030 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12349_
timestamp 0
transform 1 0 11530 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12350_
timestamp 0
transform -1 0 11430 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12351_
timestamp 0
transform -1 0 10630 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12352_
timestamp 0
transform -1 0 10750 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12353_
timestamp 0
transform 1 0 11110 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12354_
timestamp 0
transform 1 0 11130 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12355_
timestamp 0
transform -1 0 11050 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12356_
timestamp 0
transform 1 0 10650 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12357_
timestamp 0
transform -1 0 9950 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12358_
timestamp 0
transform -1 0 10470 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12359_
timestamp 0
transform -1 0 10330 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12360_
timestamp 0
transform -1 0 10030 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12361_
timestamp 0
transform -1 0 9690 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12362_
timestamp 0
transform -1 0 9830 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12363_
timestamp 0
transform -1 0 9770 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12364_
timestamp 0
transform -1 0 10890 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12365_
timestamp 0
transform 1 0 9950 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12366_
timestamp 0
transform 1 0 10110 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12367_
timestamp 0
transform 1 0 10250 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12368_
timestamp 0
transform -1 0 9550 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12369_
timestamp 0
transform -1 0 9930 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12370_
timestamp 0
transform 1 0 12670 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12371_
timestamp 0
transform 1 0 12030 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12372_
timestamp 0
transform 1 0 12170 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12373_
timestamp 0
transform -1 0 12350 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12374_
timestamp 0
transform -1 0 10190 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12375_
timestamp 0
transform -1 0 10230 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12376_
timestamp 0
transform 1 0 10270 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12377_
timestamp 0
transform 1 0 9890 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12378_
timestamp 0
transform -1 0 9290 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12379_
timestamp 0
transform -1 0 9410 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12380_
timestamp 0
transform -1 0 9510 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12381_
timestamp 0
transform -1 0 9350 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12382_
timestamp 0
transform 1 0 10650 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12383_
timestamp 0
transform 1 0 9670 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12384_
timestamp 0
transform 1 0 9770 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12385_
timestamp 0
transform 1 0 10030 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12386_
timestamp 0
transform -1 0 9930 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12387_
timestamp 0
transform -1 0 9750 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12388_
timestamp 0
transform -1 0 12490 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12389_
timestamp 0
transform 1 0 12470 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12390_
timestamp 0
transform 1 0 12190 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12391_
timestamp 0
transform -1 0 12330 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12392_
timestamp 0
transform -1 0 12090 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12393_
timestamp 0
transform 1 0 11010 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12394_
timestamp 0
transform -1 0 10870 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12395_
timestamp 0
transform 1 0 10850 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12396_
timestamp 0
transform -1 0 10030 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12397_
timestamp 0
transform -1 0 10050 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12398_
timestamp 0
transform -1 0 9910 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12399_
timestamp 0
transform -1 0 10170 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12400_
timestamp 0
transform 1 0 10270 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12401_
timestamp 0
transform 1 0 10370 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12402_
timestamp 0
transform 1 0 10730 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12403_
timestamp 0
transform 1 0 11310 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12404_
timestamp 0
transform -1 0 10550 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12405_
timestamp 0
transform -1 0 10410 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12406_
timestamp 0
transform 1 0 10650 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12407_
timestamp 0
transform -1 0 10810 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12408_
timestamp 0
transform -1 0 10610 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12409_
timestamp 0
transform -1 0 10930 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12410_
timestamp 0
transform -1 0 10470 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12411_
timestamp 0
transform 1 0 10590 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12412_
timestamp 0
transform -1 0 10470 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12413_
timestamp 0
transform 1 0 10490 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12414_
timestamp 0
transform 1 0 11130 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12415_
timestamp 0
transform 1 0 11870 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12416_
timestamp 0
transform -1 0 11790 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12417_
timestamp 0
transform -1 0 11650 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12418_
timestamp 0
transform 1 0 11630 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12419_
timestamp 0
transform 1 0 11790 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12420_
timestamp 0
transform -1 0 11750 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12421_
timestamp 0
transform -1 0 10330 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12422_
timestamp 0
transform -1 0 10330 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12423_
timestamp 0
transform 1 0 10170 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12424_
timestamp 0
transform 1 0 10010 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12425_
timestamp 0
transform 1 0 10150 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12426_
timestamp 0
transform 1 0 11250 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12427_
timestamp 0
transform -1 0 11090 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12428_
timestamp 0
transform -1 0 10970 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12429_
timestamp 0
transform 1 0 10970 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12430_
timestamp 0
transform -1 0 11650 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12431_
timestamp 0
transform -1 0 11750 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12432_
timestamp 0
transform -1 0 11610 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12433_
timestamp 0
transform -1 0 11230 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12434_
timestamp 0
transform -1 0 11230 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12435_
timestamp 0
transform 1 0 11370 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12436_
timestamp 0
transform -1 0 11350 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12437_
timestamp 0
transform -1 0 11790 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12438_
timestamp 0
transform 1 0 11490 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12439_
timestamp 0
transform -1 0 11350 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12440_
timestamp 0
transform -1 0 11390 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12441_
timestamp 0
transform 1 0 11470 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12442_
timestamp 0
transform -1 0 12150 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12443_
timestamp 0
transform 1 0 12190 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12444_
timestamp 0
transform -1 0 12010 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12445_
timestamp 0
transform 1 0 12370 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12446_
timestamp 0
transform -1 0 12090 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12447_
timestamp 0
transform -1 0 12030 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12448_
timestamp 0
transform -1 0 11930 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12449_
timestamp 0
transform 1 0 12190 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12450_
timestamp 0
transform 1 0 12230 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__12451_
timestamp 0
transform 1 0 12030 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__12452_
timestamp 0
transform 1 0 11770 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__12453_
timestamp 0
transform -1 0 11690 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__12454_
timestamp 0
transform 1 0 11810 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__12455_
timestamp 0
transform -1 0 13870 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12456_
timestamp 0
transform -1 0 13990 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12457_
timestamp 0
transform -1 0 13950 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12458_
timestamp 0
transform -1 0 14070 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12459_
timestamp 0
transform 1 0 14030 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12460_
timestamp 0
transform -1 0 11710 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__12461_
timestamp 0
transform 1 0 13990 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12462_
timestamp 0
transform 1 0 13850 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12463_
timestamp 0
transform 1 0 14130 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12464_
timestamp 0
transform 1 0 13710 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12465_
timestamp 0
transform -1 0 13550 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12466_
timestamp 0
transform 1 0 12290 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12467_
timestamp 0
transform -1 0 14810 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12468_
timestamp 0
transform 1 0 14250 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12469_
timestamp 0
transform 1 0 14330 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12470_
timestamp 0
transform 1 0 13930 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12471_
timestamp 0
transform 1 0 12170 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12472_
timestamp 0
transform 1 0 16410 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__12473_
timestamp 0
transform -1 0 16570 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__12474_
timestamp 0
transform 1 0 15170 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__12475_
timestamp 0
transform -1 0 15550 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__12476_
timestamp 0
transform 1 0 13550 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12477_
timestamp 0
transform -1 0 13710 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12478_
timestamp 0
transform 1 0 13610 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12479_
timestamp 0
transform -1 0 13770 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__12480_
timestamp 0
transform -1 0 12890 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12481_
timestamp 0
transform 1 0 12990 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12482_
timestamp 0
transform 1 0 13650 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12483_
timestamp 0
transform 1 0 13510 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12484_
timestamp 0
transform -1 0 14010 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__12485_
timestamp 0
transform -1 0 14150 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__12486_
timestamp 0
transform 1 0 14150 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12487_
timestamp 0
transform -1 0 14290 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12488_
timestamp 0
transform -1 0 13910 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__12489_
timestamp 0
transform -1 0 13750 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__12490_
timestamp 0
transform 1 0 13590 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__12491_
timestamp 0
transform -1 0 14050 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12492_
timestamp 0
transform 1 0 13390 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__12493_
timestamp 0
transform -1 0 13550 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__12494_
timestamp 0
transform -1 0 14470 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12495_
timestamp 0
transform 1 0 14070 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12496_
timestamp 0
transform -1 0 14750 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12497_
timestamp 0
transform 1 0 14590 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12498_
timestamp 0
transform 1 0 16350 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12499_
timestamp 0
transform -1 0 16610 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12500_
timestamp 0
transform 1 0 16510 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12501_
timestamp 0
transform -1 0 16650 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12502_
timestamp 0
transform -1 0 13330 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12503_
timestamp 0
transform -1 0 13470 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12504_
timestamp 0
transform 1 0 13550 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12505_
timestamp 0
transform -1 0 13710 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12506_
timestamp 0
transform -1 0 12090 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12507_
timestamp 0
transform -1 0 12230 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12508_
timestamp 0
transform -1 0 11790 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12509_
timestamp 0
transform -1 0 11930 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12510_
timestamp 0
transform 1 0 12450 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12511_
timestamp 0
transform 1 0 12310 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__12512_
timestamp 0
transform 1 0 11870 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12513_
timestamp 0
transform -1 0 11950 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__12514_
timestamp 0
transform 1 0 12050 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12515_
timestamp 0
transform -1 0 12310 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12516_
timestamp 0
transform 1 0 12150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12517_
timestamp 0
transform 1 0 11670 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12518_
timestamp 0
transform -1 0 12150 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12519_
timestamp 0
transform 1 0 11990 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12520_
timestamp 0
transform 1 0 10990 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12521_
timestamp 0
transform -1 0 11150 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__12522_
timestamp 0
transform 1 0 11390 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12523_
timestamp 0
transform -1 0 11550 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__12524_
timestamp 0
transform -1 0 9410 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12525_
timestamp 0
transform -1 0 9530 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__12526_
timestamp 0
transform -1 0 9650 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12527_
timestamp 0
transform -1 0 9770 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__12528_
timestamp 0
transform 1 0 11350 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12529_
timestamp 0
transform -1 0 11750 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__12530_
timestamp 0
transform -1 0 11590 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12531_
timestamp 0
transform -1 0 11750 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__12532_
timestamp 0
transform 1 0 11170 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12533_
timestamp 0
transform 1 0 11030 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12534_
timestamp 0
transform 1 0 10790 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12535_
timestamp 0
transform -1 0 10670 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__12616_
timestamp 0
transform 1 0 11270 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12617_
timestamp 0
transform -1 0 11390 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12618_
timestamp 0
transform 1 0 12350 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12619_
timestamp 0
transform 1 0 11490 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12620_
timestamp 0
transform -1 0 11090 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12621_
timestamp 0
transform -1 0 10830 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12622_
timestamp 0
transform 1 0 10930 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12623_
timestamp 0
transform -1 0 11050 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12624_
timestamp 0
transform -1 0 11530 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12625_
timestamp 0
transform -1 0 11710 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12626_
timestamp 0
transform -1 0 11550 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12627_
timestamp 0
transform -1 0 10610 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__12628_
timestamp 0
transform -1 0 11510 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12629_
timestamp 0
transform 1 0 11330 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12630_
timestamp 0
transform -1 0 11210 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12631_
timestamp 0
transform 1 0 11190 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12632_
timestamp 0
transform 1 0 11150 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12633_
timestamp 0
transform 1 0 11630 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12634_
timestamp 0
transform -1 0 11150 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12635_
timestamp 0
transform -1 0 11290 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12636_
timestamp 0
transform -1 0 11630 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12637_
timestamp 0
transform -1 0 11810 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12638_
timestamp 0
transform 1 0 11630 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12639_
timestamp 0
transform -1 0 11250 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12640_
timestamp 0
transform -1 0 11650 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__12641_
timestamp 0
transform -1 0 11310 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12642_
timestamp 0
transform 1 0 10950 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__12643_
timestamp 0
transform -1 0 11310 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__12644_
timestamp 0
transform -1 0 11010 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__12645_
timestamp 0
transform -1 0 11150 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12646_
timestamp 0
transform -1 0 11530 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12647_
timestamp 0
transform 1 0 11370 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12648_
timestamp 0
transform 1 0 11070 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12649_
timestamp 0
transform 1 0 11410 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12650_
timestamp 0
transform -1 0 10930 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12651_
timestamp 0
transform -1 0 10450 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__12652_
timestamp 0
transform 1 0 11130 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__12653_
timestamp 0
transform 1 0 11190 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12654_
timestamp 0
transform -1 0 11490 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__12655_
timestamp 0
transform 1 0 11190 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__12656_
timestamp 0
transform -1 0 11350 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__12657_
timestamp 0
transform 1 0 11330 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12658_
timestamp 0
transform 1 0 12090 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12659_
timestamp 0
transform -1 0 11390 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12660_
timestamp 0
transform -1 0 12510 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12661_
timestamp 0
transform 1 0 12130 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__12662_
timestamp 0
transform -1 0 12370 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__12663_
timestamp 0
transform -1 0 11990 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__12664_
timestamp 0
transform -1 0 12090 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__12665_
timestamp 0
transform 1 0 11950 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__12666_
timestamp 0
transform -1 0 11830 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__12667_
timestamp 0
transform -1 0 12010 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12668_
timestamp 0
transform -1 0 13330 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__12669_
timestamp 0
transform -1 0 17010 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12670_
timestamp 0
transform 1 0 16030 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__12671_
timestamp 0
transform 1 0 16690 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12672_
timestamp 0
transform -1 0 16550 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12673_
timestamp 0
transform -1 0 16670 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12674_
timestamp 0
transform 1 0 16870 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12675_
timestamp 0
transform 1 0 17070 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__12676_
timestamp 0
transform 1 0 16910 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__12677_
timestamp 0
transform -1 0 16590 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__12678_
timestamp 0
transform 1 0 16430 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__12679_
timestamp 0
transform -1 0 16170 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__12680_
timestamp 0
transform -1 0 16310 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__12681_
timestamp 0
transform 1 0 15930 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__12682_
timestamp 0
transform 1 0 16690 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__12683_
timestamp 0
transform 1 0 16530 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__12684_
timestamp 0
transform 1 0 16350 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__12685_
timestamp 0
transform -1 0 16250 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__12686_
timestamp 0
transform -1 0 13110 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12687_
timestamp 0
transform -1 0 13250 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12688_
timestamp 0
transform -1 0 12650 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12689_
timestamp 0
transform -1 0 14910 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__12690_
timestamp 0
transform -1 0 12770 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__12691_
timestamp 0
transform 1 0 12890 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__12692_
timestamp 0
transform -1 0 12510 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12693_
timestamp 0
transform 1 0 12050 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12694_
timestamp 0
transform -1 0 11570 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12695_
timestamp 0
transform 1 0 11350 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__12696_
timestamp 0
transform -1 0 12870 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12697_
timestamp 0
transform -1 0 16050 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12698_
timestamp 0
transform -1 0 16410 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__12699_
timestamp 0
transform -1 0 15890 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12700_
timestamp 0
transform 1 0 16170 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__12701_
timestamp 0
transform 1 0 16030 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__12702_
timestamp 0
transform -1 0 15890 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__12703_
timestamp 0
transform -1 0 15790 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__12704_
timestamp 0
transform -1 0 16530 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__12705_
timestamp 0
transform -1 0 16210 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__12706_
timestamp 0
transform -1 0 15630 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__12707_
timestamp 0
transform 1 0 14470 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__12708_
timestamp 0
transform 1 0 14450 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12709_
timestamp 0
transform 1 0 16370 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12710_
timestamp 0
transform 1 0 15750 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12711_
timestamp 0
transform 1 0 15890 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12712_
timestamp 0
transform -1 0 16670 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__12713_
timestamp 0
transform 1 0 16810 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12714_
timestamp 0
transform 1 0 16650 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12715_
timestamp 0
transform 1 0 16310 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12716_
timestamp 0
transform 1 0 17030 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__12717_
timestamp 0
transform 1 0 17070 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12718_
timestamp 0
transform 1 0 16930 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12719_
timestamp 0
transform 1 0 16690 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__12720_
timestamp 0
transform 1 0 16790 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__12721_
timestamp 0
transform 1 0 16990 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__12722_
timestamp 0
transform 1 0 16930 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12723_
timestamp 0
transform 1 0 16530 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12724_
timestamp 0
transform -1 0 14430 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12725_
timestamp 0
transform -1 0 15770 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12726_
timestamp 0
transform -1 0 16970 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12727_
timestamp 0
transform 1 0 16370 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12728_
timestamp 0
transform -1 0 16490 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__12729_
timestamp 0
transform 1 0 16730 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__12730_
timestamp 0
transform -1 0 16810 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12731_
timestamp 0
transform -1 0 16210 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12732_
timestamp 0
transform 1 0 14110 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__12733_
timestamp 0
transform -1 0 13910 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12734_
timestamp 0
transform -1 0 13810 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12735_
timestamp 0
transform -1 0 14070 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12736_
timestamp 0
transform -1 0 13650 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12737_
timestamp 0
transform -1 0 13570 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__12738_
timestamp 0
transform -1 0 13030 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12739_
timestamp 0
transform -1 0 12770 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12740_
timestamp 0
transform -1 0 11510 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__12741_
timestamp 0
transform -1 0 9010 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12742_
timestamp 0
transform 1 0 9230 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__12743_
timestamp 0
transform 1 0 9110 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__12744_
timestamp 0
transform -1 0 11730 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12745_
timestamp 0
transform -1 0 13370 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12746_
timestamp 0
transform 1 0 15550 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12747_
timestamp 0
transform -1 0 15730 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12748_
timestamp 0
transform -1 0 15690 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__12749_
timestamp 0
transform -1 0 15390 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__12750_
timestamp 0
transform 1 0 15490 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__12751_
timestamp 0
transform 1 0 15230 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__12752_
timestamp 0
transform -1 0 13830 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__12753_
timestamp 0
transform 1 0 13690 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__12754_
timestamp 0
transform 1 0 14190 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12755_
timestamp 0
transform -1 0 14590 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12756_
timestamp 0
transform 1 0 14290 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__12757_
timestamp 0
transform -1 0 13450 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12758_
timestamp 0
transform -1 0 13610 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12759_
timestamp 0
transform -1 0 13210 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12760_
timestamp 0
transform -1 0 12910 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12761_
timestamp 0
transform -1 0 12910 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12762_
timestamp 0
transform -1 0 12390 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12763_
timestamp 0
transform 1 0 13050 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12764_
timestamp 0
transform -1 0 12230 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12765_
timestamp 0
transform 1 0 12490 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12766_
timestamp 0
transform -1 0 12250 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12767_
timestamp 0
transform -1 0 12090 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12768_
timestamp 0
transform 1 0 11810 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12769_
timestamp 0
transform 1 0 12370 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12770_
timestamp 0
transform 1 0 13290 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12771_
timestamp 0
transform -1 0 12770 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12772_
timestamp 0
transform 1 0 14970 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12773_
timestamp 0
transform -1 0 13990 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__12774_
timestamp 0
transform 1 0 15150 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12775_
timestamp 0
transform -1 0 15350 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12776_
timestamp 0
transform 1 0 15450 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12777_
timestamp 0
transform 1 0 15630 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12778_
timestamp 0
transform 1 0 15490 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12779_
timestamp 0
transform 1 0 17010 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12780_
timestamp 0
transform 1 0 16810 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12781_
timestamp 0
transform 1 0 16470 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12782_
timestamp 0
transform 1 0 15230 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12783_
timestamp 0
transform -1 0 13190 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12784_
timestamp 0
transform -1 0 12990 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12785_
timestamp 0
transform -1 0 13250 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12786_
timestamp 0
transform 1 0 13070 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12787_
timestamp 0
transform -1 0 13230 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12788_
timestamp 0
transform 1 0 13350 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12789_
timestamp 0
transform -1 0 12990 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12790_
timestamp 0
transform -1 0 12870 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12791_
timestamp 0
transform -1 0 12610 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12792_
timestamp 0
transform -1 0 12470 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12793_
timestamp 0
transform 1 0 11910 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12794_
timestamp 0
transform -1 0 13090 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12795_
timestamp 0
transform -1 0 14070 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12796_
timestamp 0
transform 1 0 14970 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12797_
timestamp 0
transform 1 0 15390 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12798_
timestamp 0
transform 1 0 15230 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12799_
timestamp 0
transform -1 0 15390 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12800_
timestamp 0
transform -1 0 15390 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12801_
timestamp 0
transform 1 0 15590 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12802_
timestamp 0
transform -1 0 15110 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12803_
timestamp 0
transform -1 0 13490 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12804_
timestamp 0
transform -1 0 13650 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12805_
timestamp 0
transform -1 0 13490 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12806_
timestamp 0
transform 1 0 13930 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12807_
timestamp 0
transform 1 0 12790 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__12808_
timestamp 0
transform 1 0 13390 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12809_
timestamp 0
transform 1 0 13510 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12810_
timestamp 0
transform 1 0 13630 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12811_
timestamp 0
transform 1 0 13790 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12812_
timestamp 0
transform 1 0 12730 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12813_
timestamp 0
transform -1 0 12870 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12814_
timestamp 0
transform 1 0 12690 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12815_
timestamp 0
transform 1 0 11970 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12816_
timestamp 0
transform -1 0 12610 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12817_
timestamp 0
transform -1 0 14550 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__12818_
timestamp 0
transform 1 0 13330 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12819_
timestamp 0
transform 1 0 15650 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12820_
timestamp 0
transform 1 0 15810 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12821_
timestamp 0
transform 1 0 15670 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12822_
timestamp 0
transform 1 0 16390 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12823_
timestamp 0
transform -1 0 15530 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12824_
timestamp 0
transform -1 0 13790 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12825_
timestamp 0
transform 1 0 13590 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__12826_
timestamp 0
transform -1 0 14090 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12827_
timestamp 0
transform -1 0 13570 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__12828_
timestamp 0
transform -1 0 13270 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__12829_
timestamp 0
transform -1 0 13110 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__12830_
timestamp 0
transform -1 0 13310 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12831_
timestamp 0
transform 1 0 13110 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12832_
timestamp 0
transform -1 0 12570 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12833_
timestamp 0
transform -1 0 12430 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12834_
timestamp 0
transform -1 0 12270 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12835_
timestamp 0
transform 1 0 11490 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12836_
timestamp 0
transform 1 0 12150 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12837_
timestamp 0
transform -1 0 13550 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12838_
timestamp 0
transform 1 0 13390 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__12839_
timestamp 0
transform -1 0 15550 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12840_
timestamp 0
transform 1 0 15330 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12841_
timestamp 0
transform -1 0 15330 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__12842_
timestamp 0
transform -1 0 13490 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12843_
timestamp 0
transform -1 0 14110 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12844_
timestamp 0
transform 1 0 13930 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12845_
timestamp 0
transform 1 0 13810 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12846_
timestamp 0
transform -1 0 13270 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12847_
timestamp 0
transform -1 0 13690 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12848_
timestamp 0
transform 1 0 13950 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12849_
timestamp 0
transform -1 0 13550 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12850_
timestamp 0
transform -1 0 12750 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12851_
timestamp 0
transform -1 0 12970 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__12852_
timestamp 0
transform 1 0 13010 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12853_
timestamp 0
transform 1 0 12870 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12854_
timestamp 0
transform -1 0 13010 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12855_
timestamp 0
transform -1 0 12430 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12856_
timestamp 0
transform -1 0 12470 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12857_
timestamp 0
transform 1 0 12270 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12858_
timestamp 0
transform 1 0 11870 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12859_
timestamp 0
transform 1 0 13390 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12860_
timestamp 0
transform -1 0 13330 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12861_
timestamp 0
transform -1 0 13190 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12862_
timestamp 0
transform 1 0 13130 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12863_
timestamp 0
transform 1 0 13030 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12864_
timestamp 0
transform -1 0 13130 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12865_
timestamp 0
transform -1 0 13930 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12866_
timestamp 0
transform 1 0 13690 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__12867_
timestamp 0
transform 1 0 15210 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12868_
timestamp 0
transform -1 0 15350 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12869_
timestamp 0
transform -1 0 15250 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12870_
timestamp 0
transform 1 0 14710 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12871_
timestamp 0
transform -1 0 13790 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12872_
timestamp 0
transform -1 0 14330 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12873_
timestamp 0
transform 1 0 13610 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12874_
timestamp 0
transform 1 0 13750 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12875_
timestamp 0
transform -1 0 13650 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12876_
timestamp 0
transform 1 0 14030 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12877_
timestamp 0
transform 1 0 14190 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12878_
timestamp 0
transform -1 0 13910 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12879_
timestamp 0
transform -1 0 13010 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12880_
timestamp 0
transform -1 0 12890 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12881_
timestamp 0
transform 1 0 12970 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12882_
timestamp 0
transform 1 0 12590 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12883_
timestamp 0
transform -1 0 12290 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12884_
timestamp 0
transform -1 0 12070 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12885_
timestamp 0
transform -1 0 11970 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12886_
timestamp 0
transform -1 0 12130 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12887_
timestamp 0
transform 1 0 11970 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12888_
timestamp 0
transform -1 0 11430 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12889_
timestamp 0
transform 1 0 12850 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12890_
timestamp 0
transform -1 0 12590 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12891_
timestamp 0
transform -1 0 12710 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12892_
timestamp 0
transform 1 0 13570 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12893_
timestamp 0
transform -1 0 13850 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12894_
timestamp 0
transform 1 0 14670 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12895_
timestamp 0
transform -1 0 13690 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12896_
timestamp 0
transform 1 0 13990 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12897_
timestamp 0
transform 1 0 14150 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12898_
timestamp 0
transform 1 0 13990 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12899_
timestamp 0
transform -1 0 13450 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12900_
timestamp 0
transform -1 0 13850 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12901_
timestamp 0
transform -1 0 13710 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12902_
timestamp 0
transform -1 0 13570 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12903_
timestamp 0
transform -1 0 13370 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12904_
timestamp 0
transform -1 0 12530 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12905_
timestamp 0
transform -1 0 12370 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12906_
timestamp 0
transform -1 0 12230 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12907_
timestamp 0
transform 1 0 11770 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12908_
timestamp 0
transform 1 0 13570 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12909_
timestamp 0
transform -1 0 13450 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12910_
timestamp 0
transform 1 0 13270 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12911_
timestamp 0
transform -1 0 13310 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12912_
timestamp 0
transform 1 0 13130 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12913_
timestamp 0
transform -1 0 13350 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12914_
timestamp 0
transform 1 0 13210 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12915_
timestamp 0
transform 1 0 14250 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12916_
timestamp 0
transform 1 0 14010 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12917_
timestamp 0
transform 1 0 14670 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12918_
timestamp 0
transform 1 0 14950 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12919_
timestamp 0
transform -1 0 14530 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12920_
timestamp 0
transform 1 0 14790 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12921_
timestamp 0
transform 1 0 14550 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12922_
timestamp 0
transform 1 0 14390 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12923_
timestamp 0
transform 1 0 14370 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12924_
timestamp 0
transform 1 0 14510 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12925_
timestamp 0
transform -1 0 14130 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__12926_
timestamp 0
transform -1 0 13530 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12927_
timestamp 0
transform -1 0 12090 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12928_
timestamp 0
transform -1 0 12230 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12929_
timestamp 0
transform -1 0 11930 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12930_
timestamp 0
transform 1 0 11050 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__12931_
timestamp 0
transform 1 0 15070 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12932_
timestamp 0
transform -1 0 15210 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12933_
timestamp 0
transform -1 0 15110 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12934_
timestamp 0
transform 1 0 14930 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12935_
timestamp 0
transform 1 0 14790 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12936_
timestamp 0
transform -1 0 13990 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12937_
timestamp 0
transform 1 0 15190 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12938_
timestamp 0
transform -1 0 14530 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12939_
timestamp 0
transform 1 0 14390 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12940_
timestamp 0
transform 1 0 14690 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12941_
timestamp 0
transform -1 0 13830 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12942_
timestamp 0
transform -1 0 14130 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12943_
timestamp 0
transform -1 0 14250 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12944_
timestamp 0
transform -1 0 12910 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12945_
timestamp 0
transform -1 0 14270 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__12946_
timestamp 0
transform -1 0 13190 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12947_
timestamp 0
transform -1 0 13090 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12948_
timestamp 0
transform -1 0 12930 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12949_
timestamp 0
transform -1 0 12770 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12950_
timestamp 0
transform -1 0 13030 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12951_
timestamp 0
transform -1 0 12630 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12952_
timestamp 0
transform -1 0 12530 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12953_
timestamp 0
transform -1 0 12370 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12954_
timestamp 0
transform 1 0 11750 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12955_
timestamp 0
transform 1 0 11930 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__12956_
timestamp 0
transform -1 0 12830 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12957_
timestamp 0
transform 1 0 15090 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12958_
timestamp 0
transform 1 0 15450 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12959_
timestamp 0
transform -1 0 14870 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12960_
timestamp 0
transform -1 0 14830 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__12961_
timestamp 0
transform 1 0 13790 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12962_
timestamp 0
transform 1 0 13890 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12963_
timestamp 0
transform -1 0 13710 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__12964_
timestamp 0
transform -1 0 13690 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12965_
timestamp 0
transform 1 0 13170 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__12966_
timestamp 0
transform -1 0 12830 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__12967_
timestamp 0
transform 1 0 12650 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__12968_
timestamp 0
transform -1 0 13050 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__12969_
timestamp 0
transform -1 0 12670 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__12970_
timestamp 0
transform 1 0 12230 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__12971_
timestamp 0
transform -1 0 12910 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12972_
timestamp 0
transform 1 0 15710 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12973_
timestamp 0
transform -1 0 15850 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12974_
timestamp 0
transform -1 0 15970 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12975_
timestamp 0
transform 1 0 16270 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12976_
timestamp 0
transform 1 0 14050 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__12977_
timestamp 0
transform -1 0 14070 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__12978_
timestamp 0
transform 1 0 14170 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__12979_
timestamp 0
transform -1 0 16130 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12980_
timestamp 0
transform -1 0 14450 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12981_
timestamp 0
transform 1 0 14550 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12982_
timestamp 0
transform -1 0 14750 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12983_
timestamp 0
transform -1 0 14870 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12984_
timestamp 0
transform 1 0 16210 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12985_
timestamp 0
transform -1 0 16410 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12986_
timestamp 0
transform 1 0 16630 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__12987_
timestamp 0
transform -1 0 15810 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__12988_
timestamp 0
transform -1 0 15850 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12989_
timestamp 0
transform 1 0 16090 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12990_
timestamp 0
transform 1 0 15970 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__12991_
timestamp 0
transform 1 0 16030 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12992_
timestamp 0
transform -1 0 15790 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12993_
timestamp 0
transform -1 0 15630 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12994_
timestamp 0
transform 1 0 12350 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__12995_
timestamp 0
transform -1 0 15930 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__12996_
timestamp 0
transform -1 0 15110 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12997_
timestamp 0
transform -1 0 15250 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__12998_
timestamp 0
transform -1 0 15470 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__12999_
timestamp 0
transform 1 0 15190 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13000_
timestamp 0
transform -1 0 16470 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13001_
timestamp 0
transform 1 0 16590 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13002_
timestamp 0
transform 1 0 14390 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13003_
timestamp 0
transform 1 0 14230 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13004_
timestamp 0
transform 1 0 16030 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13005_
timestamp 0
transform -1 0 14210 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13006_
timestamp 0
transform -1 0 14350 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13007_
timestamp 0
transform 1 0 16430 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13008_
timestamp 0
transform 1 0 16290 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13009_
timestamp 0
transform 1 0 16450 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13010_
timestamp 0
transform -1 0 16990 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13011_
timestamp 0
transform 1 0 16130 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13012_
timestamp 0
transform -1 0 16710 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13013_
timestamp 0
transform 1 0 16510 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13014_
timestamp 0
transform -1 0 16190 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13015_
timestamp 0
transform 1 0 15910 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13016_
timestamp 0
transform -1 0 16330 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13017_
timestamp 0
transform -1 0 15770 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13018_
timestamp 0
transform 1 0 15630 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13019_
timestamp 0
transform -1 0 15490 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13020_
timestamp 0
transform 1 0 14390 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13021_
timestamp 0
transform -1 0 12490 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13022_
timestamp 0
transform -1 0 12270 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13023_
timestamp 0
transform 1 0 16030 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13024_
timestamp 0
transform 1 0 16630 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13025_
timestamp 0
transform 1 0 15030 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13026_
timestamp 0
transform 1 0 14890 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13027_
timestamp 0
transform 1 0 16110 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13028_
timestamp 0
transform 1 0 15970 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13029_
timestamp 0
transform -1 0 16190 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13030_
timestamp 0
transform 1 0 16330 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13031_
timestamp 0
transform -1 0 16210 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13032_
timestamp 0
transform -1 0 16190 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13033_
timestamp 0
transform 1 0 17070 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13034_
timestamp 0
transform -1 0 16790 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13035_
timestamp 0
transform 1 0 16790 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13036_
timestamp 0
transform 1 0 16930 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13037_
timestamp 0
transform 1 0 16750 0 1 250
box -6 -8 26 248
use FILL  FILL_1__13038_
timestamp 0
transform 1 0 16830 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13039_
timestamp 0
transform 1 0 16950 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13040_
timestamp 0
transform -1 0 16730 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13041_
timestamp 0
transform -1 0 16370 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13042_
timestamp 0
transform 1 0 15030 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13043_
timestamp 0
transform -1 0 16210 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13044_
timestamp 0
transform -1 0 12770 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13045_
timestamp 0
transform 1 0 16650 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13046_
timestamp 0
transform -1 0 16690 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13047_
timestamp 0
transform -1 0 15330 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13048_
timestamp 0
transform -1 0 15450 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13049_
timestamp 0
transform -1 0 15510 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13050_
timestamp 0
transform 1 0 16030 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13051_
timestamp 0
transform 1 0 16630 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13052_
timestamp 0
transform -1 0 16770 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13053_
timestamp 0
transform -1 0 16890 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13054_
timestamp 0
transform 1 0 16950 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13055_
timestamp 0
transform 1 0 16930 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13056_
timestamp 0
transform -1 0 16510 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13057_
timestamp 0
transform 1 0 17010 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__13058_
timestamp 0
transform 1 0 17010 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13059_
timestamp 0
transform 1 0 16930 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13060_
timestamp 0
transform -1 0 16870 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13061_
timestamp 0
transform 1 0 17030 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13062_
timestamp 0
transform -1 0 16590 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13063_
timestamp 0
transform 1 0 16730 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13064_
timestamp 0
transform 1 0 16450 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13065_
timestamp 0
transform 1 0 12610 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13066_
timestamp 0
transform 1 0 16790 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13067_
timestamp 0
transform -1 0 15370 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13068_
timestamp 0
transform 1 0 15270 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13069_
timestamp 0
transform -1 0 15710 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13070_
timestamp 0
transform -1 0 15850 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13071_
timestamp 0
transform 1 0 16390 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13072_
timestamp 0
transform 1 0 16510 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13073_
timestamp 0
transform 1 0 17050 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13074_
timestamp 0
transform 1 0 16510 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13075_
timestamp 0
transform -1 0 16910 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13076_
timestamp 0
transform -1 0 16930 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13077_
timestamp 0
transform -1 0 17050 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13078_
timestamp 0
transform -1 0 16790 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13079_
timestamp 0
transform -1 0 16630 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13080_
timestamp 0
transform -1 0 16910 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13081_
timestamp 0
transform -1 0 16750 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13082_
timestamp 0
transform -1 0 16710 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13083_
timestamp 0
transform -1 0 16590 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13084_
timestamp 0
transform 1 0 14450 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13085_
timestamp 0
transform -1 0 16310 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13086_
timestamp 0
transform -1 0 16170 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13087_
timestamp 0
transform 1 0 11810 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13088_
timestamp 0
transform -1 0 12270 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13089_
timestamp 0
transform 1 0 16410 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13090_
timestamp 0
transform 1 0 17030 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13091_
timestamp 0
transform -1 0 15570 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13092_
timestamp 0
transform -1 0 15430 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13093_
timestamp 0
transform 1 0 16310 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13094_
timestamp 0
transform 1 0 16250 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13095_
timestamp 0
transform -1 0 16490 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13096_
timestamp 0
transform 1 0 16990 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13097_
timestamp 0
transform -1 0 16850 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13098_
timestamp 0
transform 1 0 16670 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13099_
timestamp 0
transform 1 0 16750 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13100_
timestamp 0
transform 1 0 16610 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13101_
timestamp 0
transform -1 0 16590 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13102_
timestamp 0
transform -1 0 16070 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13103_
timestamp 0
transform 1 0 16710 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13104_
timestamp 0
transform 1 0 15930 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13105_
timestamp 0
transform 1 0 15790 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13106_
timestamp 0
transform -1 0 15670 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13107_
timestamp 0
transform -1 0 15530 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13108_
timestamp 0
transform 1 0 12590 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13109_
timestamp 0
transform 1 0 9530 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13110_
timestamp 0
transform 1 0 16570 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13111_
timestamp 0
transform 1 0 15550 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13112_
timestamp 0
transform -1 0 16110 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13113_
timestamp 0
transform 1 0 16230 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13114_
timestamp 0
transform -1 0 16250 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13115_
timestamp 0
transform -1 0 16390 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13116_
timestamp 0
transform 1 0 16370 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13117_
timestamp 0
transform 1 0 16210 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13118_
timestamp 0
transform -1 0 15990 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13119_
timestamp 0
transform 1 0 15950 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13120_
timestamp 0
transform -1 0 16110 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13121_
timestamp 0
transform 1 0 13630 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13122_
timestamp 0
transform 1 0 16830 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13123_
timestamp 0
transform 1 0 14910 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13124_
timestamp 0
transform -1 0 14310 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13125_
timestamp 0
transform -1 0 14030 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13126_
timestamp 0
transform 1 0 13750 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13127_
timestamp 0
transform -1 0 13070 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13128_
timestamp 0
transform -1 0 16450 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13129_
timestamp 0
transform -1 0 14630 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13130_
timestamp 0
transform -1 0 14790 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13131_
timestamp 0
transform -1 0 14150 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13132_
timestamp 0
transform -1 0 12950 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13133_
timestamp 0
transform -1 0 12130 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13134_
timestamp 0
transform 1 0 9770 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13135_
timestamp 0
transform 1 0 9630 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13136_
timestamp 0
transform 1 0 11290 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13137_
timestamp 0
transform -1 0 12430 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13138_
timestamp 0
transform 1 0 15970 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13139_
timestamp 0
transform -1 0 15710 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13140_
timestamp 0
transform 1 0 15650 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13141_
timestamp 0
transform 1 0 15530 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13142_
timestamp 0
transform -1 0 15630 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13143_
timestamp 0
transform 1 0 16090 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13144_
timestamp 0
transform -1 0 16310 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13145_
timestamp 0
transform 1 0 16170 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13146_
timestamp 0
transform -1 0 15370 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13147_
timestamp 0
transform -1 0 15770 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13148_
timestamp 0
transform -1 0 16050 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13149_
timestamp 0
transform 1 0 15890 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13150_
timestamp 0
transform 1 0 13870 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13151_
timestamp 0
transform -1 0 11870 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13152_
timestamp 0
transform 1 0 11990 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13153_
timestamp 0
transform -1 0 11750 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13154_
timestamp 0
transform -1 0 11610 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13155_
timestamp 0
transform 1 0 11410 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13156_
timestamp 0
transform 1 0 13370 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13157_
timestamp 0
transform -1 0 13530 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13158_
timestamp 0
transform -1 0 13230 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13159_
timestamp 0
transform -1 0 15110 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13160_
timestamp 0
transform -1 0 15830 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13161_
timestamp 0
transform -1 0 15870 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13162_
timestamp 0
transform -1 0 15710 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13163_
timestamp 0
transform -1 0 15110 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13164_
timestamp 0
transform 1 0 15190 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13165_
timestamp 0
transform -1 0 15470 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13166_
timestamp 0
transform 1 0 15330 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13167_
timestamp 0
transform -1 0 15210 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13168_
timestamp 0
transform -1 0 14970 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13169_
timestamp 0
transform -1 0 14990 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13170_
timestamp 0
transform -1 0 14830 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13171_
timestamp 0
transform -1 0 12530 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13172_
timestamp 0
transform -1 0 10950 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13173_
timestamp 0
transform 1 0 12650 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13174_
timestamp 0
transform -1 0 12270 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13175_
timestamp 0
transform 1 0 10770 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13176_
timestamp 0
transform -1 0 13310 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13177_
timestamp 0
transform 1 0 12790 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13178_
timestamp 0
transform -1 0 13850 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13179_
timestamp 0
transform -1 0 15250 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13180_
timestamp 0
transform 1 0 15430 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13181_
timestamp 0
transform 1 0 15650 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13182_
timestamp 0
transform 1 0 15530 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13183_
timestamp 0
transform -1 0 15310 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13184_
timestamp 0
transform -1 0 15030 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13185_
timestamp 0
transform 1 0 15170 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13186_
timestamp 0
transform 1 0 14810 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13187_
timestamp 0
transform -1 0 14470 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13188_
timestamp 0
transform -1 0 13810 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13189_
timestamp 0
transform 1 0 13930 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13190_
timestamp 0
transform -1 0 13670 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13191_
timestamp 0
transform -1 0 10170 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13192_
timestamp 0
transform -1 0 14590 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13193_
timestamp 0
transform -1 0 14550 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13194_
timestamp 0
transform 1 0 14690 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13195_
timestamp 0
transform -1 0 14690 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13196_
timestamp 0
transform 1 0 14370 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13197_
timestamp 0
transform -1 0 15730 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13198_
timestamp 0
transform -1 0 15610 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13199_
timestamp 0
transform -1 0 15410 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13200_
timestamp 0
transform -1 0 15110 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13201_
timestamp 0
transform 1 0 14870 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13202_
timestamp 0
transform -1 0 14750 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13203_
timestamp 0
transform -1 0 14590 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13204_
timestamp 0
transform -1 0 14830 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13205_
timestamp 0
transform 1 0 14950 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13206_
timestamp 0
transform -1 0 14690 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13207_
timestamp 0
transform 1 0 14330 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13208_
timestamp 0
transform -1 0 14110 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13209_
timestamp 0
transform 1 0 14250 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13210_
timestamp 0
transform -1 0 13970 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13211_
timestamp 0
transform 1 0 10270 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13212_
timestamp 0
transform -1 0 13030 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13213_
timestamp 0
transform -1 0 14250 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13214_
timestamp 0
transform -1 0 14110 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13215_
timestamp 0
transform -1 0 14450 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13216_
timestamp 0
transform 1 0 14310 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13217_
timestamp 0
transform -1 0 14170 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13218_
timestamp 0
transform -1 0 14050 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13219_
timestamp 0
transform -1 0 13710 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13220_
timestamp 0
transform -1 0 13550 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13221_
timestamp 0
transform -1 0 13410 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13222_
timestamp 0
transform -1 0 13350 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13223_
timestamp 0
transform -1 0 13270 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13224_
timestamp 0
transform -1 0 12750 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13225_
timestamp 0
transform 1 0 11590 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13226_
timestamp 0
transform -1 0 13230 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13227_
timestamp 0
transform -1 0 13070 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13228_
timestamp 0
transform 1 0 13330 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13229_
timestamp 0
transform -1 0 13650 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13230_
timestamp 0
transform -1 0 13210 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13231_
timestamp 0
transform -1 0 12910 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13232_
timestamp 0
transform -1 0 11630 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13233_
timestamp 0
transform 1 0 11190 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13234_
timestamp 0
transform -1 0 11470 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13235_
timestamp 0
transform -1 0 11350 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13236_
timestamp 0
transform -1 0 11410 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13237_
timestamp 0
transform -1 0 11290 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13238_
timestamp 0
transform -1 0 11170 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13239_
timestamp 0
transform 1 0 11530 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13240_
timestamp 0
transform -1 0 10990 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13241_
timestamp 0
transform 1 0 10950 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13242_
timestamp 0
transform -1 0 13790 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13243_
timestamp 0
transform 1 0 11750 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13244_
timestamp 0
transform -1 0 11930 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13245_
timestamp 0
transform -1 0 11290 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13246_
timestamp 0
transform -1 0 11130 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13247_
timestamp 0
transform 1 0 10530 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13248_
timestamp 0
transform -1 0 10430 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13249_
timestamp 0
transform -1 0 10310 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13250_
timestamp 0
transform 1 0 11230 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13251_
timestamp 0
transform -1 0 10170 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13252_
timestamp 0
transform -1 0 10070 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13253_
timestamp 0
transform -1 0 12090 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13254_
timestamp 0
transform 1 0 14490 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13255_
timestamp 0
transform -1 0 14350 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13256_
timestamp 0
transform 1 0 13410 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13257_
timestamp 0
transform 1 0 13490 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13258_
timestamp 0
transform -1 0 11170 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13259_
timestamp 0
transform 1 0 11290 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13260_
timestamp 0
transform -1 0 10890 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13261_
timestamp 0
transform -1 0 10770 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13262_
timestamp 0
transform -1 0 10590 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13263_
timestamp 0
transform 1 0 10650 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13264_
timestamp 0
transform -1 0 11050 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13265_
timestamp 0
transform -1 0 12030 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13266_
timestamp 0
transform 1 0 13850 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13267_
timestamp 0
transform -1 0 14010 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13268_
timestamp 0
transform 1 0 13710 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13269_
timestamp 0
transform -1 0 11890 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13270_
timestamp 0
transform 1 0 12030 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13271_
timestamp 0
transform -1 0 11790 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13272_
timestamp 0
transform 1 0 10990 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13273_
timestamp 0
transform -1 0 11250 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13274_
timestamp 0
transform 1 0 13430 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13275_
timestamp 0
transform -1 0 13930 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13276_
timestamp 0
transform 1 0 13910 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13277_
timestamp 0
transform -1 0 13770 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13278_
timestamp 0
transform -1 0 13650 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13279_
timestamp 0
transform -1 0 12390 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13280_
timestamp 0
transform 1 0 12530 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13281_
timestamp 0
transform 1 0 11750 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13282_
timestamp 0
transform -1 0 11490 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13283_
timestamp 0
transform 1 0 11110 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13284_
timestamp 0
transform -1 0 10730 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13285_
timestamp 0
transform 1 0 10590 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13286_
timestamp 0
transform 1 0 10930 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13287_
timestamp 0
transform -1 0 11390 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13288_
timestamp 0
transform 1 0 10850 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13289_
timestamp 0
transform 1 0 11590 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13290_
timestamp 0
transform -1 0 11150 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13291_
timestamp 0
transform 1 0 10970 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13292_
timestamp 0
transform -1 0 14630 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13293_
timestamp 0
transform 1 0 14410 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13294_
timestamp 0
transform 1 0 14290 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13295_
timestamp 0
transform -1 0 14210 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13296_
timestamp 0
transform -1 0 14170 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13297_
timestamp 0
transform 1 0 12430 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13298_
timestamp 0
transform -1 0 12290 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13299_
timestamp 0
transform 1 0 12170 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13300_
timestamp 0
transform -1 0 11390 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13301_
timestamp 0
transform -1 0 11250 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13302_
timestamp 0
transform -1 0 11450 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13303_
timestamp 0
transform -1 0 12150 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13304_
timestamp 0
transform 1 0 12550 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13305_
timestamp 0
transform -1 0 13210 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13306_
timestamp 0
transform -1 0 13070 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13307_
timestamp 0
transform -1 0 12950 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13308_
timestamp 0
transform 1 0 12790 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13309_
timestamp 0
transform 1 0 12830 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13310_
timestamp 0
transform 1 0 12650 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13311_
timestamp 0
transform 1 0 12710 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13312_
timestamp 0
transform 1 0 11990 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13313_
timestamp 0
transform -1 0 11850 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13314_
timestamp 0
transform 1 0 11670 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13315_
timestamp 0
transform 1 0 13070 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13316_
timestamp 0
transform -1 0 12770 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13317_
timestamp 0
transform -1 0 12610 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13318_
timestamp 0
transform 1 0 12210 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13319_
timestamp 0
transform -1 0 12470 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13320_
timestamp 0
transform -1 0 12330 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13321_
timestamp 0
transform 1 0 12290 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13322_
timestamp 0
transform 1 0 11890 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13323_
timestamp 0
transform 1 0 11630 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13324_
timestamp 0
transform 1 0 11470 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13325_
timestamp 0
transform 1 0 11530 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13326_
timestamp 0
transform 1 0 11690 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13327_
timestamp 0
transform -1 0 12090 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13328_
timestamp 0
transform 1 0 12230 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13329_
timestamp 0
transform 1 0 11930 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13330_
timestamp 0
transform -1 0 11730 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13331_
timestamp 0
transform 1 0 11790 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13332_
timestamp 0
transform 1 0 11610 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13333_
timestamp 0
transform 1 0 11850 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13334_
timestamp 0
transform 1 0 11990 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13335_
timestamp 0
transform -1 0 12010 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13336_
timestamp 0
transform 1 0 11830 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13337_
timestamp 0
transform 1 0 12970 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13338_
timestamp 0
transform -1 0 12870 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13339_
timestamp 0
transform 1 0 12950 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13340_
timestamp 0
transform -1 0 12850 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13341_
timestamp 0
transform -1 0 11630 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13342_
timestamp 0
transform -1 0 12170 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13343_
timestamp 0
transform -1 0 11790 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13344_
timestamp 0
transform 1 0 11950 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13345_
timestamp 0
transform 1 0 12210 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13346_
timestamp 0
transform 1 0 12070 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13347_
timestamp 0
transform -1 0 14710 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13348_
timestamp 0
transform 1 0 14930 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13349_
timestamp 0
transform -1 0 15090 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13350_
timestamp 0
transform -1 0 15190 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13351_
timestamp 0
transform 1 0 15010 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13352_
timestamp 0
transform 1 0 14730 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13353_
timestamp 0
transform 1 0 14870 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13354_
timestamp 0
transform -1 0 14990 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13355_
timestamp 0
transform -1 0 15130 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13356_
timestamp 0
transform 1 0 15030 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13357_
timestamp 0
transform 1 0 15170 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13358_
timestamp 0
transform -1 0 11650 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13359_
timestamp 0
transform -1 0 15310 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13360_
timestamp 0
transform 1 0 15130 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13361_
timestamp 0
transform -1 0 15270 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13362_
timestamp 0
transform 1 0 15110 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13363_
timestamp 0
transform 1 0 12330 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13364_
timestamp 0
transform 1 0 16570 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13365_
timestamp 0
transform -1 0 16830 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13366_
timestamp 0
transform 1 0 16810 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13367_
timestamp 0
transform 1 0 16770 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13368_
timestamp 0
transform 1 0 15250 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13369_
timestamp 0
transform 1 0 15110 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13370_
timestamp 0
transform 1 0 14810 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13371_
timestamp 0
transform -1 0 14990 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13372_
timestamp 0
transform -1 0 15670 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13373_
timestamp 0
transform -1 0 15810 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13374_
timestamp 0
transform -1 0 16070 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13375_
timestamp 0
transform 1 0 16190 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13376_
timestamp 0
transform 1 0 14110 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13377_
timestamp 0
transform -1 0 14250 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13378_
timestamp 0
transform -1 0 14670 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13379_
timestamp 0
transform -1 0 14790 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13380_
timestamp 0
transform 1 0 14050 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13381_
timestamp 0
transform 1 0 14930 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13382_
timestamp 0
transform 1 0 14770 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13383_
timestamp 0
transform 1 0 14250 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13384_
timestamp 0
transform 1 0 14310 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13385_
timestamp 0
transform 1 0 14390 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13386_
timestamp 0
transform -1 0 13830 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13387_
timestamp 0
transform -1 0 13870 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13388_
timestamp 0
transform -1 0 13970 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13389_
timestamp 0
transform -1 0 14250 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13390_
timestamp 0
transform 1 0 14170 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13391_
timestamp 0
transform 1 0 14290 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13392_
timestamp 0
transform -1 0 14630 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13393_
timestamp 0
transform 1 0 14470 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13394_
timestamp 0
transform -1 0 13530 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13395_
timestamp 0
transform -1 0 13690 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13396_
timestamp 0
transform 1 0 14530 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13397_
timestamp 0
transform 1 0 14350 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13398_
timestamp 0
transform 1 0 12990 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13399_
timestamp 0
transform -1 0 13150 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13400_
timestamp 0
transform -1 0 14850 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13401_
timestamp 0
transform -1 0 14970 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13402_
timestamp 0
transform -1 0 11950 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13403_
timestamp 0
transform -1 0 12070 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13404_
timestamp 0
transform 1 0 12970 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13405_
timestamp 0
transform -1 0 13110 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13406_
timestamp 0
transform -1 0 11950 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13407_
timestamp 0
transform -1 0 12710 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13408_
timestamp 0
transform 1 0 12530 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13409_
timestamp 0
transform -1 0 12570 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13410_
timestamp 0
transform -1 0 12750 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13411_
timestamp 0
transform 1 0 12590 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13412_
timestamp 0
transform -1 0 11670 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13413_
timestamp 0
transform -1 0 11790 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13414_
timestamp 0
transform 1 0 12430 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13415_
timestamp 0
transform -1 0 12290 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13416_
timestamp 0
transform 1 0 12590 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13417_
timestamp 0
transform 1 0 12430 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13418_
timestamp 0
transform 1 0 12930 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13419_
timestamp 0
transform -1 0 13070 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13420_
timestamp 0
transform -1 0 11650 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13421_
timestamp 0
transform -1 0 11810 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13422_
timestamp 0
transform -1 0 12210 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13423_
timestamp 0
transform -1 0 12370 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13424_
timestamp 0
transform -1 0 12470 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13425_
timestamp 0
transform -1 0 12590 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13426_
timestamp 0
transform 1 0 11070 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13427_
timestamp 0
transform -1 0 10810 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13502_
timestamp 0
transform -1 0 7650 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13503_
timestamp 0
transform -1 0 7510 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13504_
timestamp 0
transform -1 0 7790 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13505_
timestamp 0
transform 1 0 7950 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13506_
timestamp 0
transform 1 0 8350 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13507_
timestamp 0
transform 1 0 8590 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13508_
timestamp 0
transform 1 0 8430 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13509_
timestamp 0
transform -1 0 7750 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13510_
timestamp 0
transform -1 0 7150 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13511_
timestamp 0
transform 1 0 7190 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13512_
timestamp 0
transform -1 0 7070 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13513_
timestamp 0
transform 1 0 6370 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13514_
timestamp 0
transform 1 0 7410 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13515_
timestamp 0
transform -1 0 7670 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13516_
timestamp 0
transform 1 0 7810 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13517_
timestamp 0
transform -1 0 7150 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13518_
timestamp 0
transform 1 0 7930 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13519_
timestamp 0
transform 1 0 7550 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13520_
timestamp 0
transform 1 0 8070 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13521_
timestamp 0
transform -1 0 7830 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13522_
timestamp 0
transform 1 0 7810 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13523_
timestamp 0
transform 1 0 7530 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13524_
timestamp 0
transform -1 0 7690 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13525_
timestamp 0
transform -1 0 7670 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13526_
timestamp 0
transform -1 0 6990 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13527_
timestamp 0
transform 1 0 7570 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__13528_
timestamp 0
transform -1 0 10110 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13529_
timestamp 0
transform 1 0 9050 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13530_
timestamp 0
transform -1 0 8910 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13531_
timestamp 0
transform -1 0 9490 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13532_
timestamp 0
transform -1 0 8730 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13533_
timestamp 0
transform 1 0 8690 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13534_
timestamp 0
transform -1 0 8750 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13535_
timestamp 0
transform -1 0 7890 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13536_
timestamp 0
transform 1 0 8230 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13537_
timestamp 0
transform 1 0 8670 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13538_
timestamp 0
transform 1 0 8910 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13539_
timestamp 0
transform -1 0 9210 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13540_
timestamp 0
transform -1 0 8570 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13541_
timestamp 0
transform -1 0 8850 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__13542_
timestamp 0
transform 1 0 8270 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13543_
timestamp 0
transform -1 0 8310 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13544_
timestamp 0
transform -1 0 7150 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13545_
timestamp 0
transform 1 0 6710 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13546_
timestamp 0
transform -1 0 7890 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13547_
timestamp 0
transform -1 0 7570 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13548_
timestamp 0
transform 1 0 10250 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13549_
timestamp 0
transform -1 0 9890 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13550_
timestamp 0
transform -1 0 10010 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13551_
timestamp 0
transform 1 0 10210 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13552_
timestamp 0
transform -1 0 9750 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13553_
timestamp 0
transform -1 0 10030 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13554_
timestamp 0
transform 1 0 9850 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13555_
timestamp 0
transform -1 0 7770 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13556_
timestamp 0
transform -1 0 8170 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13557_
timestamp 0
transform 1 0 7850 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13558_
timestamp 0
transform 1 0 8130 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13559_
timestamp 0
transform -1 0 8470 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13560_
timestamp 0
transform 1 0 8290 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13561_
timestamp 0
transform 1 0 7990 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13562_
timestamp 0
transform -1 0 7610 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13563_
timestamp 0
transform 1 0 7110 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13564_
timestamp 0
transform -1 0 6610 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13565_
timestamp 0
transform 1 0 7290 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13566_
timestamp 0
transform -1 0 8870 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13567_
timestamp 0
transform 1 0 9390 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13568_
timestamp 0
transform 1 0 9910 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13569_
timestamp 0
transform 1 0 7410 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13570_
timestamp 0
transform 1 0 7250 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13571_
timestamp 0
transform -1 0 8190 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13572_
timestamp 0
transform -1 0 6210 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13573_
timestamp 0
transform 1 0 8450 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13574_
timestamp 0
transform -1 0 9270 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13575_
timestamp 0
transform -1 0 9450 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13576_
timestamp 0
transform -1 0 8590 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13577_
timestamp 0
transform -1 0 7430 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13578_
timestamp 0
transform -1 0 7730 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13579_
timestamp 0
transform 1 0 7830 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13580_
timestamp 0
transform 1 0 8130 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13581_
timestamp 0
transform -1 0 8470 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13582_
timestamp 0
transform 1 0 8290 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13583_
timestamp 0
transform 1 0 7970 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13584_
timestamp 0
transform -1 0 7070 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13585_
timestamp 0
transform 1 0 10330 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13586_
timestamp 0
transform -1 0 9670 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13587_
timestamp 0
transform -1 0 9390 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13588_
timestamp 0
transform -1 0 9530 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13589_
timestamp 0
transform -1 0 9630 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13590_
timestamp 0
transform -1 0 9330 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13591_
timestamp 0
transform 1 0 9250 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13592_
timestamp 0
transform -1 0 8970 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13593_
timestamp 0
transform -1 0 8370 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13594_
timestamp 0
transform 1 0 9310 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13595_
timestamp 0
transform 1 0 9170 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13596_
timestamp 0
transform 1 0 8890 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13597_
timestamp 0
transform 1 0 8610 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13598_
timestamp 0
transform -1 0 8350 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13599_
timestamp 0
transform 1 0 7730 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13600_
timestamp 0
transform -1 0 7150 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13601_
timestamp 0
transform 1 0 6290 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13602_
timestamp 0
transform 1 0 9210 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13603_
timestamp 0
transform -1 0 9310 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13604_
timestamp 0
transform 1 0 9050 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13605_
timestamp 0
transform 1 0 9150 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13606_
timestamp 0
transform 1 0 8810 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13607_
timestamp 0
transform -1 0 9010 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13608_
timestamp 0
transform -1 0 7430 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13609_
timestamp 0
transform 1 0 6810 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13610_
timestamp 0
transform -1 0 6410 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13611_
timestamp 0
transform -1 0 6150 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13612_
timestamp 0
transform 1 0 6530 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13613_
timestamp 0
transform 1 0 6230 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13614_
timestamp 0
transform -1 0 6590 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13615_
timestamp 0
transform 1 0 6290 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13616_
timestamp 0
transform -1 0 6470 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13617_
timestamp 0
transform -1 0 6350 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13618_
timestamp 0
transform 1 0 9110 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__13619_
timestamp 0
transform 1 0 9390 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__13620_
timestamp 0
transform 1 0 9230 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__13621_
timestamp 0
transform 1 0 7010 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13622_
timestamp 0
transform -1 0 6090 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13623_
timestamp 0
transform -1 0 9290 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13624_
timestamp 0
transform 1 0 9230 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13625_
timestamp 0
transform -1 0 8410 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13626_
timestamp 0
transform -1 0 8110 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13627_
timestamp 0
transform 1 0 8210 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13628_
timestamp 0
transform -1 0 7970 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13629_
timestamp 0
transform -1 0 6690 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13630_
timestamp 0
transform -1 0 5550 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13631_
timestamp 0
transform -1 0 6050 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13632_
timestamp 0
transform -1 0 6150 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13633_
timestamp 0
transform -1 0 5930 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13634_
timestamp 0
transform -1 0 5250 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13635_
timestamp 0
transform -1 0 5410 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13636_
timestamp 0
transform -1 0 4770 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13637_
timestamp 0
transform -1 0 4610 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13638_
timestamp 0
transform -1 0 5290 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13639_
timestamp 0
transform 1 0 5390 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13640_
timestamp 0
transform 1 0 4850 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13641_
timestamp 0
transform 1 0 5510 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13642_
timestamp 0
transform 1 0 6750 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13643_
timestamp 0
transform 1 0 6570 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13644_
timestamp 0
transform 1 0 6710 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13645_
timestamp 0
transform 1 0 6870 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13646_
timestamp 0
transform -1 0 6670 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13647_
timestamp 0
transform -1 0 5110 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13648_
timestamp 0
transform -1 0 5010 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13649_
timestamp 0
transform -1 0 5810 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13650_
timestamp 0
transform 1 0 6810 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13651_
timestamp 0
transform 1 0 9890 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13652_
timestamp 0
transform 1 0 10110 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13653_
timestamp 0
transform 1 0 9950 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13654_
timestamp 0
transform 1 0 8990 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13655_
timestamp 0
transform 1 0 8850 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13656_
timestamp 0
transform 1 0 7290 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13657_
timestamp 0
transform 1 0 6330 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13658_
timestamp 0
transform -1 0 7570 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13659_
timestamp 0
transform 1 0 7650 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13660_
timestamp 0
transform -1 0 6010 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13661_
timestamp 0
transform -1 0 5890 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13662_
timestamp 0
transform 1 0 6050 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13663_
timestamp 0
transform -1 0 5730 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13664_
timestamp 0
transform -1 0 5650 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13665_
timestamp 0
transform 1 0 5770 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13666_
timestamp 0
transform -1 0 4390 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13667_
timestamp 0
transform -1 0 4490 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13668_
timestamp 0
transform 1 0 4970 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13669_
timestamp 0
transform 1 0 5130 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13670_
timestamp 0
transform -1 0 5610 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13671_
timestamp 0
transform 1 0 5650 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13672_
timestamp 0
transform -1 0 5610 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13673_
timestamp 0
transform 1 0 10250 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13674_
timestamp 0
transform 1 0 9950 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13675_
timestamp 0
transform 1 0 9790 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13676_
timestamp 0
transform 1 0 9290 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13677_
timestamp 0
transform 1 0 9130 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13678_
timestamp 0
transform 1 0 7830 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13679_
timestamp 0
transform -1 0 7710 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13680_
timestamp 0
transform -1 0 7070 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13681_
timestamp 0
transform 1 0 6270 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13682_
timestamp 0
transform -1 0 5970 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13683_
timestamp 0
transform -1 0 6570 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13684_
timestamp 0
transform -1 0 6410 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13685_
timestamp 0
transform -1 0 6130 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13686_
timestamp 0
transform 1 0 6150 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13687_
timestamp 0
transform -1 0 6010 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13688_
timestamp 0
transform -1 0 5870 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13689_
timestamp 0
transform 1 0 6030 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13690_
timestamp 0
transform -1 0 6090 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13691_
timestamp 0
transform 1 0 5930 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13692_
timestamp 0
transform -1 0 5970 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13693_
timestamp 0
transform -1 0 6230 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13694_
timestamp 0
transform -1 0 6990 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13695_
timestamp 0
transform 1 0 6150 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13696_
timestamp 0
transform 1 0 9650 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13697_
timestamp 0
transform -1 0 9430 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13698_
timestamp 0
transform -1 0 8730 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13699_
timestamp 0
transform 1 0 7470 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13700_
timestamp 0
transform -1 0 7350 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13701_
timestamp 0
transform 1 0 6270 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13702_
timestamp 0
transform -1 0 6850 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13703_
timestamp 0
transform 1 0 6590 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13704_
timestamp 0
transform -1 0 6750 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13705_
timestamp 0
transform 1 0 6470 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13706_
timestamp 0
transform -1 0 6450 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13707_
timestamp 0
transform -1 0 5770 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13708_
timestamp 0
transform 1 0 6850 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13709_
timestamp 0
transform 1 0 6290 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13710_
timestamp 0
transform 1 0 6430 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13711_
timestamp 0
transform 1 0 6490 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13712_
timestamp 0
transform -1 0 7310 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__13713_
timestamp 0
transform -1 0 5790 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13714_
timestamp 0
transform 1 0 7670 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13715_
timestamp 0
transform 1 0 6670 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13716_
timestamp 0
transform -1 0 9010 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13717_
timestamp 0
transform 1 0 8330 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13718_
timestamp 0
transform 1 0 8170 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13719_
timestamp 0
transform -1 0 6670 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13720_
timestamp 0
transform 1 0 7410 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13721_
timestamp 0
transform -1 0 6150 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13722_
timestamp 0
transform -1 0 6630 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13723_
timestamp 0
transform -1 0 6370 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13724_
timestamp 0
transform -1 0 7150 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13725_
timestamp 0
transform 1 0 7010 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13726_
timestamp 0
transform -1 0 7010 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13727_
timestamp 0
transform -1 0 6210 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13728_
timestamp 0
transform 1 0 6250 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13729_
timestamp 0
transform -1 0 5870 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13730_
timestamp 0
transform 1 0 6570 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13731_
timestamp 0
transform -1 0 6750 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13732_
timestamp 0
transform -1 0 6050 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13733_
timestamp 0
transform -1 0 6070 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13734_
timestamp 0
transform 1 0 5890 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13735_
timestamp 0
transform -1 0 6850 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13736_
timestamp 0
transform -1 0 6530 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13737_
timestamp 0
transform 1 0 6170 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13738_
timestamp 0
transform 1 0 6330 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13739_
timestamp 0
transform -1 0 5990 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13740_
timestamp 0
transform 1 0 6430 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13741_
timestamp 0
transform 1 0 6450 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13742_
timestamp 0
transform -1 0 7350 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13743_
timestamp 0
transform 1 0 6870 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13744_
timestamp 0
transform -1 0 9690 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13745_
timestamp 0
transform 1 0 9650 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13746_
timestamp 0
transform -1 0 9550 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13747_
timestamp 0
transform 1 0 8710 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13748_
timestamp 0
transform 1 0 7270 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13749_
timestamp 0
transform -1 0 7090 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13750_
timestamp 0
transform 1 0 6790 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13751_
timestamp 0
transform -1 0 6950 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13752_
timestamp 0
transform -1 0 7210 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13753_
timestamp 0
transform 1 0 7170 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13754_
timestamp 0
transform -1 0 6910 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13755_
timestamp 0
transform -1 0 7050 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13756_
timestamp 0
transform -1 0 6750 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13757_
timestamp 0
transform 1 0 7030 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13758_
timestamp 0
transform -1 0 6910 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13759_
timestamp 0
transform 1 0 6450 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13760_
timestamp 0
transform 1 0 6590 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13761_
timestamp 0
transform -1 0 6890 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13762_
timestamp 0
transform -1 0 6890 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13763_
timestamp 0
transform 1 0 6730 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13764_
timestamp 0
transform -1 0 6710 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13765_
timestamp 0
transform -1 0 6950 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13766_
timestamp 0
transform 1 0 6610 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13767_
timestamp 0
transform 1 0 6330 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13768_
timestamp 0
transform 1 0 6450 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13769_
timestamp 0
transform -1 0 8110 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13770_
timestamp 0
transform 1 0 7890 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13771_
timestamp 0
transform 1 0 8570 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13772_
timestamp 0
transform -1 0 8370 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13773_
timestamp 0
transform -1 0 8070 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13774_
timestamp 0
transform 1 0 8330 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13775_
timestamp 0
transform -1 0 8050 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13776_
timestamp 0
transform -1 0 7970 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13777_
timestamp 0
transform -1 0 8210 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13778_
timestamp 0
transform 1 0 8190 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13779_
timestamp 0
transform -1 0 7790 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13780_
timestamp 0
transform 1 0 7510 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13781_
timestamp 0
transform -1 0 7290 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13782_
timestamp 0
transform -1 0 7130 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13783_
timestamp 0
transform -1 0 6990 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13784_
timestamp 0
transform -1 0 6890 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13785_
timestamp 0
transform 1 0 6770 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13786_
timestamp 0
transform -1 0 6650 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13787_
timestamp 0
transform 1 0 6290 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13788_
timestamp 0
transform -1 0 6610 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13789_
timestamp 0
transform 1 0 6470 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13790_
timestamp 0
transform -1 0 7690 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13791_
timestamp 0
transform -1 0 7390 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13792_
timestamp 0
transform -1 0 8970 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13793_
timestamp 0
transform 1 0 8190 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13794_
timestamp 0
transform -1 0 8550 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13795_
timestamp 0
transform 1 0 8570 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13796_
timestamp 0
transform -1 0 8390 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13797_
timestamp 0
transform 1 0 8630 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13798_
timestamp 0
transform 1 0 8490 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13799_
timestamp 0
transform -1 0 8090 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13800_
timestamp 0
transform 1 0 8650 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13801_
timestamp 0
transform -1 0 8750 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13802_
timestamp 0
transform -1 0 8830 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13803_
timestamp 0
transform -1 0 7810 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13804_
timestamp 0
transform -1 0 7310 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13805_
timestamp 0
transform 1 0 7450 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13806_
timestamp 0
transform -1 0 7310 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13807_
timestamp 0
transform -1 0 7430 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__13808_
timestamp 0
transform -1 0 9810 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13809_
timestamp 0
transform -1 0 8870 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13810_
timestamp 0
transform 1 0 9010 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13811_
timestamp 0
transform 1 0 9110 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13812_
timestamp 0
transform 1 0 9070 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13813_
timestamp 0
transform 1 0 9210 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13814_
timestamp 0
transform -1 0 8910 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13815_
timestamp 0
transform -1 0 8930 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13816_
timestamp 0
transform -1 0 8810 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13817_
timestamp 0
transform 1 0 9230 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13818_
timestamp 0
transform 1 0 9350 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13819_
timestamp 0
transform -1 0 9350 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13820_
timestamp 0
transform 1 0 9070 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13821_
timestamp 0
transform 1 0 8530 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13822_
timestamp 0
transform -1 0 8250 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13823_
timestamp 0
transform 1 0 7910 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13824_
timestamp 0
transform 1 0 7650 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13825_
timestamp 0
transform 1 0 8230 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13826_
timestamp 0
transform -1 0 8410 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13827_
timestamp 0
transform 1 0 7930 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13828_
timestamp 0
transform 1 0 8090 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13829_
timestamp 0
transform -1 0 8050 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13830_
timestamp 0
transform -1 0 7630 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13831_
timestamp 0
transform 1 0 7090 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13832_
timestamp 0
transform -1 0 7350 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13833_
timestamp 0
transform -1 0 8350 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13834_
timestamp 0
transform -1 0 10110 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13835_
timestamp 0
transform 1 0 10430 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13836_
timestamp 0
transform 1 0 10030 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13837_
timestamp 0
transform -1 0 9970 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__13838_
timestamp 0
transform 1 0 9770 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13839_
timestamp 0
transform -1 0 9470 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13840_
timestamp 0
transform -1 0 9470 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13841_
timestamp 0
transform 1 0 9330 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13842_
timestamp 0
transform -1 0 8010 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13843_
timestamp 0
transform -1 0 7790 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13844_
timestamp 0
transform 1 0 8170 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13845_
timestamp 0
transform -1 0 7910 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13846_
timestamp 0
transform -1 0 7470 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__13847_
timestamp 0
transform 1 0 7470 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13848_
timestamp 0
transform -1 0 8450 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__13849_
timestamp 0
transform -1 0 5810 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13850_
timestamp 0
transform -1 0 5690 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13851_
timestamp 0
transform -1 0 5930 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13852_
timestamp 0
transform -1 0 6090 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13853_
timestamp 0
transform -1 0 6730 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13854_
timestamp 0
transform 1 0 6990 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13855_
timestamp 0
transform 1 0 6830 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13856_
timestamp 0
transform -1 0 6730 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13857_
timestamp 0
transform -1 0 7790 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13858_
timestamp 0
transform -1 0 7910 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13859_
timestamp 0
transform 1 0 6710 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13860_
timestamp 0
transform 1 0 6670 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13861_
timestamp 0
transform -1 0 7930 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13862_
timestamp 0
transform 1 0 7970 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13863_
timestamp 0
transform 1 0 7810 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13864_
timestamp 0
transform -1 0 8030 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13865_
timestamp 0
transform -1 0 7430 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13866_
timestamp 0
transform 1 0 7910 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13867_
timestamp 0
transform 1 0 7530 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13868_
timestamp 0
transform 1 0 7650 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13869_
timestamp 0
transform 1 0 8590 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13870_
timestamp 0
transform 1 0 8650 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__13871_
timestamp 0
transform -1 0 8170 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13872_
timestamp 0
transform -1 0 8250 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13873_
timestamp 0
transform 1 0 5490 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13874_
timestamp 0
transform -1 0 5950 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13875_
timestamp 0
transform -1 0 6270 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13876_
timestamp 0
transform -1 0 6410 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13877_
timestamp 0
transform -1 0 6550 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13878_
timestamp 0
transform -1 0 7170 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13879_
timestamp 0
transform 1 0 7770 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13880_
timestamp 0
transform 1 0 7610 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13881_
timestamp 0
transform -1 0 7110 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13882_
timestamp 0
transform 1 0 7530 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13883_
timestamp 0
transform 1 0 7290 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13884_
timestamp 0
transform -1 0 6890 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13885_
timestamp 0
transform -1 0 7010 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13886_
timestamp 0
transform -1 0 7290 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13887_
timestamp 0
transform -1 0 8110 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13888_
timestamp 0
transform -1 0 7390 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13889_
timestamp 0
transform 1 0 7190 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13890_
timestamp 0
transform -1 0 8210 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13891_
timestamp 0
transform 1 0 8470 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13892_
timestamp 0
transform 1 0 8770 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13893_
timestamp 0
transform 1 0 8330 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13894_
timestamp 0
transform -1 0 8630 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13895_
timestamp 0
transform 1 0 8210 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13896_
timestamp 0
transform -1 0 8070 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13897_
timestamp 0
transform -1 0 7930 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13898_
timestamp 0
transform 1 0 8010 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13899_
timestamp 0
transform -1 0 7510 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13900_
timestamp 0
transform 1 0 8470 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13901_
timestamp 0
transform 1 0 8410 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13902_
timestamp 0
transform 1 0 9550 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13903_
timestamp 0
transform 1 0 9510 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13904_
timestamp 0
transform -1 0 8790 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13905_
timestamp 0
transform -1 0 9130 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13906_
timestamp 0
transform -1 0 6210 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13907_
timestamp 0
transform -1 0 6610 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13908_
timestamp 0
transform 1 0 6450 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13909_
timestamp 0
transform -1 0 7250 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13910_
timestamp 0
transform 1 0 8550 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13911_
timestamp 0
transform 1 0 8650 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13912_
timestamp 0
transform 1 0 8050 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13913_
timestamp 0
transform 1 0 8890 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13914_
timestamp 0
transform 1 0 9030 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13915_
timestamp 0
transform 1 0 8850 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13916_
timestamp 0
transform -1 0 8890 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13917_
timestamp 0
transform 1 0 8730 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13918_
timestamp 0
transform -1 0 8470 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13919_
timestamp 0
transform -1 0 8630 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13920_
timestamp 0
transform 1 0 8730 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13921_
timestamp 0
transform -1 0 7650 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__13922_
timestamp 0
transform 1 0 8730 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13923_
timestamp 0
transform -1 0 7130 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13924_
timestamp 0
transform -1 0 9530 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13925_
timestamp 0
transform -1 0 9650 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__13926_
timestamp 0
transform 1 0 10030 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13927_
timestamp 0
transform 1 0 9410 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13928_
timestamp 0
transform 1 0 7650 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13929_
timestamp 0
transform 1 0 7530 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13930_
timestamp 0
transform 1 0 7770 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13931_
timestamp 0
transform 1 0 9470 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13932_
timestamp 0
transform 1 0 8810 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13933_
timestamp 0
transform -1 0 8990 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13934_
timestamp 0
transform -1 0 9070 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13935_
timestamp 0
transform -1 0 7910 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13936_
timestamp 0
transform -1 0 7510 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13937_
timestamp 0
transform -1 0 7750 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13938_
timestamp 0
transform -1 0 7390 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13939_
timestamp 0
transform -1 0 6730 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13940_
timestamp 0
transform -1 0 7010 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13941_
timestamp 0
transform -1 0 6890 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13942_
timestamp 0
transform -1 0 8130 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13943_
timestamp 0
transform 1 0 7590 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13944_
timestamp 0
transform 1 0 10290 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13945_
timestamp 0
transform 1 0 10150 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__13946_
timestamp 0
transform -1 0 10330 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13947_
timestamp 0
transform 1 0 10430 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13948_
timestamp 0
transform 1 0 10590 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__13949_
timestamp 0
transform 1 0 10490 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13950_
timestamp 0
transform 1 0 10210 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13951_
timestamp 0
transform 1 0 8250 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13952_
timestamp 0
transform 1 0 9510 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13953_
timestamp 0
transform 1 0 9970 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13954_
timestamp 0
transform 1 0 9370 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13955_
timestamp 0
transform -1 0 10290 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13956_
timestamp 0
transform -1 0 10130 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13957_
timestamp 0
transform 1 0 10730 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13958_
timestamp 0
transform 1 0 10410 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13959_
timestamp 0
transform 1 0 10590 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13960_
timestamp 0
transform 1 0 9770 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13961_
timestamp 0
transform -1 0 8070 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13962_
timestamp 0
transform 1 0 9250 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13963_
timestamp 0
transform -1 0 9130 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13964_
timestamp 0
transform -1 0 9370 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13965_
timestamp 0
transform 1 0 9090 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13966_
timestamp 0
transform 1 0 9610 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13967_
timestamp 0
transform -1 0 9190 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13968_
timestamp 0
transform 1 0 10210 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13969_
timestamp 0
transform 1 0 10070 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13970_
timestamp 0
transform -1 0 9130 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13971_
timestamp 0
transform 1 0 9830 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13972_
timestamp 0
transform -1 0 8830 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13973_
timestamp 0
transform -1 0 8550 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13974_
timestamp 0
transform 1 0 9350 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13975_
timestamp 0
transform 1 0 9190 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13976_
timestamp 0
transform -1 0 9670 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13977_
timestamp 0
transform -1 0 8710 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13978_
timestamp 0
transform -1 0 8230 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13979_
timestamp 0
transform -1 0 9910 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__13980_
timestamp 0
transform 1 0 8370 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1__13981_
timestamp 0
transform 1 0 9850 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13982_
timestamp 0
transform -1 0 9610 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__13983_
timestamp 0
transform 1 0 9690 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13984_
timestamp 0
transform -1 0 9570 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13985_
timestamp 0
transform 1 0 9190 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__13986_
timestamp 0
transform 1 0 9510 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__13987_
timestamp 0
transform 1 0 10310 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__13988_
timestamp 0
transform 1 0 10350 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13989_
timestamp 0
transform 1 0 10490 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__13990_
timestamp 0
transform 1 0 10370 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__13991_
timestamp 0
transform -1 0 10770 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13992_
timestamp 0
transform 1 0 9970 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1__13993_
timestamp 0
transform 1 0 10890 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13994_
timestamp 0
transform 1 0 10670 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__13995_
timestamp 0
transform 1 0 10630 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13996_
timestamp 0
transform 1 0 10350 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13997_
timestamp 0
transform -1 0 10490 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__13998_
timestamp 0
transform -1 0 10150 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__13999_
timestamp 0
transform -1 0 10450 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__14000_
timestamp 0
transform -1 0 9970 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__14001_
timestamp 0
transform 1 0 9790 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__14002_
timestamp 0
transform -1 0 9750 0 1 16090
box -6 -8 26 248
use FILL  FILL_1__14003_
timestamp 0
transform -1 0 9770 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__14004_
timestamp 0
transform -1 0 10270 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__14005_
timestamp 0
transform -1 0 10310 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__14006_
timestamp 0
transform -1 0 10150 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__14007_
timestamp 0
transform -1 0 10090 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__14008_
timestamp 0
transform 1 0 9990 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1__14009_
timestamp 0
transform -1 0 9950 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__14010_
timestamp 0
transform -1 0 9590 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__14011_
timestamp 0
transform -1 0 9650 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__14012_
timestamp 0
transform 1 0 9610 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__14013_
timestamp 0
transform -1 0 8670 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__14014_
timestamp 0
transform -1 0 9850 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__14015_
timestamp 0
transform -1 0 10530 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__14016_
timestamp 0
transform 1 0 10710 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__14017_
timestamp 0
transform -1 0 10650 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__14018_
timestamp 0
transform 1 0 10850 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__14019_
timestamp 0
transform -1 0 10710 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__14020_
timestamp 0
transform -1 0 10810 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__14021_
timestamp 0
transform 1 0 10990 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__14022_
timestamp 0
transform 1 0 11110 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__14023_
timestamp 0
transform -1 0 10550 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__14024_
timestamp 0
transform -1 0 10990 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__14025_
timestamp 0
transform 1 0 11230 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__14026_
timestamp 0
transform -1 0 10850 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__14027_
timestamp 0
transform 1 0 10410 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__14028_
timestamp 0
transform -1 0 9430 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__14029_
timestamp 0
transform -1 0 9730 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__14030_
timestamp 0
transform 1 0 10190 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__14031_
timestamp 0
transform -1 0 9790 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__14032_
timestamp 0
transform 1 0 8910 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__14033_
timestamp 0
transform 1 0 10230 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__14034_
timestamp 0
transform -1 0 10030 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__14035_
timestamp 0
transform 1 0 10070 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__14036_
timestamp 0
transform 1 0 10490 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__14037_
timestamp 0
transform -1 0 10650 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__14038_
timestamp 0
transform -1 0 10610 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__14039_
timestamp 0
transform 1 0 10610 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__14040_
timestamp 0
transform -1 0 10850 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__14041_
timestamp 0
transform 1 0 10850 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__14042_
timestamp 0
transform 1 0 11010 0 1 14650
box -6 -8 26 248
use FILL  FILL_1__14043_
timestamp 0
transform 1 0 10930 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__14044_
timestamp 0
transform -1 0 10890 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__14045_
timestamp 0
transform -1 0 10610 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__14046_
timestamp 0
transform 1 0 10730 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__14047_
timestamp 0
transform -1 0 10450 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__14048_
timestamp 0
transform -1 0 9950 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__14049_
timestamp 0
transform 1 0 9970 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__14050_
timestamp 0
transform -1 0 9770 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__14051_
timestamp 0
transform -1 0 9530 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__14052_
timestamp 0
transform -1 0 9830 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__14053_
timestamp 0
transform -1 0 9650 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__14054_
timestamp 0
transform 1 0 9670 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__14055_
timestamp 0
transform -1 0 9830 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__14056_
timestamp 0
transform 1 0 10450 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__14057_
timestamp 0
transform -1 0 9830 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__14058_
timestamp 0
transform 1 0 10730 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__14059_
timestamp 0
transform -1 0 9930 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__14060_
timestamp 0
transform -1 0 10450 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__14061_
timestamp 0
transform 1 0 10270 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__14062_
timestamp 0
transform 1 0 10150 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__14063_
timestamp 0
transform 1 0 10010 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1__14064_
timestamp 0
transform -1 0 10730 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__14065_
timestamp 0
transform 1 0 10450 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__14066_
timestamp 0
transform -1 0 10310 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__14067_
timestamp 0
transform -1 0 10170 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__14068_
timestamp 0
transform 1 0 9350 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__14069_
timestamp 0
transform 1 0 10830 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__14070_
timestamp 0
transform -1 0 10610 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__14071_
timestamp 0
transform -1 0 10090 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__14072_
timestamp 0
transform -1 0 10210 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__14073_
timestamp 0
transform 1 0 10550 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__14074_
timestamp 0
transform 1 0 10450 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__14075_
timestamp 0
transform 1 0 10470 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__14076_
timestamp 0
transform -1 0 10610 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__14077_
timestamp 0
transform -1 0 10370 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__14078_
timestamp 0
transform 1 0 10110 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__14079_
timestamp 0
transform -1 0 9110 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__14080_
timestamp 0
transform -1 0 9670 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__14081_
timestamp 0
transform 1 0 9370 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__14082_
timestamp 0
transform -1 0 9250 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__14083_
timestamp 0
transform 1 0 9510 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__14084_
timestamp 0
transform 1 0 10430 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__14085_
timestamp 0
transform -1 0 10070 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__14086_
timestamp 0
transform 1 0 10210 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__14087_
timestamp 0
transform -1 0 9930 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__14088_
timestamp 0
transform 1 0 9470 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__14089_
timestamp 0
transform 1 0 9270 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__14090_
timestamp 0
transform 1 0 11070 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__14091_
timestamp 0
transform 1 0 10930 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1__14092_
timestamp 0
transform 1 0 10050 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__14093_
timestamp 0
transform 1 0 9990 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__14094_
timestamp 0
transform -1 0 9910 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__14095_
timestamp 0
transform 1 0 9870 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__14096_
timestamp 0
transform -1 0 9790 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__14097_
timestamp 0
transform -1 0 9770 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__14098_
timestamp 0
transform -1 0 9650 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__14099_
timestamp 0
transform 1 0 8770 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__14100_
timestamp 0
transform 1 0 8430 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__14101_
timestamp 0
transform 1 0 8770 0 1 12730
box -6 -8 26 248
use FILL  FILL_1__14102_
timestamp 0
transform -1 0 10350 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__14103_
timestamp 0
transform 1 0 10310 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__14104_
timestamp 0
transform -1 0 9690 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__14105_
timestamp 0
transform -1 0 9830 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__14106_
timestamp 0
transform -1 0 9570 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__14107_
timestamp 0
transform -1 0 9510 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__14108_
timestamp 0
transform 1 0 9590 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__14109_
timestamp 0
transform 1 0 9730 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__14110_
timestamp 0
transform -1 0 9870 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__14111_
timestamp 0
transform 1 0 9330 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__14112_
timestamp 0
transform 1 0 9190 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__14113_
timestamp 0
transform 1 0 7590 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__14114_
timestamp 0
transform 1 0 9430 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__14115_
timestamp 0
transform 1 0 9290 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__14116_
timestamp 0
transform -1 0 9590 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__14117_
timestamp 0
transform 1 0 9710 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1__14118_
timestamp 0
transform -1 0 7870 0 1 12250
box -6 -8 26 248
use FILL  FILL_1__14119_
timestamp 0
transform -1 0 10150 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__14120_
timestamp 0
transform -1 0 10190 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__14121_
timestamp 0
transform 1 0 9850 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__14122_
timestamp 0
transform 1 0 9710 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__14123_
timestamp 0
transform -1 0 8430 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__14124_
timestamp 0
transform -1 0 8570 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__14125_
timestamp 0
transform 1 0 8110 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__14126_
timestamp 0
transform -1 0 8530 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__14127_
timestamp 0
transform 1 0 8650 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__14128_
timestamp 0
transform -1 0 8510 0 1 15130
box -6 -8 26 248
use FILL  FILL_1__14129_
timestamp 0
transform 1 0 9170 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__14130_
timestamp 0
transform 1 0 9010 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__14131_
timestamp 0
transform -1 0 10230 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__14132_
timestamp 0
transform 1 0 10150 0 1 13690
box -6 -8 26 248
use FILL  FILL_1__14133_
timestamp 0
transform -1 0 10950 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__14134_
timestamp 0
transform 1 0 10790 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__14135_
timestamp 0
transform -1 0 8450 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__14136_
timestamp 0
transform -1 0 9210 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__14137_
timestamp 0
transform 1 0 9030 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__14138_
timestamp 0
transform 1 0 7930 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__14139_
timestamp 0
transform -1 0 9070 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__14140_
timestamp 0
transform 1 0 8890 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1__14141_
timestamp 0
transform 1 0 7690 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__14142_
timestamp 0
transform 1 0 7630 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__14143_
timestamp 0
transform 1 0 7810 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__14144_
timestamp 0
transform -1 0 7810 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__14145_
timestamp 0
transform -1 0 6570 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__14146_
timestamp 0
transform 1 0 6410 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__14147_
timestamp 0
transform 1 0 7550 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__14148_
timestamp 0
transform 1 0 7150 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__14149_
timestamp 0
transform -1 0 7470 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1__14150_
timestamp 0
transform -1 0 7570 0 1 14170
box -6 -8 26 248
use FILL  FILL_1__14151_
timestamp 0
transform -1 0 7610 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__14152_
timestamp 0
transform -1 0 7770 0 1 13210
box -6 -8 26 248
use FILL  FILL_1__14153_
timestamp 0
transform 1 0 7170 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1__14154_
timestamp 0
transform -1 0 6970 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__14155_
timestamp 0
transform 1 0 7430 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1__14156_
timestamp 0
transform 1 0 7250 0 1 15610
box -6 -8 26 248
use FILL  FILL_1__14157_
timestamp 0
transform -1 0 11090 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__14158_
timestamp 0
transform 1 0 10930 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1__14216_
timestamp 0
transform 1 0 7470 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__14217_
timestamp 0
transform 1 0 7690 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__14218_
timestamp 0
transform -1 0 7710 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14219_
timestamp 0
transform -1 0 7530 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14220_
timestamp 0
transform 1 0 7650 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14221_
timestamp 0
transform 1 0 7510 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14222_
timestamp 0
transform -1 0 7430 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14223_
timestamp 0
transform -1 0 6910 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14224_
timestamp 0
transform 1 0 7030 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14225_
timestamp 0
transform 1 0 6830 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__14226_
timestamp 0
transform -1 0 7210 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__14227_
timestamp 0
transform 1 0 7170 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14228_
timestamp 0
transform -1 0 8530 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__14229_
timestamp 0
transform 1 0 7950 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__14230_
timestamp 0
transform -1 0 8370 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__14231_
timestamp 0
transform -1 0 10230 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__14232_
timestamp 0
transform -1 0 9950 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__14233_
timestamp 0
transform -1 0 10090 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__14234_
timestamp 0
transform -1 0 8990 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__14235_
timestamp 0
transform 1 0 8530 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__14236_
timestamp 0
transform 1 0 8430 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__14237_
timestamp 0
transform -1 0 8870 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__14238_
timestamp 0
transform -1 0 7890 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__14239_
timestamp 0
transform -1 0 8010 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__14240_
timestamp 0
transform -1 0 8450 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__14241_
timestamp 0
transform -1 0 8330 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__14242_
timestamp 0
transform -1 0 8290 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__14243_
timestamp 0
transform -1 0 8370 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14244_
timestamp 0
transform 1 0 6890 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14245_
timestamp 0
transform -1 0 6770 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14246_
timestamp 0
transform 1 0 9470 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14247_
timestamp 0
transform 1 0 8710 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__14248_
timestamp 0
transform 1 0 8570 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__14249_
timestamp 0
transform 1 0 9810 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__14250_
timestamp 0
transform 1 0 9990 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14251_
timestamp 0
transform 1 0 9830 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14252_
timestamp 0
transform 1 0 7590 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__14253_
timestamp 0
transform 1 0 7810 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__14254_
timestamp 0
transform 1 0 7650 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14255_
timestamp 0
transform 1 0 7510 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14256_
timestamp 0
transform 1 0 7150 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14257_
timestamp 0
transform -1 0 8110 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14258_
timestamp 0
transform 1 0 7050 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__14259_
timestamp 0
transform -1 0 7170 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__14260_
timestamp 0
transform 1 0 7310 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14261_
timestamp 0
transform 1 0 7730 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14262_
timestamp 0
transform 1 0 7590 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14263_
timestamp 0
transform -1 0 7810 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14264_
timestamp 0
transform 1 0 7010 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14265_
timestamp 0
transform -1 0 7030 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14266_
timestamp 0
transform -1 0 6930 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__14267_
timestamp 0
transform -1 0 7170 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14268_
timestamp 0
transform -1 0 6890 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14269_
timestamp 0
transform 1 0 7070 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__14270_
timestamp 0
transform 1 0 6910 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__14271_
timestamp 0
transform -1 0 7310 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14272_
timestamp 0
transform -1 0 7450 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14273_
timestamp 0
transform 1 0 7550 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14274_
timestamp 0
transform -1 0 7730 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14275_
timestamp 0
transform 1 0 7270 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14276_
timestamp 0
transform -1 0 7710 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14277_
timestamp 0
transform -1 0 7930 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14278_
timestamp 0
transform -1 0 7970 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14279_
timestamp 0
transform 1 0 9310 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14280_
timestamp 0
transform -1 0 9250 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14281_
timestamp 0
transform 1 0 8030 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14282_
timestamp 0
transform -1 0 9370 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14283_
timestamp 0
transform 1 0 9450 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14284_
timestamp 0
transform 1 0 8270 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14285_
timestamp 0
transform -1 0 8410 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14286_
timestamp 0
transform 1 0 8210 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__14287_
timestamp 0
transform -1 0 9170 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14288_
timestamp 0
transform 1 0 8230 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14289_
timestamp 0
transform 1 0 8070 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14290_
timestamp 0
transform 1 0 7930 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14291_
timestamp 0
transform -1 0 8090 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14292_
timestamp 0
transform -1 0 8190 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14293_
timestamp 0
transform 1 0 9210 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14294_
timestamp 0
transform -1 0 9230 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14295_
timestamp 0
transform 1 0 8970 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14296_
timestamp 0
transform 1 0 9090 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14297_
timestamp 0
transform 1 0 9070 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14298_
timestamp 0
transform -1 0 9130 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14299_
timestamp 0
transform -1 0 8830 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14300_
timestamp 0
transform -1 0 9110 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14301_
timestamp 0
transform 1 0 7830 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__14302_
timestamp 0
transform -1 0 8850 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14303_
timestamp 0
transform -1 0 8890 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14304_
timestamp 0
transform -1 0 8990 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14305_
timestamp 0
transform 1 0 8690 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14306_
timestamp 0
transform -1 0 8830 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14307_
timestamp 0
transform 1 0 8730 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14308_
timestamp 0
transform 1 0 8130 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14309_
timestamp 0
transform 1 0 9370 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14310_
timestamp 0
transform -1 0 8330 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14311_
timestamp 0
transform -1 0 8350 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14312_
timestamp 0
transform 1 0 8470 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14313_
timestamp 0
transform -1 0 9650 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14314_
timestamp 0
transform -1 0 9530 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14315_
timestamp 0
transform 1 0 9570 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14316_
timestamp 0
transform 1 0 8670 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14317_
timestamp 0
transform -1 0 8690 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__14318_
timestamp 0
transform 1 0 8430 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14319_
timestamp 0
transform -1 0 9030 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14320_
timestamp 0
transform -1 0 9710 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14321_
timestamp 0
transform -1 0 8750 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14322_
timestamp 0
transform -1 0 8890 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14323_
timestamp 0
transform 1 0 8550 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14324_
timestamp 0
transform 1 0 8910 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__14325_
timestamp 0
transform 1 0 8430 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14326_
timestamp 0
transform -1 0 8630 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14327_
timestamp 0
transform 1 0 8710 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14328_
timestamp 0
transform 1 0 8850 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14329_
timestamp 0
transform -1 0 8810 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__14330_
timestamp 0
transform 1 0 9010 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14331_
timestamp 0
transform -1 0 9170 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14332_
timestamp 0
transform -1 0 9290 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14333_
timestamp 0
transform 1 0 8950 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14334_
timestamp 0
transform -1 0 9710 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__14335_
timestamp 0
transform -1 0 8650 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__14336_
timestamp 0
transform 1 0 8510 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__14337_
timestamp 0
transform -1 0 8410 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__14338_
timestamp 0
transform 1 0 8850 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__14339_
timestamp 0
transform 1 0 9010 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__14340_
timestamp 0
transform -1 0 9010 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__14341_
timestamp 0
transform -1 0 8870 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__14342_
timestamp 0
transform 1 0 9130 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__14343_
timestamp 0
transform 1 0 8710 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__14344_
timestamp 0
transform 1 0 8970 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__14345_
timestamp 0
transform 1 0 9290 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__14346_
timestamp 0
transform 1 0 9410 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__14347_
timestamp 0
transform -1 0 9570 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__14348_
timestamp 0
transform 1 0 8010 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14349_
timestamp 0
transform 1 0 7850 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14350_
timestamp 0
transform -1 0 8170 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14351_
timestamp 0
transform -1 0 7690 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14352_
timestamp 0
transform -1 0 7450 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14353_
timestamp 0
transform -1 0 7550 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14354_
timestamp 0
transform -1 0 8010 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14355_
timestamp 0
transform 1 0 7850 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14356_
timestamp 0
transform 1 0 8290 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14357_
timestamp 0
transform -1 0 8310 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14358_
timestamp 0
transform 1 0 8310 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14359_
timestamp 0
transform 1 0 8430 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14360_
timestamp 0
transform -1 0 8430 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14361_
timestamp 0
transform 1 0 8450 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14362_
timestamp 0
transform 1 0 7550 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__14363_
timestamp 0
transform 1 0 8130 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14364_
timestamp 0
transform -1 0 8030 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14365_
timestamp 0
transform -1 0 7890 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14366_
timestamp 0
transform 1 0 8030 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14367_
timestamp 0
transform 1 0 7310 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14368_
timestamp 0
transform -1 0 9410 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14369_
timestamp 0
transform 1 0 8570 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14370_
timestamp 0
transform 1 0 8550 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14371_
timestamp 0
transform -1 0 9650 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14372_
timestamp 0
transform -1 0 10830 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14373_
timestamp 0
transform 1 0 8670 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14374_
timestamp 0
transform 1 0 10350 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14375_
timestamp 0
transform 1 0 10370 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14376_
timestamp 0
transform 1 0 8870 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__14377_
timestamp 0
transform 1 0 9990 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14378_
timestamp 0
transform 1 0 10950 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14379_
timestamp 0
transform 1 0 11270 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14380_
timestamp 0
transform -1 0 11130 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14381_
timestamp 0
transform 1 0 11030 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14382_
timestamp 0
transform 1 0 9510 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14383_
timestamp 0
transform -1 0 10210 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14384_
timestamp 0
transform 1 0 10490 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14385_
timestamp 0
transform 1 0 10710 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14386_
timestamp 0
transform -1 0 10790 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14387_
timestamp 0
transform 1 0 10630 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14388_
timestamp 0
transform -1 0 10550 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14389_
timestamp 0
transform 1 0 9070 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__14390_
timestamp 0
transform -1 0 10330 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14391_
timestamp 0
transform 1 0 10470 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14392_
timestamp 0
transform 1 0 10610 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14393_
timestamp 0
transform 1 0 11050 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14394_
timestamp 0
transform -1 0 10910 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14395_
timestamp 0
transform 1 0 10670 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14396_
timestamp 0
transform 1 0 9570 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14397_
timestamp 0
transform 1 0 9770 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14398_
timestamp 0
transform -1 0 9970 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14399_
timestamp 0
transform 1 0 10570 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14400_
timestamp 0
transform -1 0 10010 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14401_
timestamp 0
transform 1 0 9990 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14402_
timestamp 0
transform 1 0 10070 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14403_
timestamp 0
transform 1 0 10130 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14404_
timestamp 0
transform -1 0 8950 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__14405_
timestamp 0
transform -1 0 9170 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14406_
timestamp 0
transform 1 0 10250 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14407_
timestamp 0
transform 1 0 9850 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__14408_
timestamp 0
transform -1 0 8870 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14409_
timestamp 0
transform -1 0 9010 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14410_
timestamp 0
transform 1 0 8690 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14411_
timestamp 0
transform -1 0 10430 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14412_
timestamp 0
transform 1 0 10130 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14413_
timestamp 0
transform 1 0 10250 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14414_
timestamp 0
transform 1 0 9090 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14415_
timestamp 0
transform 1 0 8890 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__14416_
timestamp 0
transform 1 0 9850 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14417_
timestamp 0
transform 1 0 9430 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14418_
timestamp 0
transform -1 0 9250 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14419_
timestamp 0
transform -1 0 9430 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14420_
timestamp 0
transform 1 0 9790 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14421_
timestamp 0
transform -1 0 8170 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__14422_
timestamp 0
transform -1 0 8290 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__14423_
timestamp 0
transform 1 0 8970 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__14424_
timestamp 0
transform 1 0 9270 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__14425_
timestamp 0
transform 1 0 9590 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14426_
timestamp 0
transform -1 0 8990 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__14427_
timestamp 0
transform 1 0 9710 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__14428_
timestamp 0
transform -1 0 10050 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14429_
timestamp 0
transform -1 0 9910 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__14430_
timestamp 0
transform 1 0 9790 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14431_
timestamp 0
transform -1 0 9950 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14432_
timestamp 0
transform 1 0 9910 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14433_
timestamp 0
transform 1 0 8030 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__14434_
timestamp 0
transform -1 0 8410 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__14435_
timestamp 0
transform 1 0 8490 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__14436_
timestamp 0
transform 1 0 7890 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__14437_
timestamp 0
transform -1 0 8130 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__14438_
timestamp 0
transform -1 0 8370 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__14439_
timestamp 0
transform 1 0 8470 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__14440_
timestamp 0
transform 1 0 9130 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__14441_
timestamp 0
transform -1 0 9150 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__14442_
timestamp 0
transform 1 0 8310 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__14443_
timestamp 0
transform -1 0 8470 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__14444_
timestamp 0
transform 1 0 9010 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__14445_
timestamp 0
transform -1 0 8770 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__14446_
timestamp 0
transform 1 0 8890 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__14447_
timestamp 0
transform 1 0 8650 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__14448_
timestamp 0
transform 1 0 8510 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__14449_
timestamp 0
transform 1 0 8010 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__14450_
timestamp 0
transform 1 0 9070 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__14451_
timestamp 0
transform 1 0 8930 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__14452_
timestamp 0
transform 1 0 8870 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__14453_
timestamp 0
transform 1 0 8290 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__14454_
timestamp 0
transform 1 0 8130 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__14455_
timestamp 0
transform 1 0 8590 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14456_
timestamp 0
transform 1 0 8550 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__14457_
timestamp 0
transform 1 0 8250 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__14458_
timestamp 0
transform 1 0 8350 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__14459_
timestamp 0
transform 1 0 8130 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__14460_
timestamp 0
transform -1 0 8010 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__14461_
timestamp 0
transform 1 0 8170 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__14462_
timestamp 0
transform 1 0 8030 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__14463_
timestamp 0
transform 1 0 8210 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__14464_
timestamp 0
transform -1 0 7950 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__14465_
timestamp 0
transform -1 0 8090 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__14466_
timestamp 0
transform -1 0 7730 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__14467_
timestamp 0
transform -1 0 7890 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__14468_
timestamp 0
transform 1 0 7890 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__14469_
timestamp 0
transform 1 0 7750 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__14470_
timestamp 0
transform -1 0 7370 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__14471_
timestamp 0
transform 1 0 7150 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__14472_
timestamp 0
transform 1 0 9350 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__14473_
timestamp 0
transform 1 0 9190 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__14474_
timestamp 0
transform 1 0 7770 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__14475_
timestamp 0
transform -1 0 8010 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__14476_
timestamp 0
transform 1 0 9470 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__14477_
timestamp 0
transform -1 0 9130 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__14478_
timestamp 0
transform -1 0 9250 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__14479_
timestamp 0
transform -1 0 7790 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__14480_
timestamp 0
transform 1 0 9710 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__14481_
timestamp 0
transform 1 0 9570 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__14482_
timestamp 0
transform 1 0 9970 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__14483_
timestamp 0
transform 1 0 9810 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__14484_
timestamp 0
transform 1 0 9910 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__14485_
timestamp 0
transform 1 0 9510 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__14486_
timestamp 0
transform 1 0 9850 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__14487_
timestamp 0
transform 1 0 9870 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__14488_
timestamp 0
transform -1 0 9530 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__14489_
timestamp 0
transform 1 0 9370 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__14490_
timestamp 0
transform 1 0 8390 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__14491_
timestamp 0
transform -1 0 8570 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__14492_
timestamp 0
transform 1 0 8230 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__14493_
timestamp 0
transform 1 0 8090 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__14494_
timestamp 0
transform -1 0 7490 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__14495_
timestamp 0
transform -1 0 7630 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__14496_
timestamp 0
transform 1 0 7410 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__14497_
timestamp 0
transform -1 0 7330 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__14498_
timestamp 0
transform 1 0 9550 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__14499_
timestamp 0
transform -1 0 9570 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__14556_
timestamp 0
transform -1 0 14750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__14557_
timestamp 0
transform -1 0 14490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__14558_
timestamp 0
transform -1 0 14050 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14559_
timestamp 0
transform -1 0 12930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14560_
timestamp 0
transform -1 0 12150 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14561_
timestamp 0
transform -1 0 13070 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14562_
timestamp 0
transform 1 0 11710 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14563_
timestamp 0
transform -1 0 12010 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14564_
timestamp 0
transform -1 0 12530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14565_
timestamp 0
transform -1 0 12650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14566_
timestamp 0
transform -1 0 14570 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14567_
timestamp 0
transform -1 0 14590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__14568_
timestamp 0
transform -1 0 15470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__14569_
timestamp 0
transform 1 0 15070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__14570_
timestamp 0
transform 1 0 15050 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__14571_
timestamp 0
transform 1 0 14070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__14572_
timestamp 0
transform -1 0 14130 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__14573_
timestamp 0
transform -1 0 12510 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14574_
timestamp 0
transform 1 0 11650 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14575_
timestamp 0
transform 1 0 11850 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14576_
timestamp 0
transform -1 0 13330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14577_
timestamp 0
transform -1 0 13170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14578_
timestamp 0
transform 1 0 13010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14579_
timestamp 0
transform -1 0 13410 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14580_
timestamp 0
transform -1 0 12990 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14581_
timestamp 0
transform 1 0 14330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__14582_
timestamp 0
transform -1 0 14210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__14583_
timestamp 0
transform -1 0 13810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__14584_
timestamp 0
transform -1 0 13930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__14585_
timestamp 0
transform -1 0 12370 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14586_
timestamp 0
transform -1 0 9750 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14587_
timestamp 0
transform -1 0 10010 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14588_
timestamp 0
transform 1 0 10030 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14589_
timestamp 0
transform -1 0 9910 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14590_
timestamp 0
transform 1 0 9870 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14591_
timestamp 0
transform -1 0 11990 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14592_
timestamp 0
transform 1 0 11970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14593_
timestamp 0
transform 1 0 13030 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14594_
timestamp 0
transform -1 0 13950 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14595_
timestamp 0
transform 1 0 11290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14596_
timestamp 0
transform 1 0 14270 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__14597_
timestamp 0
transform -1 0 14930 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__14598_
timestamp 0
transform 1 0 13790 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14599_
timestamp 0
transform -1 0 12810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14600_
timestamp 0
transform -1 0 12950 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14601_
timestamp 0
transform -1 0 11850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14602_
timestamp 0
transform 1 0 14910 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14603_
timestamp 0
transform 1 0 15310 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14604_
timestamp 0
transform 1 0 15170 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14605_
timestamp 0
transform -1 0 15030 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14606_
timestamp 0
transform -1 0 14570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14607_
timestamp 0
transform -1 0 14970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14608_
timestamp 0
transform -1 0 14850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14609_
timestamp 0
transform 1 0 15070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14610_
timestamp 0
transform -1 0 15770 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14611_
timestamp 0
transform 1 0 16030 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14612_
timestamp 0
transform 1 0 16170 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14613_
timestamp 0
transform 1 0 16310 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14614_
timestamp 0
transform 1 0 15910 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14615_
timestamp 0
transform 1 0 15190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14616_
timestamp 0
transform -1 0 15630 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14617_
timestamp 0
transform -1 0 14690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14618_
timestamp 0
transform 1 0 13730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14619_
timestamp 0
transform -1 0 13630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14620_
timestamp 0
transform 1 0 14330 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14621_
timestamp 0
transform -1 0 14210 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14622_
timestamp 0
transform 1 0 13910 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14623_
timestamp 0
transform -1 0 14070 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14624_
timestamp 0
transform -1 0 13790 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14625_
timestamp 0
transform -1 0 13950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14626_
timestamp 0
transform 1 0 13870 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14627_
timestamp 0
transform 1 0 14670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14628_
timestamp 0
transform -1 0 14570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14629_
timestamp 0
transform 1 0 14410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14630_
timestamp 0
transform 1 0 13990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14631_
timestamp 0
transform -1 0 14150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14632_
timestamp 0
transform -1 0 14290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14633_
timestamp 0
transform -1 0 13890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14634_
timestamp 0
transform -1 0 13730 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14635_
timestamp 0
transform 1 0 14470 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14636_
timestamp 0
transform 1 0 14610 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14637_
timestamp 0
transform 1 0 14730 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14638_
timestamp 0
transform 1 0 14990 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14639_
timestamp 0
transform 1 0 15510 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14640_
timestamp 0
transform -1 0 15410 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14641_
timestamp 0
transform -1 0 15690 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14642_
timestamp 0
transform -1 0 14890 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14643_
timestamp 0
transform 1 0 15830 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14644_
timestamp 0
transform 1 0 16010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14645_
timestamp 0
transform -1 0 15910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14646_
timestamp 0
transform -1 0 15610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14647_
timestamp 0
transform 1 0 15750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14648_
timestamp 0
transform 1 0 16130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14649_
timestamp 0
transform -1 0 17050 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14650_
timestamp 0
transform 1 0 16870 0 1 16570
box -6 -8 26 248
use FILL  FILL_1__14651_
timestamp 0
transform 1 0 16950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14652_
timestamp 0
transform -1 0 16570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14653_
timestamp 0
transform 1 0 16410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14654_
timestamp 0
transform 1 0 16290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14655_
timestamp 0
transform -1 0 16810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14656_
timestamp 0
transform 1 0 16650 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14657_
timestamp 0
transform 1 0 16390 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14658_
timestamp 0
transform 1 0 16670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14659_
timestamp 0
transform -1 0 16510 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14660_
timestamp 0
transform 1 0 16090 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14661_
timestamp 0
transform 1 0 16250 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14662_
timestamp 0
transform -1 0 16890 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14663_
timestamp 0
transform 1 0 17010 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14664_
timestamp 0
transform 1 0 16650 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14665_
timestamp 0
transform 1 0 17030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14666_
timestamp 0
transform 1 0 16770 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14667_
timestamp 0
transform 1 0 17010 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14668_
timestamp 0
transform 1 0 16870 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14669_
timestamp 0
transform 1 0 16910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14670_
timestamp 0
transform -1 0 16630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14671_
timestamp 0
transform -1 0 16790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14672_
timestamp 0
transform -1 0 16730 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14673_
timestamp 0
transform -1 0 16090 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14674_
timestamp 0
transform -1 0 16350 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14675_
timestamp 0
transform 1 0 16210 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14676_
timestamp 0
transform 1 0 16110 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14677_
timestamp 0
transform -1 0 15970 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14678_
timestamp 0
transform 1 0 16270 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14679_
timestamp 0
transform 1 0 16250 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14680_
timestamp 0
transform -1 0 15990 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14681_
timestamp 0
transform 1 0 16490 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14682_
timestamp 0
transform -1 0 15950 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14683_
timestamp 0
transform 1 0 16630 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14684_
timestamp 0
transform -1 0 16570 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14685_
timestamp 0
transform 1 0 15950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14686_
timestamp 0
transform -1 0 16790 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14687_
timestamp 0
transform -1 0 16650 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14688_
timestamp 0
transform -1 0 16430 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14689_
timestamp 0
transform 1 0 16350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14690_
timestamp 0
transform -1 0 16490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14691_
timestamp 0
transform -1 0 15810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14692_
timestamp 0
transform -1 0 14350 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14693_
timestamp 0
transform 1 0 14450 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14694_
timestamp 0
transform -1 0 14770 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14695_
timestamp 0
transform -1 0 14950 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14696_
timestamp 0
transform 1 0 14670 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14697_
timestamp 0
transform 1 0 14810 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14698_
timestamp 0
transform -1 0 14850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14699_
timestamp 0
transform 1 0 14990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14700_
timestamp 0
transform -1 0 14630 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14701_
timestamp 0
transform 1 0 14830 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14702_
timestamp 0
transform -1 0 14550 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14703_
timestamp 0
transform -1 0 14310 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14704_
timestamp 0
transform -1 0 14430 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14705_
timestamp 0
transform 1 0 14970 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14706_
timestamp 0
transform 1 0 14210 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14707_
timestamp 0
transform -1 0 14110 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14708_
timestamp 0
transform -1 0 13970 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14709_
timestamp 0
transform 1 0 14010 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14710_
timestamp 0
transform 1 0 14150 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14711_
timestamp 0
transform -1 0 14650 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14712_
timestamp 0
transform 1 0 15110 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14713_
timestamp 0
transform 1 0 15250 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14714_
timestamp 0
transform 1 0 14990 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14715_
timestamp 0
transform 1 0 15130 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14716_
timestamp 0
transform -1 0 15550 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14717_
timestamp 0
transform 1 0 15670 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14718_
timestamp 0
transform -1 0 15550 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14719_
timestamp 0
transform -1 0 15310 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14720_
timestamp 0
transform 1 0 15530 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14721_
timestamp 0
transform 1 0 15410 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14722_
timestamp 0
transform 1 0 15450 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14723_
timestamp 0
transform -1 0 15330 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14724_
timestamp 0
transform -1 0 15830 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14725_
timestamp 0
transform -1 0 15710 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14726_
timestamp 0
transform -1 0 15670 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14727_
timestamp 0
transform 1 0 15790 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14728_
timestamp 0
transform 1 0 15410 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14729_
timestamp 0
transform 1 0 16090 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14730_
timestamp 0
transform 1 0 15950 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14731_
timestamp 0
transform 1 0 15810 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14732_
timestamp 0
transform 1 0 15990 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14733_
timestamp 0
transform -1 0 15870 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14734_
timestamp 0
transform 1 0 12750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14735_
timestamp 0
transform 1 0 14870 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14736_
timestamp 0
transform -1 0 15390 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14737_
timestamp 0
transform -1 0 15030 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14738_
timestamp 0
transform -1 0 15330 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14739_
timestamp 0
transform -1 0 15170 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14740_
timestamp 0
transform -1 0 14770 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14741_
timestamp 0
transform 1 0 14670 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14742_
timestamp 0
transform 1 0 12170 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14743_
timestamp 0
transform -1 0 12030 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14744_
timestamp 0
transform 1 0 11890 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14745_
timestamp 0
transform -1 0 12450 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14746_
timestamp 0
transform -1 0 12570 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14747_
timestamp 0
transform -1 0 12410 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14748_
timestamp 0
transform -1 0 12610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14749_
timestamp 0
transform -1 0 11670 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14750_
timestamp 0
transform -1 0 11770 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14751_
timestamp 0
transform -1 0 11250 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14752_
timestamp 0
transform 1 0 12150 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14753_
timestamp 0
transform 1 0 12290 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14754_
timestamp 0
transform -1 0 12110 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14755_
timestamp 0
transform 1 0 12230 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14756_
timestamp 0
transform -1 0 11830 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14757_
timestamp 0
transform -1 0 11970 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14758_
timestamp 0
transform 1 0 12710 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14759_
timestamp 0
transform -1 0 11390 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14760_
timestamp 0
transform -1 0 11510 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14761_
timestamp 0
transform 1 0 12710 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14762_
timestamp 0
transform 1 0 12430 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14763_
timestamp 0
transform -1 0 12310 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14764_
timestamp 0
transform 1 0 12570 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14765_
timestamp 0
transform 1 0 13410 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14766_
timestamp 0
transform 1 0 12850 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14767_
timestamp 0
transform 1 0 12990 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14768_
timestamp 0
transform 1 0 12770 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14769_
timestamp 0
transform -1 0 12790 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14770_
timestamp 0
transform 1 0 12850 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14771_
timestamp 0
transform -1 0 13610 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14772_
timestamp 0
transform 1 0 13470 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14773_
timestamp 0
transform -1 0 13870 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14774_
timestamp 0
transform -1 0 13730 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14775_
timestamp 0
transform -1 0 13150 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14776_
timestamp 0
transform -1 0 13290 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14777_
timestamp 0
transform 1 0 13970 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14778_
timestamp 0
transform -1 0 13370 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14779_
timestamp 0
transform -1 0 13210 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14780_
timestamp 0
transform -1 0 12930 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14781_
timestamp 0
transform -1 0 13070 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14782_
timestamp 0
transform 1 0 12990 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14783_
timestamp 0
transform 1 0 13270 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14784_
timestamp 0
transform -1 0 14390 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14785_
timestamp 0
transform 1 0 14890 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14786_
timestamp 0
transform 1 0 13570 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14787_
timestamp 0
transform 1 0 13570 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14788_
timestamp 0
transform 1 0 13130 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14789_
timestamp 0
transform 1 0 13410 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14790_
timestamp 0
transform -1 0 13730 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14791_
timestamp 0
transform 1 0 13970 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14792_
timestamp 0
transform -1 0 14110 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14793_
timestamp 0
transform -1 0 10970 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14794_
timestamp 0
transform 1 0 11090 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14795_
timestamp 0
transform 1 0 11490 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14796_
timestamp 0
transform 1 0 11610 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14797_
timestamp 0
transform 1 0 16150 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14798_
timestamp 0
transform 1 0 16070 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14799_
timestamp 0
transform 1 0 16210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14800_
timestamp 0
transform -1 0 15670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14801_
timestamp 0
transform 1 0 14530 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14802_
timestamp 0
transform 1 0 13830 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14803_
timestamp 0
transform -1 0 14150 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14804_
timestamp 0
transform -1 0 14250 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14805_
timestamp 0
transform 1 0 11870 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14806_
timestamp 0
transform -1 0 11770 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14807_
timestamp 0
transform -1 0 11530 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14808_
timestamp 0
transform -1 0 11670 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14809_
timestamp 0
transform 1 0 11190 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14810_
timestamp 0
transform 1 0 10790 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14811_
timestamp 0
transform 1 0 10670 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14812_
timestamp 0
transform -1 0 10570 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14813_
timestamp 0
transform 1 0 11330 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14814_
timestamp 0
transform 1 0 11230 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14815_
timestamp 0
transform -1 0 11090 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14816_
timestamp 0
transform 1 0 11370 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14817_
timestamp 0
transform -1 0 11070 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14818_
timestamp 0
transform -1 0 10430 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14819_
timestamp 0
transform -1 0 10930 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14820_
timestamp 0
transform -1 0 10270 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14821_
timestamp 0
transform 1 0 10130 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14822_
timestamp 0
transform 1 0 10370 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14823_
timestamp 0
transform -1 0 9930 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14824_
timestamp 0
transform 1 0 10790 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14825_
timestamp 0
transform -1 0 10210 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14826_
timestamp 0
transform -1 0 10330 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14827_
timestamp 0
transform -1 0 10050 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14828_
timestamp 0
transform 1 0 9770 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14829_
timestamp 0
transform -1 0 10110 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14830_
timestamp 0
transform 1 0 10630 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14831_
timestamp 0
transform 1 0 10350 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14832_
timestamp 0
transform -1 0 10910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14833_
timestamp 0
transform 1 0 10650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14834_
timestamp 0
transform -1 0 9530 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14835_
timestamp 0
transform -1 0 9650 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14836_
timestamp 0
transform -1 0 9130 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14837_
timestamp 0
transform 1 0 9250 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14838_
timestamp 0
transform -1 0 9410 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14839_
timestamp 0
transform 1 0 10510 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14840_
timestamp 0
transform -1 0 10670 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14841_
timestamp 0
transform 1 0 10230 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14842_
timestamp 0
transform 1 0 10490 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14843_
timestamp 0
transform -1 0 10550 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14844_
timestamp 0
transform -1 0 12250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14845_
timestamp 0
transform -1 0 12330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14846_
timestamp 0
transform 1 0 12370 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14847_
timestamp 0
transform -1 0 11670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14848_
timestamp 0
transform -1 0 13470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14849_
timestamp 0
transform 1 0 11770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14850_
timestamp 0
transform -1 0 15270 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14851_
timestamp 0
transform 1 0 15450 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14852_
timestamp 0
transform -1 0 13650 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14853_
timestamp 0
transform -1 0 13330 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14854_
timestamp 0
transform 1 0 12830 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14855_
timestamp 0
transform 1 0 14390 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__14856_
timestamp 0
transform -1 0 12170 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14857_
timestamp 0
transform 1 0 12450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14858_
timestamp 0
transform 1 0 13030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14859_
timestamp 0
transform 1 0 13790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14860_
timestamp 0
transform -1 0 13490 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14861_
timestamp 0
transform 1 0 13410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__14862_
timestamp 0
transform 1 0 12010 0 1 730
box -6 -8 26 248
use FILL  FILL_1__14863_
timestamp 0
transform 1 0 12150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14864_
timestamp 0
transform 1 0 10770 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14865_
timestamp 0
transform -1 0 10930 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__14866_
timestamp 0
transform 1 0 11590 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14867_
timestamp 0
transform 1 0 11010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__14868_
timestamp 0
transform -1 0 11250 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__14908_
timestamp 0
transform -1 0 7610 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__14909_
timestamp 0
transform -1 0 50 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__14910_
timestamp 0
transform -1 0 8510 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14911_
timestamp 0
transform -1 0 9770 0 1 250
box -6 -8 26 248
use FILL  FILL_1__14912_
timestamp 0
transform -1 0 6790 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14913_
timestamp 0
transform -1 0 50 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__14914_
timestamp 0
transform 1 0 8230 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__14915_
timestamp 0
transform 1 0 16190 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__14916_
timestamp 0
transform 1 0 8430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__14917_
timestamp 0
transform -1 0 7970 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__14918_
timestamp 0
transform -1 0 8110 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__14919_
timestamp 0
transform -1 0 6310 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__14920_
timestamp 0
transform 1 0 8990 0 -1 250
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert0
timestamp 0
transform 1 0 8210 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert1
timestamp 0
transform 1 0 9490 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert2
timestamp 0
transform -1 0 7850 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert3
timestamp 0
transform 1 0 9450 0 1 8410
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert4
timestamp 0
transform -1 0 9350 0 1 8410
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert5
timestamp 0
transform 1 0 5410 0 1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert6
timestamp 0
transform 1 0 4630 0 1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert7
timestamp 0
transform -1 0 1330 0 1 10810
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert8
timestamp 0
transform -1 0 1170 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert9
timestamp 0
transform 1 0 4530 0 1 6010
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert10
timestamp 0
transform 1 0 4130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert11
timestamp 0
transform 1 0 3590 0 1 6010
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert12
timestamp 0
transform -1 0 3310 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert13
timestamp 0
transform -1 0 4430 0 1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert14
timestamp 0
transform -1 0 4110 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert15
timestamp 0
transform 1 0 6850 0 1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert16
timestamp 0
transform -1 0 4790 0 1 7450
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert17
timestamp 0
transform -1 0 3230 0 1 7450
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert18
timestamp 0
transform -1 0 4530 0 1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert19
timestamp 0
transform -1 0 16150 0 1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert20
timestamp 0
transform -1 0 16270 0 1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert21
timestamp 0
transform -1 0 12890 0 1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert22
timestamp 0
transform -1 0 12110 0 1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert23
timestamp 0
transform -1 0 3030 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert24
timestamp 0
transform 1 0 4670 0 1 10330
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert25
timestamp 0
transform 1 0 1050 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert26
timestamp 0
transform -1 0 50 0 1 10810
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert27
timestamp 0
transform -1 0 1190 0 1 10810
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert28
timestamp 0
transform -1 0 50 0 1 10330
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert108
timestamp 0
transform -1 0 7810 0 1 7450
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert109
timestamp 0
transform 1 0 9290 0 1 7450
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert110
timestamp 0
transform -1 0 9030 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert111
timestamp 0
transform 1 0 8810 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert112
timestamp 0
transform 1 0 8310 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert113
timestamp 0
transform -1 0 13850 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert114
timestamp 0
transform -1 0 13530 0 1 13210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert115
timestamp 0
transform -1 0 14350 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert116
timestamp 0
transform 1 0 15090 0 1 14650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert117
timestamp 0
transform -1 0 6970 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert118
timestamp 0
transform 1 0 8150 0 1 6490
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert119
timestamp 0
transform 1 0 7710 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert120
timestamp 0
transform 1 0 7090 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert121
timestamp 0
transform -1 0 5810 0 1 6490
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert122
timestamp 0
transform -1 0 7590 0 1 6010
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert123
timestamp 0
transform 1 0 7750 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert124
timestamp 0
transform -1 0 6590 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert125
timestamp 0
transform -1 0 6010 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert126
timestamp 0
transform 1 0 5350 0 1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert127
timestamp 0
transform -1 0 4090 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert128
timestamp 0
transform 1 0 4610 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert129
timestamp 0
transform -1 0 4190 0 1 7450
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert130
timestamp 0
transform -1 0 5110 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert131
timestamp 0
transform -1 0 2570 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert132
timestamp 0
transform 1 0 2670 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert133
timestamp 0
transform 1 0 890 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert134
timestamp 0
transform -1 0 430 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert135
timestamp 0
transform 1 0 610 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert136
timestamp 0
transform 1 0 13590 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert137
timestamp 0
transform -1 0 11910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert138
timestamp 0
transform -1 0 12050 0 1 250
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert139
timestamp 0
transform 1 0 15510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert140
timestamp 0
transform 1 0 14550 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert141
timestamp 0
transform -1 0 10970 0 1 11290
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert142
timestamp 0
transform 1 0 12130 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert143
timestamp 0
transform -1 0 11310 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert144
timestamp 0
transform 1 0 12190 0 1 11290
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert145
timestamp 0
transform 1 0 12310 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert146
timestamp 0
transform -1 0 10530 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert147
timestamp 0
transform 1 0 10650 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert148
timestamp 0
transform 1 0 8490 0 1 250
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert149
timestamp 0
transform 1 0 8090 0 -1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert150
timestamp 0
transform -1 0 7930 0 1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert151
timestamp 0
transform -1 0 16070 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert152
timestamp 0
transform 1 0 16050 0 1 13690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert153
timestamp 0
transform -1 0 15930 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert154
timestamp 0
transform -1 0 15930 0 1 12730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert155
timestamp 0
transform -1 0 15990 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert156
timestamp 0
transform -1 0 15730 0 1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert157
timestamp 0
transform -1 0 15030 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert158
timestamp 0
transform 1 0 16950 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert159
timestamp 0
transform 1 0 15890 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert160
timestamp 0
transform 1 0 16410 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert161
timestamp 0
transform 1 0 11950 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert162
timestamp 0
transform 1 0 12730 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert163
timestamp 0
transform 1 0 12730 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert164
timestamp 0
transform -1 0 10530 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert165
timestamp 0
transform -1 0 11690 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert166
timestamp 0
transform -1 0 1190 0 1 9850
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert167
timestamp 0
transform -1 0 1150 0 1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert168
timestamp 0
transform 1 0 3650 0 1 9850
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert169
timestamp 0
transform 1 0 3710 0 1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert170
timestamp 0
transform 1 0 1510 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert171
timestamp 0
transform -1 0 14430 0 1 12730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert172
timestamp 0
transform 1 0 12850 0 1 12730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert173
timestamp 0
transform -1 0 11950 0 1 13690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert174
timestamp 0
transform -1 0 12110 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert175
timestamp 0
transform 1 0 14750 0 1 12250
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert176
timestamp 0
transform -1 0 14030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert177
timestamp 0
transform 1 0 15850 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert178
timestamp 0
transform -1 0 14050 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert179
timestamp 0
transform 1 0 15830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert180
timestamp 0
transform 1 0 15250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert181
timestamp 0
transform 1 0 11490 0 1 6490
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert182
timestamp 0
transform -1 0 10050 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert183
timestamp 0
transform 1 0 11730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert184
timestamp 0
transform 1 0 11810 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert185
timestamp 0
transform -1 0 10330 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert186
timestamp 0
transform -1 0 6010 0 1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert187
timestamp 0
transform 1 0 8230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert188
timestamp 0
transform -1 0 6830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert189
timestamp 0
transform -1 0 5970 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert190
timestamp 0
transform 1 0 9610 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert191
timestamp 0
transform 1 0 12510 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert192
timestamp 0
transform 1 0 12390 0 1 14650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert193
timestamp 0
transform 1 0 12130 0 1 15130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert194
timestamp 0
transform -1 0 11430 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert195
timestamp 0
transform -1 0 11850 0 1 14170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert196
timestamp 0
transform -1 0 1390 0 1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert197
timestamp 0
transform -1 0 1870 0 1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert198
timestamp 0
transform -1 0 730 0 1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert199
timestamp 0
transform 1 0 1890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert200
timestamp 0
transform 1 0 12750 0 1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert201
timestamp 0
transform -1 0 11890 0 1 10810
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert202
timestamp 0
transform 1 0 12830 0 1 10810
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert203
timestamp 0
transform -1 0 12610 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert204
timestamp 0
transform -1 0 12510 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert205
timestamp 0
transform 1 0 12050 0 1 5530
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert206
timestamp 0
transform 1 0 14030 0 1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert207
timestamp 0
transform -1 0 11830 0 1 5530
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert208
timestamp 0
transform 1 0 15490 0 1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert209
timestamp 0
transform 1 0 150 0 1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert210
timestamp 0
transform 1 0 1130 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert211
timestamp 0
transform 1 0 310 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert212
timestamp 0
transform -1 0 790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert213
timestamp 0
transform -1 0 50 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert214
timestamp 0
transform 1 0 6410 0 1 6970
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert215
timestamp 0
transform -1 0 5730 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert216
timestamp 0
transform -1 0 4810 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert217
timestamp 0
transform -1 0 3490 0 1 6970
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert218
timestamp 0
transform 1 0 6690 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert219
timestamp 0
transform -1 0 11570 0 1 5530
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert220
timestamp 0
transform 1 0 11750 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert221
timestamp 0
transform -1 0 12110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert222
timestamp 0
transform -1 0 9970 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert223
timestamp 0
transform 1 0 12290 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert224
timestamp 0
transform -1 0 8950 0 1 14170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert225
timestamp 0
transform 1 0 6950 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert226
timestamp 0
transform -1 0 10570 0 1 15610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert227
timestamp 0
transform -1 0 6850 0 1 15130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert228
timestamp 0
transform -1 0 7550 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert229
timestamp 0
transform 1 0 8970 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert230
timestamp 0
transform 1 0 8730 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert231
timestamp 0
transform -1 0 7450 0 1 16090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert232
timestamp 0
transform -1 0 8930 0 1 15130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert233
timestamp 0
transform -1 0 15150 0 1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert234
timestamp 0
transform 1 0 15370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert235
timestamp 0
transform -1 0 12930 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert236
timestamp 0
transform -1 0 12130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert237
timestamp 0
transform -1 0 13230 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert238
timestamp 0
transform -1 0 2290 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert239
timestamp 0
transform -1 0 4670 0 1 13210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert240
timestamp 0
transform 1 0 5210 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert241
timestamp 0
transform 1 0 5630 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert242
timestamp 0
transform 1 0 5410 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert243
timestamp 0
transform -1 0 1850 0 1 5530
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert244
timestamp 0
transform -1 0 1410 0 1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert245
timestamp 0
transform 1 0 4470 0 1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert246
timestamp 0
transform 1 0 2430 0 1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert247
timestamp 0
transform 1 0 3870 0 1 5530
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert248
timestamp 0
transform 1 0 2270 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert249
timestamp 0
transform 1 0 3250 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert250
timestamp 0
transform -1 0 450 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert251
timestamp 0
transform -1 0 1910 0 -1 15610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert252
timestamp 0
transform 1 0 3050 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert253
timestamp 0
transform 1 0 8630 0 1 6010
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert254
timestamp 0
transform 1 0 11370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert255
timestamp 0
transform -1 0 10230 0 1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert256
timestamp 0
transform 1 0 11110 0 1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert257
timestamp 0
transform 1 0 12050 0 1 6010
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert258
timestamp 0
transform -1 0 13990 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert259
timestamp 0
transform -1 0 13750 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert260
timestamp 0
transform 1 0 16470 0 1 15610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert261
timestamp 0
transform -1 0 15870 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert262
timestamp 0
transform -1 0 13450 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert263
timestamp 0
transform -1 0 13350 0 1 13690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert264
timestamp 0
transform 1 0 4550 0 1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert265
timestamp 0
transform 1 0 5430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert266
timestamp 0
transform -1 0 4290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert267
timestamp 0
transform -1 0 4410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert268
timestamp 0
transform -1 0 4370 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert269
timestamp 0
transform -1 0 7530 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert270
timestamp 0
transform -1 0 7190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert271
timestamp 0
transform 1 0 9850 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert272
timestamp 0
transform 1 0 8070 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert273
timestamp 0
transform 1 0 9010 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert274
timestamp 0
transform -1 0 8270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert275
timestamp 0
transform 1 0 9870 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert276
timestamp 0
transform 1 0 9690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert277
timestamp 0
transform -1 0 7030 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert278
timestamp 0
transform 1 0 7450 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert279
timestamp 0
transform 1 0 9910 0 1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert280
timestamp 0
transform -1 0 15930 0 1 14170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert281
timestamp 0
transform -1 0 15870 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert282
timestamp 0
transform 1 0 15910 0 1 13690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert283
timestamp 0
transform -1 0 16590 0 1 14170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert284
timestamp 0
transform 1 0 16090 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert285
timestamp 0
transform -1 0 15870 0 1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert286
timestamp 0
transform -1 0 16330 0 1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert287
timestamp 0
transform 1 0 16370 0 1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert288
timestamp 0
transform 1 0 15070 0 1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert289
timestamp 0
transform -1 0 13010 0 1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert290
timestamp 0
transform 1 0 6730 0 1 12730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert291
timestamp 0
transform 1 0 6590 0 1 12730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert292
timestamp 0
transform -1 0 6490 0 1 12730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert293
timestamp 0
transform 1 0 8290 0 1 12730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert294
timestamp 0
transform -1 0 11870 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert295
timestamp 0
transform -1 0 11890 0 1 10330
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert296
timestamp 0
transform 1 0 15230 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert297
timestamp 0
transform 1 0 15010 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert298
timestamp 0
transform 1 0 17070 0 1 10330
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert299
timestamp 0
transform 1 0 16910 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert300
timestamp 0
transform 1 0 9110 0 1 14650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert301
timestamp 0
transform -1 0 7990 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert302
timestamp 0
transform -1 0 8070 0 1 14650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert303
timestamp 0
transform -1 0 8050 0 1 12730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert304
timestamp 0
transform -1 0 8570 0 1 6970
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert305
timestamp 0
transform 1 0 8610 0 1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert306
timestamp 0
transform -1 0 9690 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert307
timestamp 0
transform 1 0 9710 0 1 6970
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert308
timestamp 0
transform 1 0 10210 0 1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert309
timestamp 0
transform -1 0 13650 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert310
timestamp 0
transform 1 0 13750 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert311
timestamp 0
transform -1 0 15910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert312
timestamp 0
transform -1 0 15990 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert313
timestamp 0
transform -1 0 15090 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert314
timestamp 0
transform 1 0 15610 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert315
timestamp 0
transform 1 0 16390 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert316
timestamp 0
transform 1 0 14250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert317
timestamp 0
transform 1 0 16370 0 1 5530
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert318
timestamp 0
transform -1 0 11690 0 1 5530
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert319
timestamp 0
transform 1 0 11930 0 1 5530
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert320
timestamp 0
transform 1 0 8570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert321
timestamp 0
transform -1 0 6950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert322
timestamp 0
transform 1 0 7030 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert323
timestamp 0
transform 1 0 8650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert324
timestamp 0
transform -1 0 650 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert325
timestamp 0
transform 1 0 2970 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert326
timestamp 0
transform 1 0 2090 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert327
timestamp 0
transform -1 0 2890 0 1 15130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert328
timestamp 0
transform 1 0 1050 0 1 15610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert329
timestamp 0
transform 1 0 2070 0 1 16570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert330
timestamp 0
transform -1 0 2850 0 1 15610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert331
timestamp 0
transform 1 0 3750 0 1 14170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert332
timestamp 0
transform -1 0 2830 0 1 12730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert333
timestamp 0
transform -1 0 1810 0 1 15130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert334
timestamp 0
transform 1 0 2810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert335
timestamp 0
transform 1 0 2570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert336
timestamp 0
transform 1 0 310 0 1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert337
timestamp 0
transform -1 0 1170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert338
timestamp 0
transform -1 0 1530 0 1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert339
timestamp 0
transform -1 0 810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert340
timestamp 0
transform 1 0 310 0 1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert341
timestamp 0
transform -1 0 550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert342
timestamp 0
transform 1 0 1190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert343
timestamp 0
transform 1 0 190 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert344
timestamp 0
transform -1 0 50 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert345
timestamp 0
transform 1 0 10870 0 -1 16570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert346
timestamp 0
transform -1 0 11070 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert347
timestamp 0
transform 1 0 11490 0 1 15130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert348
timestamp 0
transform -1 0 10930 0 1 13690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert349
timestamp 0
transform 1 0 8090 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert350
timestamp 0
transform -1 0 7810 0 -1 16090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert351
timestamp 0
transform -1 0 7630 0 1 15130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert352
timestamp 0
transform 1 0 7750 0 1 15130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert353
timestamp 0
transform 1 0 10730 0 -1 14650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert354
timestamp 0
transform -1 0 6470 0 1 16090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert355
timestamp 0
transform -1 0 9450 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert356
timestamp 0
transform 1 0 9450 0 1 16090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert357
timestamp 0
transform -1 0 7050 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert358
timestamp 0
transform 1 0 10770 0 1 13690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert359
timestamp 0
transform -1 0 9470 0 1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert360
timestamp 0
transform -1 0 7510 0 1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert361
timestamp 0
transform -1 0 6310 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert362
timestamp 0
transform -1 0 8170 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert363
timestamp 0
transform 1 0 6670 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert364
timestamp 0
transform 1 0 3470 0 1 11770
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert365
timestamp 0
transform -1 0 4810 0 1 13210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert366
timestamp 0
transform -1 0 3670 0 1 13210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert367
timestamp 0
transform -1 0 2970 0 -1 13210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert368
timestamp 0
transform -1 0 4750 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert369
timestamp 0
transform 1 0 13330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert370
timestamp 0
transform -1 0 12910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert371
timestamp 0
transform 1 0 12030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert372
timestamp 0
transform 1 0 13190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert373
timestamp 0
transform -1 0 11190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert374
timestamp 0
transform 1 0 2870 0 1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert375
timestamp 0
transform 1 0 2990 0 1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert376
timestamp 0
transform -1 0 1450 0 1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert377
timestamp 0
transform -1 0 1990 0 1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert378
timestamp 0
transform -1 0 1330 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert379
timestamp 0
transform 1 0 6350 0 1 11770
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert380
timestamp 0
transform 1 0 4930 0 1 13210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert381
timestamp 0
transform -1 0 2870 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert382
timestamp 0
transform 1 0 5750 0 1 11290
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert383
timestamp 0
transform -1 0 4510 0 1 11290
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert29
timestamp 0
transform -1 0 9410 0 1 4570
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert30
timestamp 0
transform 1 0 10470 0 1 16570
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert31
timestamp 0
transform -1 0 1750 0 1 5050
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert32
timestamp 0
transform -1 0 6210 0 1 12250
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert33
timestamp 0
transform -1 0 5790 0 -1 14170
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert34
timestamp 0
transform -1 0 10050 0 1 7450
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert35
timestamp 0
transform -1 0 13190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert36
timestamp 0
transform 1 0 3510 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert37
timestamp 0
transform -1 0 14690 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert38
timestamp 0
transform 1 0 5630 0 1 10810
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert39
timestamp 0
transform -1 0 5870 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert40
timestamp 0
transform 1 0 15890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert41
timestamp 0
transform -1 0 11310 0 1 3130
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert42
timestamp 0
transform 1 0 9470 0 1 11290
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert43
timestamp 0
transform 1 0 7370 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert44
timestamp 0
transform 1 0 2750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert45
timestamp 0
transform 1 0 11050 0 -1 15130
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert46
timestamp 0
transform 1 0 3490 0 1 6490
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert47
timestamp 0
transform 1 0 12990 0 1 7930
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert48
timestamp 0
transform -1 0 2090 0 -1 12730
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert49
timestamp 0
transform 1 0 6110 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert50
timestamp 0
transform -1 0 13490 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert51
timestamp 0
transform 1 0 14710 0 1 13690
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert52
timestamp 0
transform -1 0 7030 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert53
timestamp 0
transform -1 0 4250 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert54
timestamp 0
transform 1 0 13110 0 1 6970
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert55
timestamp 0
transform 1 0 14150 0 1 12730
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert56
timestamp 0
transform -1 0 11190 0 1 7930
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert57
timestamp 0
transform -1 0 14690 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert58
timestamp 0
transform 1 0 7150 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert59
timestamp 0
transform -1 0 5850 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert60
timestamp 0
transform -1 0 8850 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert61
timestamp 0
transform 1 0 6350 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert62
timestamp 0
transform 1 0 11190 0 1 7450
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert63
timestamp 0
transform 1 0 10330 0 1 12250
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert64
timestamp 0
transform 1 0 3790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert65
timestamp 0
transform 1 0 6930 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert66
timestamp 0
transform 1 0 10570 0 1 16090
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert67
timestamp 0
transform -1 0 15210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert68
timestamp 0
transform -1 0 6250 0 1 14170
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert69
timestamp 0
transform 1 0 6930 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert70
timestamp 0
transform 1 0 3030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert71
timestamp 0
transform -1 0 2610 0 1 11770
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert72
timestamp 0
transform 1 0 9410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert73
timestamp 0
transform 1 0 12390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert74
timestamp 0
transform 1 0 15290 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert75
timestamp 0
transform 1 0 10330 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert76
timestamp 0
transform 1 0 8310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert77
timestamp 0
transform 1 0 11410 0 1 7930
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert78
timestamp 0
transform 1 0 10830 0 1 15610
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert79
timestamp 0
transform 1 0 11370 0 1 4570
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert80
timestamp 0
transform 1 0 4510 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert81
timestamp 0
transform -1 0 5330 0 1 13210
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert82
timestamp 0
transform 1 0 11950 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert83
timestamp 0
transform -1 0 1810 0 1 6490
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert84
timestamp 0
transform 1 0 8450 0 1 11290
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert85
timestamp 0
transform -1 0 5290 0 -1 13690
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert86
timestamp 0
transform 1 0 12590 0 1 3130
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert87
timestamp 0
transform -1 0 12050 0 1 7450
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert88
timestamp 0
transform 1 0 8070 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert89
timestamp 0
transform 1 0 6510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert90
timestamp 0
transform -1 0 2790 0 1 13210
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert91
timestamp 0
transform -1 0 2130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert92
timestamp 0
transform 1 0 9370 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert93
timestamp 0
transform -1 0 2130 0 1 7450
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert94
timestamp 0
transform -1 0 4110 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert95
timestamp 0
transform -1 0 3090 0 1 11770
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert96
timestamp 0
transform -1 0 8990 0 1 5050
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert97
timestamp 0
transform -1 0 9250 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert98
timestamp 0
transform -1 0 8110 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert99
timestamp 0
transform -1 0 9910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert100
timestamp 0
transform 1 0 11630 0 1 4570
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert101
timestamp 0
transform -1 0 14930 0 -1 12250
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert102
timestamp 0
transform 1 0 12270 0 1 7450
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert103
timestamp 0
transform -1 0 10130 0 1 6970
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert104
timestamp 0
transform -1 0 6190 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert105
timestamp 0
transform -1 0 6590 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert106
timestamp 0
transform -1 0 2190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert107
timestamp 0
transform 1 0 9710 0 1 11290
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert384
timestamp 0
transform 1 0 8910 0 -1 17050
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert385
timestamp 0
transform -1 0 5570 0 1 6490
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert386
timestamp 0
transform -1 0 4670 0 1 5050
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert387
timestamp 0
transform 1 0 10770 0 1 7450
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert388
timestamp 0
transform -1 0 7850 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert389
timestamp 0
transform 1 0 8370 0 1 6010
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert390
timestamp 0
transform -1 0 10350 0 1 4570
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert391
timestamp 0
transform -1 0 7030 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__7072_
timestamp 0
transform 1 0 6170 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__7074_
timestamp 0
transform 1 0 6710 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__7076_
timestamp 0
transform -1 0 5850 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__7079_
timestamp 0
transform -1 0 6810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__7081_
timestamp 0
transform -1 0 5430 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__7084_
timestamp 0
transform 1 0 8690 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__7086_
timestamp 0
transform -1 0 5630 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__7088_
timestamp 0
transform -1 0 5210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__7091_
timestamp 0
transform -1 0 5450 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__7093_
timestamp 0
transform -1 0 5270 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__7096_
timestamp 0
transform -1 0 5710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__7098_
timestamp 0
transform -1 0 5830 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__7100_
timestamp 0
transform 1 0 5470 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__7103_
timestamp 0
transform 1 0 6410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__7105_
timestamp 0
transform 1 0 5350 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__7107_
timestamp 0
transform 1 0 4910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__7110_
timestamp 0
transform -1 0 5370 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__7112_
timestamp 0
transform -1 0 6250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__7115_
timestamp 0
transform -1 0 8990 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__7117_
timestamp 0
transform -1 0 10810 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__7119_
timestamp 0
transform 1 0 8670 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__7122_
timestamp 0
transform -1 0 7910 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__7124_
timestamp 0
transform 1 0 9130 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__7127_
timestamp 0
transform 1 0 9110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__7129_
timestamp 0
transform -1 0 8970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__7131_
timestamp 0
transform 1 0 8490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__7134_
timestamp 0
transform 1 0 13070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7136_
timestamp 0
transform 1 0 13130 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7138_
timestamp 0
transform -1 0 10490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7141_
timestamp 0
transform -1 0 9310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__7143_
timestamp 0
transform -1 0 9150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__7146_
timestamp 0
transform 1 0 9570 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7148_
timestamp 0
transform -1 0 10010 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7150_
timestamp 0
transform 1 0 8910 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7153_
timestamp 0
transform 1 0 9750 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__7155_
timestamp 0
transform 1 0 7970 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__7158_
timestamp 0
transform -1 0 6490 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__7160_
timestamp 0
transform -1 0 10190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7162_
timestamp 0
transform 1 0 9210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7165_
timestamp 0
transform 1 0 8670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__7167_
timestamp 0
transform -1 0 9210 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7169_
timestamp 0
transform 1 0 8830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__7172_
timestamp 0
transform 1 0 11150 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7174_
timestamp 0
transform -1 0 9890 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7177_
timestamp 0
transform 1 0 8350 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__7179_
timestamp 0
transform 1 0 10350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7181_
timestamp 0
transform 1 0 9150 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7184_
timestamp 0
transform -1 0 9010 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7186_
timestamp 0
transform 1 0 8530 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7188_
timestamp 0
transform -1 0 8010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__7191_
timestamp 0
transform 1 0 10350 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7193_
timestamp 0
transform -1 0 10190 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7196_
timestamp 0
transform -1 0 7970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__7198_
timestamp 0
transform 1 0 8110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__7200_
timestamp 0
transform 1 0 8470 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7203_
timestamp 0
transform -1 0 6630 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__7205_
timestamp 0
transform 1 0 9410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__7208_
timestamp 0
transform -1 0 7810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__7210_
timestamp 0
transform -1 0 8910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7212_
timestamp 0
transform -1 0 9410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7215_
timestamp 0
transform 1 0 8910 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7217_
timestamp 0
transform 1 0 9190 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7219_
timestamp 0
transform 1 0 9310 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7222_
timestamp 0
transform -1 0 8370 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7224_
timestamp 0
transform -1 0 7710 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7227_
timestamp 0
transform -1 0 7450 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7229_
timestamp 0
transform -1 0 6150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__7231_
timestamp 0
transform -1 0 5930 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__7234_
timestamp 0
transform 1 0 8370 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7236_
timestamp 0
transform -1 0 8750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7239_
timestamp 0
transform -1 0 9470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__7241_
timestamp 0
transform 1 0 7650 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__7243_
timestamp 0
transform -1 0 8110 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__7246_
timestamp 0
transform -1 0 6490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__7248_
timestamp 0
transform 1 0 6530 0 1 730
box -6 -8 26 248
use FILL  FILL_2__7250_
timestamp 0
transform -1 0 6190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__7253_
timestamp 0
transform 1 0 6430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__7255_
timestamp 0
transform -1 0 8090 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7258_
timestamp 0
transform -1 0 5790 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__7260_
timestamp 0
transform -1 0 7950 0 1 730
box -6 -8 26 248
use FILL  FILL_2__7262_
timestamp 0
transform -1 0 8250 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7265_
timestamp 0
transform -1 0 6690 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__7267_
timestamp 0
transform -1 0 5690 0 1 250
box -6 -8 26 248
use FILL  FILL_2__7270_
timestamp 0
transform -1 0 5190 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__7272_
timestamp 0
transform -1 0 5490 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__7274_
timestamp 0
transform 1 0 5610 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__7277_
timestamp 0
transform 1 0 5830 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__7279_
timestamp 0
transform 1 0 6130 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__7281_
timestamp 0
transform -1 0 6250 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__7284_
timestamp 0
transform -1 0 7370 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__7286_
timestamp 0
transform 1 0 6790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__7289_
timestamp 0
transform -1 0 5570 0 1 250
box -6 -8 26 248
use FILL  FILL_2__7291_
timestamp 0
transform -1 0 5810 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__7293_
timestamp 0
transform 1 0 5970 0 1 730
box -6 -8 26 248
use FILL  FILL_2__7296_
timestamp 0
transform 1 0 7910 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7298_
timestamp 0
transform 1 0 6070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__7300_
timestamp 0
transform -1 0 4290 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__7303_
timestamp 0
transform 1 0 7090 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__7305_
timestamp 0
transform -1 0 4830 0 1 250
box -6 -8 26 248
use FILL  FILL_2__7308_
timestamp 0
transform -1 0 4150 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__7310_
timestamp 0
transform -1 0 4670 0 1 250
box -6 -8 26 248
use FILL  FILL_2__7312_
timestamp 0
transform -1 0 4510 0 1 250
box -6 -8 26 248
use FILL  FILL_2__7315_
timestamp 0
transform 1 0 5510 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__7317_
timestamp 0
transform -1 0 5370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__7320_
timestamp 0
transform 1 0 5510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__7322_
timestamp 0
transform -1 0 3850 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__7324_
timestamp 0
transform -1 0 5910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__7327_
timestamp 0
transform -1 0 4770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__7329_
timestamp 0
transform 1 0 5190 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__7331_
timestamp 0
transform -1 0 7290 0 1 730
box -6 -8 26 248
use FILL  FILL_2__7334_
timestamp 0
transform -1 0 6250 0 1 730
box -6 -8 26 248
use FILL  FILL_2__7336_
timestamp 0
transform -1 0 4990 0 1 250
box -6 -8 26 248
use FILL  FILL_2__7339_
timestamp 0
transform 1 0 5350 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__7341_
timestamp 0
transform 1 0 5410 0 1 730
box -6 -8 26 248
use FILL  FILL_2__7343_
timestamp 0
transform -1 0 5030 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__7346_
timestamp 0
transform 1 0 5150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__7348_
timestamp 0
transform 1 0 5330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__7351_
timestamp 0
transform 1 0 6170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__7353_
timestamp 0
transform -1 0 5290 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__7355_
timestamp 0
transform -1 0 5450 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7358_
timestamp 0
transform -1 0 5850 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7360_
timestamp 0
transform -1 0 5730 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7362_
timestamp 0
transform 1 0 5550 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7365_
timestamp 0
transform 1 0 6130 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7367_
timestamp 0
transform -1 0 6850 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7370_
timestamp 0
transform -1 0 6010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__7372_
timestamp 0
transform -1 0 4930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__7374_
timestamp 0
transform 1 0 5130 0 1 730
box -6 -8 26 248
use FILL  FILL_2__7377_
timestamp 0
transform -1 0 6690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7379_
timestamp 0
transform 1 0 6090 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__7382_
timestamp 0
transform 1 0 6450 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7384_
timestamp 0
transform 1 0 6610 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7386_
timestamp 0
transform 1 0 6290 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7389_
timestamp 0
transform -1 0 7230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7391_
timestamp 0
transform -1 0 6510 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7393_
timestamp 0
transform -1 0 5090 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__7396_
timestamp 0
transform -1 0 7090 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7398_
timestamp 0
transform 1 0 6770 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7401_
timestamp 0
transform -1 0 7330 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7403_
timestamp 0
transform 1 0 7590 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7405_
timestamp 0
transform 1 0 8190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7408_
timestamp 0
transform 1 0 7650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7410_
timestamp 0
transform 1 0 7210 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7412_
timestamp 0
transform 1 0 6970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__7415_
timestamp 0
transform 1 0 7130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__7417_
timestamp 0
transform 1 0 5950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__7420_
timestamp 0
transform 1 0 7450 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__7422_
timestamp 0
transform 1 0 7670 0 1 250
box -6 -8 26 248
use FILL  FILL_2__7424_
timestamp 0
transform -1 0 7690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__7427_
timestamp 0
transform -1 0 7310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__7429_
timestamp 0
transform -1 0 6830 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7432_
timestamp 0
transform -1 0 6670 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7434_
timestamp 0
transform 1 0 8230 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__7436_
timestamp 0
transform -1 0 7230 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__7439_
timestamp 0
transform 1 0 8050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__7441_
timestamp 0
transform -1 0 7730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__7443_
timestamp 0
transform 1 0 5270 0 1 250
box -6 -8 26 248
use FILL  FILL_2__7446_
timestamp 0
transform 1 0 6390 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__7448_
timestamp 0
transform 1 0 8250 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__7451_
timestamp 0
transform -1 0 8090 0 1 250
box -6 -8 26 248
use FILL  FILL_2__7453_
timestamp 0
transform 1 0 8210 0 1 250
box -6 -8 26 248
use FILL  FILL_2__7455_
timestamp 0
transform -1 0 10070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__7458_
timestamp 0
transform 1 0 10370 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7460_
timestamp 0
transform -1 0 6650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__7463_
timestamp 0
transform 1 0 8070 0 1 730
box -6 -8 26 248
use FILL  FILL_2__7465_
timestamp 0
transform 1 0 6890 0 1 730
box -6 -8 26 248
use FILL  FILL_2__7467_
timestamp 0
transform 1 0 8510 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__7470_
timestamp 0
transform -1 0 8250 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__7472_
timestamp 0
transform -1 0 8730 0 1 730
box -6 -8 26 248
use FILL  FILL_2__7474_
timestamp 0
transform -1 0 8270 0 1 730
box -6 -8 26 248
use FILL  FILL_2__7477_
timestamp 0
transform 1 0 9590 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7479_
timestamp 0
transform 1 0 9430 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7482_
timestamp 0
transform -1 0 10010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__7484_
timestamp 0
transform -1 0 8650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__7486_
timestamp 0
transform 1 0 11190 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7489_
timestamp 0
transform -1 0 7790 0 1 730
box -6 -8 26 248
use FILL  FILL_2__7491_
timestamp 0
transform 1 0 8350 0 1 250
box -6 -8 26 248
use FILL  FILL_2__7494_
timestamp 0
transform -1 0 7830 0 1 250
box -6 -8 26 248
use FILL  FILL_2__7496_
timestamp 0
transform -1 0 9090 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__7498_
timestamp 0
transform 1 0 8870 0 1 730
box -6 -8 26 248
use FILL  FILL_2__7501_
timestamp 0
transform -1 0 11670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7503_
timestamp 0
transform 1 0 11630 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7505_
timestamp 0
transform 1 0 11490 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7508_
timestamp 0
transform 1 0 11770 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7510_
timestamp 0
transform -1 0 7730 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__7513_
timestamp 0
transform 1 0 9050 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__7515_
timestamp 0
transform -1 0 7970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__7517_
timestamp 0
transform 1 0 9190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__7520_
timestamp 0
transform 1 0 9350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__7522_
timestamp 0
transform 1 0 12130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7524_
timestamp 0
transform 1 0 12250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7527_
timestamp 0
transform 1 0 12590 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7529_
timestamp 0
transform -1 0 11950 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7532_
timestamp 0
transform -1 0 7990 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__7534_
timestamp 0
transform 1 0 8770 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__7536_
timestamp 0
transform -1 0 10810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__7539_
timestamp 0
transform 1 0 11690 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7541_
timestamp 0
transform -1 0 11170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__7544_
timestamp 0
transform 1 0 11310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__7546_
timestamp 0
transform 1 0 12650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__7548_
timestamp 0
transform 1 0 12650 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7551_
timestamp 0
transform -1 0 9710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__7553_
timestamp 0
transform 1 0 11110 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__7555_
timestamp 0
transform 1 0 8790 0 1 250
box -6 -8 26 248
use FILL  FILL_2__7558_
timestamp 0
transform 1 0 10430 0 1 730
box -6 -8 26 248
use FILL  FILL_2__7560_
timestamp 0
transform 1 0 9290 0 1 730
box -6 -8 26 248
use FILL  FILL_2__7563_
timestamp 0
transform -1 0 10310 0 1 730
box -6 -8 26 248
use FILL  FILL_2__7565_
timestamp 0
transform 1 0 13710 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7567_
timestamp 0
transform 1 0 13570 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7570_
timestamp 0
transform -1 0 11590 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__7572_
timestamp 0
transform 1 0 9130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__7575_
timestamp 0
transform 1 0 9490 0 1 250
box -6 -8 26 248
use FILL  FILL_2__7577_
timestamp 0
transform 1 0 10370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__7579_
timestamp 0
transform -1 0 9650 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__7582_
timestamp 0
transform -1 0 13010 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7584_
timestamp 0
transform -1 0 12030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__7586_
timestamp 0
transform -1 0 12670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7589_
timestamp 0
transform 1 0 12090 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7591_
timestamp 0
transform 1 0 13970 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7594_
timestamp 0
transform 1 0 13410 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7596_
timestamp 0
transform -1 0 10770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__7598_
timestamp 0
transform 1 0 9250 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__7601_
timestamp 0
transform -1 0 9670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__7603_
timestamp 0
transform 1 0 9210 0 1 250
box -6 -8 26 248
use FILL  FILL_2__7606_
timestamp 0
transform 1 0 10030 0 1 730
box -6 -8 26 248
use FILL  FILL_2__7608_
timestamp 0
transform 1 0 10090 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__7610_
timestamp 0
transform 1 0 9930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__7613_
timestamp 0
transform 1 0 11410 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7615_
timestamp 0
transform 1 0 11150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__7617_
timestamp 0
transform -1 0 10890 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__7620_
timestamp 0
transform 1 0 12230 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7622_
timestamp 0
transform 1 0 11910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7625_
timestamp 0
transform 1 0 9330 0 1 250
box -6 -8 26 248
use FILL  FILL_2__7627_
timestamp 0
transform 1 0 10330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__7629_
timestamp 0
transform 1 0 11550 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7632_
timestamp 0
transform 1 0 10730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__7634_
timestamp 0
transform 1 0 11930 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7637_
timestamp 0
transform -1 0 11350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__7639_
timestamp 0
transform -1 0 10290 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__7641_
timestamp 0
transform 1 0 11490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__7644_
timestamp 0
transform -1 0 10050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__7646_
timestamp 0
transform 1 0 10990 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7648_
timestamp 0
transform 1 0 12850 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__7651_
timestamp 0
transform -1 0 11050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__7653_
timestamp 0
transform -1 0 10430 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__7656_
timestamp 0
transform -1 0 11650 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7658_
timestamp 0
transform 1 0 11330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__7660_
timestamp 0
transform 1 0 9470 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__7663_
timestamp 0
transform 1 0 9670 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__7665_
timestamp 0
transform 1 0 10430 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__7667_
timestamp 0
transform -1 0 9630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__7670_
timestamp 0
transform 1 0 10790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__7672_
timestamp 0
transform 1 0 10890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__7675_
timestamp 0
transform 1 0 9970 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__7677_
timestamp 0
transform 1 0 11130 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7679_
timestamp 0
transform 1 0 10270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__7682_
timestamp 0
transform -1 0 10610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__7684_
timestamp 0
transform -1 0 10130 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__7687_
timestamp 0
transform -1 0 6290 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__7689_
timestamp 0
transform -1 0 6150 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__7691_
timestamp 0
transform -1 0 5730 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__7694_
timestamp 0
transform -1 0 5510 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__7696_
timestamp 0
transform -1 0 6090 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__7698_
timestamp 0
transform -1 0 6390 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__7701_
timestamp 0
transform -1 0 5830 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__7703_
timestamp 0
transform -1 0 5690 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__7706_
timestamp 0
transform -1 0 5310 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__7708_
timestamp 0
transform -1 0 6070 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__7710_
timestamp 0
transform 1 0 7230 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__7713_
timestamp 0
transform 1 0 7630 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__7715_
timestamp 0
transform 1 0 7350 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__7718_
timestamp 0
transform -1 0 6810 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__7720_
timestamp 0
transform 1 0 6290 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__7722_
timestamp 0
transform -1 0 6950 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__7725_
timestamp 0
transform -1 0 7710 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__7727_
timestamp 0
transform 1 0 7070 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__7729_
timestamp 0
transform -1 0 6550 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__7732_
timestamp 0
transform -1 0 6370 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__7734_
timestamp 0
transform -1 0 6290 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__7737_
timestamp 0
transform -1 0 8110 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__7739_
timestamp 0
transform 1 0 7190 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__7741_
timestamp 0
transform 1 0 7710 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__7744_
timestamp 0
transform -1 0 6570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__7746_
timestamp 0
transform 1 0 7130 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__7749_
timestamp 0
transform -1 0 8150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__7751_
timestamp 0
transform 1 0 8850 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__7753_
timestamp 0
transform 1 0 8290 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__7756_
timestamp 0
transform -1 0 8030 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__7758_
timestamp 0
transform 1 0 7470 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__7760_
timestamp 0
transform 1 0 7170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__7763_
timestamp 0
transform -1 0 7510 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__7765_
timestamp 0
transform 1 0 7850 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__7768_
timestamp 0
transform 1 0 7890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__7770_
timestamp 0
transform 1 0 7850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__7772_
timestamp 0
transform -1 0 7730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__7775_
timestamp 0
transform 1 0 6930 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__7777_
timestamp 0
transform 1 0 7350 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__7779_
timestamp 0
transform 1 0 7090 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__7782_
timestamp 0
transform 1 0 6650 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__7784_
timestamp 0
transform -1 0 4910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__7787_
timestamp 0
transform -1 0 5170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__7789_
timestamp 0
transform 1 0 5290 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__7791_
timestamp 0
transform -1 0 6090 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__7794_
timestamp 0
transform -1 0 8490 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__7796_
timestamp 0
transform 1 0 7110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__7799_
timestamp 0
transform -1 0 7250 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__7801_
timestamp 0
transform -1 0 6510 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__7803_
timestamp 0
transform -1 0 6930 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__7806_
timestamp 0
transform -1 0 7450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__7808_
timestamp 0
transform 1 0 8210 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__7810_
timestamp 0
transform -1 0 7070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__7813_
timestamp 0
transform 1 0 7890 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__7815_
timestamp 0
transform -1 0 6410 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__7818_
timestamp 0
transform 1 0 7470 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__7820_
timestamp 0
transform 1 0 7630 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__7822_
timestamp 0
transform 1 0 7070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__7825_
timestamp 0
transform -1 0 6350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__7827_
timestamp 0
transform 1 0 6170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__7830_
timestamp 0
transform 1 0 6330 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__7832_
timestamp 0
transform 1 0 6770 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__7834_
timestamp 0
transform 1 0 6910 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__7837_
timestamp 0
transform 1 0 6910 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__7839_
timestamp 0
transform -1 0 10530 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7841_
timestamp 0
transform 1 0 9610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__7844_
timestamp 0
transform 1 0 9290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__7846_
timestamp 0
transform -1 0 6670 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__7849_
timestamp 0
transform 1 0 9770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__7851_
timestamp 0
transform -1 0 6170 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__7853_
timestamp 0
transform 1 0 10990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__7856_
timestamp 0
transform 1 0 8930 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__7858_
timestamp 0
transform -1 0 8790 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__7861_
timestamp 0
transform -1 0 9130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__7863_
timestamp 0
transform 1 0 10090 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__7865_
timestamp 0
transform -1 0 7090 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__7868_
timestamp 0
transform -1 0 6810 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__7870_
timestamp 0
transform -1 0 7070 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__7872_
timestamp 0
transform -1 0 7950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__7875_
timestamp 0
transform -1 0 6650 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__7877_
timestamp 0
transform -1 0 6830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__7880_
timestamp 0
transform -1 0 6090 0 1 250
box -6 -8 26 248
use FILL  FILL_2__7882_
timestamp 0
transform -1 0 7190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__7884_
timestamp 0
transform -1 0 7230 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__7887_
timestamp 0
transform 1 0 8210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__7889_
timestamp 0
transform -1 0 7470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__7891_
timestamp 0
transform 1 0 7190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__7894_
timestamp 0
transform 1 0 8350 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__7896_
timestamp 0
transform -1 0 8230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__7899_
timestamp 0
transform 1 0 7530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__7901_
timestamp 0
transform -1 0 8090 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__7903_
timestamp 0
transform -1 0 4930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__7906_
timestamp 0
transform 1 0 8850 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__7908_
timestamp 0
transform -1 0 8310 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__7911_
timestamp 0
transform -1 0 6950 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__7913_
timestamp 0
transform 1 0 6790 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__7915_
timestamp 0
transform 1 0 6170 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__7998_
timestamp 0
transform -1 0 4950 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8000_
timestamp 0
transform 1 0 4350 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__8002_
timestamp 0
transform -1 0 4510 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__8005_
timestamp 0
transform -1 0 4370 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__8007_
timestamp 0
transform 1 0 4490 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__8010_
timestamp 0
transform -1 0 3790 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__8012_
timestamp 0
transform -1 0 4030 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__8014_
timestamp 0
transform 1 0 6570 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__8017_
timestamp 0
transform 1 0 4870 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__8019_
timestamp 0
transform -1 0 4510 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__8022_
timestamp 0
transform -1 0 4250 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8024_
timestamp 0
transform 1 0 2990 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__8026_
timestamp 0
transform -1 0 3570 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__8029_
timestamp 0
transform 1 0 3370 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__8031_
timestamp 0
transform -1 0 3670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__8033_
timestamp 0
transform 1 0 3130 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__8036_
timestamp 0
transform -1 0 4370 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__8038_
timestamp 0
transform 1 0 3090 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__8041_
timestamp 0
transform 1 0 4450 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8043_
timestamp 0
transform 1 0 4530 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8045_
timestamp 0
transform 1 0 3930 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8048_
timestamp 0
transform -1 0 3570 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__8050_
timestamp 0
transform 1 0 4570 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8053_
timestamp 0
transform 1 0 2910 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__8055_
timestamp 0
transform -1 0 5410 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8057_
timestamp 0
transform 1 0 1570 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__8060_
timestamp 0
transform 1 0 2490 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__8062_
timestamp 0
transform -1 0 3950 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__8064_
timestamp 0
transform 1 0 3610 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__8067_
timestamp 0
transform -1 0 4030 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__8069_
timestamp 0
transform -1 0 2950 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__8072_
timestamp 0
transform 1 0 3810 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8074_
timestamp 0
transform 1 0 5250 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8076_
timestamp 0
transform 1 0 5570 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__8079_
timestamp 0
transform -1 0 4990 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8081_
timestamp 0
transform 1 0 6850 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8084_
timestamp 0
transform -1 0 2890 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8086_
timestamp 0
transform -1 0 2630 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8088_
timestamp 0
transform 1 0 3670 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8091_
timestamp 0
transform 1 0 3150 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__8093_
timestamp 0
transform -1 0 3370 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8095_
timestamp 0
transform -1 0 70 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__8098_
timestamp 0
transform -1 0 2730 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8100_
timestamp 0
transform 1 0 3370 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__8103_
timestamp 0
transform -1 0 3230 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8105_
timestamp 0
transform 1 0 3190 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8107_
timestamp 0
transform -1 0 2250 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__8110_
timestamp 0
transform -1 0 3650 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8112_
timestamp 0
transform -1 0 2150 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__8114_
timestamp 0
transform 1 0 2150 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8117_
timestamp 0
transform -1 0 3350 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8119_
timestamp 0
transform 1 0 4830 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8122_
timestamp 0
transform -1 0 4950 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8124_
timestamp 0
transform -1 0 4830 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8126_
timestamp 0
transform -1 0 4530 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8129_
timestamp 0
transform 1 0 7210 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__8131_
timestamp 0
transform 1 0 4510 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__8134_
timestamp 0
transform -1 0 1990 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8136_
timestamp 0
transform -1 0 4090 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8138_
timestamp 0
transform 1 0 4370 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8141_
timestamp 0
transform -1 0 4290 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8143_
timestamp 0
transform 1 0 4390 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8145_
timestamp 0
transform -1 0 4830 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__8148_
timestamp 0
transform 1 0 5290 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8150_
timestamp 0
transform 1 0 4890 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8153_
timestamp 0
transform 1 0 3930 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8155_
timestamp 0
transform 1 0 3570 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__8157_
timestamp 0
transform -1 0 4650 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8160_
timestamp 0
transform -1 0 4550 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8162_
timestamp 0
transform -1 0 1570 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__8165_
timestamp 0
transform 1 0 1570 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__8167_
timestamp 0
transform 1 0 5970 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__8169_
timestamp 0
transform 1 0 1590 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8172_
timestamp 0
transform 1 0 1010 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__8174_
timestamp 0
transform 1 0 1990 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__8176_
timestamp 0
transform 1 0 2370 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__8179_
timestamp 0
transform -1 0 2830 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__8181_
timestamp 0
transform -1 0 2310 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__8184_
timestamp 0
transform -1 0 450 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__8186_
timestamp 0
transform -1 0 1750 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__8188_
timestamp 0
transform 1 0 1670 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8191_
timestamp 0
transform 1 0 810 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__8193_
timestamp 0
transform -1 0 870 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__8196_
timestamp 0
transform 1 0 570 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__8198_
timestamp 0
transform 1 0 710 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__8200_
timestamp 0
transform 1 0 1130 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__8203_
timestamp 0
transform -1 0 990 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__8205_
timestamp 0
transform -1 0 490 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__8207_
timestamp 0
transform 1 0 1030 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__8210_
timestamp 0
transform 1 0 550 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8212_
timestamp 0
transform -1 0 690 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__8215_
timestamp 0
transform 1 0 50 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__8217_
timestamp 0
transform 1 0 190 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__8219_
timestamp 0
transform 1 0 1130 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__8222_
timestamp 0
transform -1 0 2510 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__8224_
timestamp 0
transform 1 0 510 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8226_
timestamp 0
transform -1 0 630 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__8229_
timestamp 0
transform -1 0 70 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8231_
timestamp 0
transform -1 0 330 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__8234_
timestamp 0
transform -1 0 70 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__8236_
timestamp 0
transform 1 0 510 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__8238_
timestamp 0
transform -1 0 590 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__8241_
timestamp 0
transform 1 0 530 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__8243_
timestamp 0
transform 1 0 1210 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8246_
timestamp 0
transform -1 0 230 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8248_
timestamp 0
transform 1 0 210 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__8250_
timestamp 0
transform -1 0 390 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__8253_
timestamp 0
transform -1 0 230 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__8255_
timestamp 0
transform -1 0 810 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__8257_
timestamp 0
transform -1 0 870 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__8260_
timestamp 0
transform 1 0 170 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__8262_
timestamp 0
transform 1 0 530 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8265_
timestamp 0
transform 1 0 190 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8267_
timestamp 0
transform -1 0 830 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8269_
timestamp 0
transform -1 0 870 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__8272_
timestamp 0
transform -1 0 2190 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8274_
timestamp 0
transform -1 0 2670 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8277_
timestamp 0
transform -1 0 1030 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__8279_
timestamp 0
transform -1 0 410 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__8281_
timestamp 0
transform -1 0 570 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__8284_
timestamp 0
transform -1 0 70 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__8286_
timestamp 0
transform -1 0 250 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__8288_
timestamp 0
transform 1 0 330 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__8291_
timestamp 0
transform 1 0 1050 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8293_
timestamp 0
transform 1 0 1550 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8296_
timestamp 0
transform 1 0 350 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8298_
timestamp 0
transform -1 0 670 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8300_
timestamp 0
transform 1 0 630 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__8303_
timestamp 0
transform 1 0 170 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__8305_
timestamp 0
transform 1 0 750 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__8308_
timestamp 0
transform -1 0 310 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8310_
timestamp 0
transform 1 0 150 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8312_
timestamp 0
transform 1 0 450 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8315_
timestamp 0
transform 1 0 1290 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__8317_
timestamp 0
transform -1 0 3230 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__8319_
timestamp 0
transform 1 0 450 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__8322_
timestamp 0
transform 1 0 330 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__8324_
timestamp 0
transform -1 0 610 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__8327_
timestamp 0
transform -1 0 70 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8329_
timestamp 0
transform -1 0 70 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__8331_
timestamp 0
transform -1 0 570 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8334_
timestamp 0
transform 1 0 730 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__8336_
timestamp 0
transform 1 0 690 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8338_
timestamp 0
transform 1 0 890 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8341_
timestamp 0
transform -1 0 2910 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8343_
timestamp 0
transform -1 0 590 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__8346_
timestamp 0
transform 1 0 550 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__8348_
timestamp 0
transform -1 0 190 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__8350_
timestamp 0
transform -1 0 70 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__8353_
timestamp 0
transform 1 0 790 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__8355_
timestamp 0
transform 1 0 1270 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8358_
timestamp 0
transform 1 0 3390 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8360_
timestamp 0
transform -1 0 4330 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__8362_
timestamp 0
transform 1 0 4130 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8365_
timestamp 0
transform 1 0 5710 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8367_
timestamp 0
transform 1 0 770 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8369_
timestamp 0
transform 1 0 1270 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__8372_
timestamp 0
transform -1 0 1750 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8374_
timestamp 0
transform -1 0 2710 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__8377_
timestamp 0
transform -1 0 1050 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8379_
timestamp 0
transform 1 0 2870 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__8381_
timestamp 0
transform -1 0 2790 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__8384_
timestamp 0
transform -1 0 1850 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__8386_
timestamp 0
transform -1 0 5510 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__8389_
timestamp 0
transform -1 0 330 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__8391_
timestamp 0
transform 1 0 850 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8393_
timestamp 0
transform -1 0 1050 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__8396_
timestamp 0
transform 1 0 1750 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8398_
timestamp 0
transform 1 0 1230 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8400_
timestamp 0
transform -1 0 2630 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__8403_
timestamp 0
transform -1 0 2410 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__8405_
timestamp 0
transform -1 0 2410 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8408_
timestamp 0
transform -1 0 2630 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__8410_
timestamp 0
transform -1 0 2370 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__8412_
timestamp 0
transform -1 0 1030 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__8415_
timestamp 0
transform -1 0 1430 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__8417_
timestamp 0
transform 1 0 1450 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8420_
timestamp 0
transform 1 0 2050 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8422_
timestamp 0
transform 1 0 2170 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8424_
timestamp 0
transform -1 0 2330 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__8427_
timestamp 0
transform -1 0 2130 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__8429_
timestamp 0
transform -1 0 2090 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__8431_
timestamp 0
transform 1 0 3410 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8434_
timestamp 0
transform -1 0 890 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8436_
timestamp 0
transform 1 0 910 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__8439_
timestamp 0
transform 1 0 1690 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__8441_
timestamp 0
transform -1 0 1970 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__8443_
timestamp 0
transform 1 0 2250 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__8446_
timestamp 0
transform -1 0 2610 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8448_
timestamp 0
transform -1 0 2470 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8450_
timestamp 0
transform 1 0 1850 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__8453_
timestamp 0
transform 1 0 2690 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__8455_
timestamp 0
transform 1 0 1150 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__8458_
timestamp 0
transform 1 0 1710 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__8460_
timestamp 0
transform 1 0 2190 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__8462_
timestamp 0
transform -1 0 1890 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8465_
timestamp 0
transform 1 0 2450 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8467_
timestamp 0
transform 1 0 2150 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8470_
timestamp 0
transform 1 0 3430 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8472_
timestamp 0
transform -1 0 4130 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8474_
timestamp 0
transform -1 0 4290 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8477_
timestamp 0
transform -1 0 2330 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__8479_
timestamp 0
transform 1 0 1290 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__8481_
timestamp 0
transform -1 0 1450 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8484_
timestamp 0
transform 1 0 1910 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8486_
timestamp 0
transform -1 0 1590 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__8489_
timestamp 0
transform 1 0 3450 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__8491_
timestamp 0
transform 1 0 3570 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__8493_
timestamp 0
transform 1 0 4110 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__8496_
timestamp 0
transform -1 0 4250 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__8498_
timestamp 0
transform 1 0 1330 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__8501_
timestamp 0
transform 1 0 2230 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__8503_
timestamp 0
transform -1 0 1590 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__8505_
timestamp 0
transform -1 0 2410 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__8508_
timestamp 0
transform -1 0 3070 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__8510_
timestamp 0
transform -1 0 2890 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__8512_
timestamp 0
transform 1 0 3710 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__8515_
timestamp 0
transform 1 0 3270 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8517_
timestamp 0
transform 1 0 3010 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__8520_
timestamp 0
transform 1 0 3570 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__8522_
timestamp 0
transform -1 0 4090 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__8524_
timestamp 0
transform -1 0 2790 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__8527_
timestamp 0
transform 1 0 1230 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8529_
timestamp 0
transform 1 0 1230 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__8532_
timestamp 0
transform -1 0 1530 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__8534_
timestamp 0
transform 1 0 1790 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__8536_
timestamp 0
transform -1 0 1970 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__8539_
timestamp 0
transform 1 0 3030 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__8541_
timestamp 0
transform 1 0 3830 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__8543_
timestamp 0
transform -1 0 2250 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__8546_
timestamp 0
transform -1 0 2170 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8548_
timestamp 0
transform -1 0 1650 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__8551_
timestamp 0
transform 1 0 1710 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8553_
timestamp 0
transform 1 0 1870 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8555_
timestamp 0
transform 1 0 1750 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__8558_
timestamp 0
transform 1 0 2030 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__8560_
timestamp 0
transform 1 0 1870 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__8563_
timestamp 0
transform 1 0 3030 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__8565_
timestamp 0
transform 1 0 2290 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__8567_
timestamp 0
transform 1 0 1710 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8570_
timestamp 0
transform 1 0 1950 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8572_
timestamp 0
transform 1 0 2110 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8574_
timestamp 0
transform -1 0 2230 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__8577_
timestamp 0
transform 1 0 2630 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__8579_
timestamp 0
transform -1 0 2110 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__8582_
timestamp 0
transform -1 0 1990 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__8584_
timestamp 0
transform -1 0 1370 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8586_
timestamp 0
transform -1 0 1610 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__8589_
timestamp 0
transform 1 0 1590 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__8591_
timestamp 0
transform -1 0 1070 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__8593_
timestamp 0
transform 1 0 1210 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__8596_
timestamp 0
transform 1 0 1890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__8598_
timestamp 0
transform -1 0 3710 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__8601_
timestamp 0
transform -1 0 1610 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__8603_
timestamp 0
transform 1 0 430 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__8605_
timestamp 0
transform 1 0 290 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__8608_
timestamp 0
transform 1 0 2430 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__8610_
timestamp 0
transform -1 0 6050 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8613_
timestamp 0
transform 1 0 5730 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8615_
timestamp 0
transform -1 0 4630 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__8617_
timestamp 0
transform 1 0 6630 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8620_
timestamp 0
transform 1 0 6650 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__8622_
timestamp 0
transform 1 0 6190 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8624_
timestamp 0
transform -1 0 6150 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8627_
timestamp 0
transform 1 0 6330 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__8629_
timestamp 0
transform 1 0 6250 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__8632_
timestamp 0
transform -1 0 6090 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__8634_
timestamp 0
transform 1 0 5270 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__8636_
timestamp 0
transform 1 0 5390 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__8639_
timestamp 0
transform -1 0 5210 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__8641_
timestamp 0
transform -1 0 6610 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8644_
timestamp 0
transform 1 0 6570 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__8646_
timestamp 0
transform 1 0 6450 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8648_
timestamp 0
transform 1 0 5810 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8651_
timestamp 0
transform 1 0 6070 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8653_
timestamp 0
transform 1 0 6050 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8655_
timestamp 0
transform -1 0 6210 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8658_
timestamp 0
transform -1 0 5890 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8660_
timestamp 0
transform -1 0 7270 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__8663_
timestamp 0
transform 1 0 6610 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8665_
timestamp 0
transform 1 0 6970 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8667_
timestamp 0
transform -1 0 6810 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__8670_
timestamp 0
transform 1 0 7190 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8672_
timestamp 0
transform 1 0 7370 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8675_
timestamp 0
transform -1 0 6270 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__8677_
timestamp 0
transform 1 0 6130 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8679_
timestamp 0
transform -1 0 7350 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8682_
timestamp 0
transform 1 0 6770 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8684_
timestamp 0
transform -1 0 7590 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8686_
timestamp 0
transform -1 0 6930 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8689_
timestamp 0
transform 1 0 7130 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8691_
timestamp 0
transform 1 0 6870 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__8694_
timestamp 0
transform -1 0 5910 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__8696_
timestamp 0
transform 1 0 6030 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__8698_
timestamp 0
transform 1 0 6170 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__8701_
timestamp 0
transform 1 0 6410 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__8703_
timestamp 0
transform 1 0 7110 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8705_
timestamp 0
transform 1 0 6210 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__8708_
timestamp 0
transform 1 0 6650 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8710_
timestamp 0
transform 1 0 6930 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8713_
timestamp 0
transform 1 0 7190 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8715_
timestamp 0
transform 1 0 7410 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8717_
timestamp 0
transform 1 0 6430 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__8720_
timestamp 0
transform 1 0 6590 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8722_
timestamp 0
transform 1 0 5710 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__8725_
timestamp 0
transform 1 0 6510 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__8727_
timestamp 0
transform -1 0 6690 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__8729_
timestamp 0
transform -1 0 6590 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__8732_
timestamp 0
transform -1 0 6190 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__8734_
timestamp 0
transform -1 0 5570 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__8736_
timestamp 0
transform 1 0 6030 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__8739_
timestamp 0
transform -1 0 5450 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__8741_
timestamp 0
transform -1 0 4850 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__8744_
timestamp 0
transform -1 0 6330 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__8746_
timestamp 0
transform 1 0 5270 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__8748_
timestamp 0
transform 1 0 5390 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__8751_
timestamp 0
transform 1 0 5250 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__8753_
timestamp 0
transform 1 0 4310 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__8756_
timestamp 0
transform 1 0 4090 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__8758_
timestamp 0
transform -1 0 4070 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__8760_
timestamp 0
transform 1 0 1050 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__8763_
timestamp 0
transform 1 0 4290 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8765_
timestamp 0
transform -1 0 4010 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8767_
timestamp 0
transform -1 0 4990 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__8770_
timestamp 0
transform 1 0 5230 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8772_
timestamp 0
transform -1 0 3570 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__8775_
timestamp 0
transform 1 0 5370 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__8777_
timestamp 0
transform 1 0 3810 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8779_
timestamp 0
transform -1 0 2810 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8782_
timestamp 0
transform -1 0 5250 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__8784_
timestamp 0
transform 1 0 3290 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__8787_
timestamp 0
transform 1 0 2990 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__8789_
timestamp 0
transform 1 0 1150 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__8791_
timestamp 0
transform 1 0 1310 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__8794_
timestamp 0
transform -1 0 4810 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8796_
timestamp 0
transform -1 0 3850 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8798_
timestamp 0
transform 1 0 5270 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__8801_
timestamp 0
transform -1 0 3590 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__8803_
timestamp 0
transform 1 0 2210 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__8806_
timestamp 0
transform 1 0 4190 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__8808_
timestamp 0
transform -1 0 4050 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__8810_
timestamp 0
transform 1 0 5650 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__8813_
timestamp 0
transform 1 0 5430 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__8815_
timestamp 0
transform -1 0 4770 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__8817_
timestamp 0
transform 1 0 5150 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__8820_
timestamp 0
transform 1 0 5450 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__8822_
timestamp 0
transform 1 0 5670 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__8825_
timestamp 0
transform 1 0 5330 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__8827_
timestamp 0
transform 1 0 6270 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__8829_
timestamp 0
transform -1 0 6710 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8832_
timestamp 0
transform 1 0 4750 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__8834_
timestamp 0
transform 1 0 5510 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__8837_
timestamp 0
transform -1 0 5490 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__8839_
timestamp 0
transform -1 0 5850 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__8921_
timestamp 0
transform -1 0 2830 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__8924_
timestamp 0
transform -1 0 4070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__8926_
timestamp 0
transform -1 0 4310 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__8928_
timestamp 0
transform 1 0 4550 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__8931_
timestamp 0
transform 1 0 4190 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__8933_
timestamp 0
transform 1 0 4010 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__8936_
timestamp 0
transform 1 0 4330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__8938_
timestamp 0
transform 1 0 4910 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__8940_
timestamp 0
transform -1 0 4950 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__8943_
timestamp 0
transform 1 0 4650 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__8945_
timestamp 0
transform 1 0 5610 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__8948_
timestamp 0
transform -1 0 6050 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__8950_
timestamp 0
transform -1 0 5390 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__8952_
timestamp 0
transform 1 0 4770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__8955_
timestamp 0
transform 1 0 5590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__8957_
timestamp 0
transform -1 0 4950 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__8959_
timestamp 0
transform -1 0 5130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__8962_
timestamp 0
transform 1 0 3590 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__8964_
timestamp 0
transform 1 0 4530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__8967_
timestamp 0
transform -1 0 5550 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__8969_
timestamp 0
transform -1 0 4010 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__8971_
timestamp 0
transform 1 0 5970 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__8974_
timestamp 0
transform 1 0 4230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__8976_
timestamp 0
transform 1 0 4170 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__8979_
timestamp 0
transform -1 0 2410 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__8981_
timestamp 0
transform -1 0 310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__8983_
timestamp 0
transform -1 0 1250 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__8986_
timestamp 0
transform -1 0 930 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__8988_
timestamp 0
transform -1 0 1210 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__8990_
timestamp 0
transform -1 0 670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__8993_
timestamp 0
transform 1 0 1450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__8995_
timestamp 0
transform 1 0 1070 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__8998_
timestamp 0
transform -1 0 2270 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__9000_
timestamp 0
transform -1 0 470 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__9002_
timestamp 0
transform 1 0 3450 0 1 250
box -6 -8 26 248
use FILL  FILL_2__9005_
timestamp 0
transform 1 0 4530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__9007_
timestamp 0
transform -1 0 3610 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__9009_
timestamp 0
transform -1 0 590 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__9012_
timestamp 0
transform -1 0 210 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__9014_
timestamp 0
transform -1 0 630 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__9017_
timestamp 0
transform 1 0 470 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__9019_
timestamp 0
transform -1 0 170 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__9021_
timestamp 0
transform -1 0 830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__9024_
timestamp 0
transform -1 0 1270 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9026_
timestamp 0
transform 1 0 1070 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9029_
timestamp 0
transform -1 0 1530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9031_
timestamp 0
transform 1 0 1710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__9033_
timestamp 0
transform 1 0 1490 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__9036_
timestamp 0
transform 1 0 750 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9038_
timestamp 0
transform -1 0 790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9040_
timestamp 0
transform -1 0 1050 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__9043_
timestamp 0
transform -1 0 1710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__9045_
timestamp 0
transform 1 0 1850 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__9048_
timestamp 0
transform 1 0 2670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__9050_
timestamp 0
transform 1 0 2970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__9052_
timestamp 0
transform 1 0 7530 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__9055_
timestamp 0
transform -1 0 3990 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__9057_
timestamp 0
transform -1 0 470 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9060_
timestamp 0
transform -1 0 330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__9062_
timestamp 0
transform 1 0 590 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__9064_
timestamp 0
transform 1 0 2130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__9067_
timestamp 0
transform 1 0 1970 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__9069_
timestamp 0
transform 1 0 2270 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__9071_
timestamp 0
transform 1 0 3550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__9074_
timestamp 0
transform -1 0 3410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__9076_
timestamp 0
transform 1 0 4030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9079_
timestamp 0
transform 1 0 4870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__9081_
timestamp 0
transform 1 0 3130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__9083_
timestamp 0
transform -1 0 2950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__9086_
timestamp 0
transform -1 0 350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__9088_
timestamp 0
transform -1 0 950 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9091_
timestamp 0
transform 1 0 1550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__9093_
timestamp 0
transform 1 0 1570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__9095_
timestamp 0
transform -1 0 2690 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__9098_
timestamp 0
transform 1 0 3190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__9100_
timestamp 0
transform 1 0 3510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__9102_
timestamp 0
transform 1 0 4090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__9105_
timestamp 0
transform 1 0 3350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__9107_
timestamp 0
transform -1 0 230 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9110_
timestamp 0
transform 1 0 650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__9112_
timestamp 0
transform -1 0 970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9114_
timestamp 0
transform 1 0 3350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9117_
timestamp 0
transform -1 0 2970 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9119_
timestamp 0
transform 1 0 3950 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9122_
timestamp 0
transform 1 0 3730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9124_
timestamp 0
transform 1 0 4930 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9126_
timestamp 0
transform -1 0 5850 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9129_
timestamp 0
transform 1 0 2950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9131_
timestamp 0
transform 1 0 570 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9133_
timestamp 0
transform -1 0 1090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__9136_
timestamp 0
transform -1 0 3130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9138_
timestamp 0
transform -1 0 2830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__9141_
timestamp 0
transform -1 0 3550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__9143_
timestamp 0
transform 1 0 4430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9145_
timestamp 0
transform 1 0 4730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9148_
timestamp 0
transform 1 0 4530 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9150_
timestamp 0
transform 1 0 690 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9152_
timestamp 0
transform -1 0 870 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9155_
timestamp 0
transform 1 0 2790 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9157_
timestamp 0
transform 1 0 4930 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9160_
timestamp 0
transform 1 0 3810 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9162_
timestamp 0
transform 1 0 3790 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9164_
timestamp 0
transform -1 0 4790 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9167_
timestamp 0
transform 1 0 5310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9169_
timestamp 0
transform 1 0 5050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9172_
timestamp 0
transform -1 0 4090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__9174_
timestamp 0
transform -1 0 3930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__9176_
timestamp 0
transform -1 0 4210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9179_
timestamp 0
transform -1 0 430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9181_
timestamp 0
transform -1 0 1510 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9183_
timestamp 0
transform -1 0 3390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9186_
timestamp 0
transform 1 0 4030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9188_
timestamp 0
transform 1 0 3770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9191_
timestamp 0
transform 1 0 4270 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__9193_
timestamp 0
transform 1 0 4890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9195_
timestamp 0
transform 1 0 4330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__9198_
timestamp 0
transform -1 0 4910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9200_
timestamp 0
transform -1 0 3750 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__9203_
timestamp 0
transform -1 0 2390 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__9205_
timestamp 0
transform 1 0 1170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9207_
timestamp 0
transform 1 0 2890 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__9210_
timestamp 0
transform 1 0 2490 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__9212_
timestamp 0
transform 1 0 3030 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__9214_
timestamp 0
transform 1 0 4210 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__9217_
timestamp 0
transform 1 0 4630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__9219_
timestamp 0
transform -1 0 4330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9222_
timestamp 0
transform 1 0 4730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9224_
timestamp 0
transform -1 0 4110 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__9226_
timestamp 0
transform -1 0 3670 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__9229_
timestamp 0
transform 1 0 1330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9231_
timestamp 0
transform 1 0 3150 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__9234_
timestamp 0
transform 1 0 3770 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__9236_
timestamp 0
transform 1 0 3930 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__9238_
timestamp 0
transform 1 0 4470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__9241_
timestamp 0
transform -1 0 5190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9243_
timestamp 0
transform 1 0 910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9245_
timestamp 0
transform 1 0 3670 0 1 730
box -6 -8 26 248
use FILL  FILL_2__9248_
timestamp 0
transform -1 0 3310 0 1 730
box -6 -8 26 248
use FILL  FILL_2__9250_
timestamp 0
transform 1 0 3750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__9253_
timestamp 0
transform -1 0 3990 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__9255_
timestamp 0
transform -1 0 4130 0 1 730
box -6 -8 26 248
use FILL  FILL_2__9257_
timestamp 0
transform -1 0 3910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__9260_
timestamp 0
transform 1 0 4250 0 1 730
box -6 -8 26 248
use FILL  FILL_2__9262_
timestamp 0
transform 1 0 4550 0 1 730
box -6 -8 26 248
use FILL  FILL_2__9264_
timestamp 0
transform 1 0 4850 0 1 730
box -6 -8 26 248
use FILL  FILL_2__9267_
timestamp 0
transform -1 0 4230 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__9269_
timestamp 0
transform 1 0 290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9272_
timestamp 0
transform -1 0 3590 0 1 250
box -6 -8 26 248
use FILL  FILL_2__9274_
timestamp 0
transform 1 0 3950 0 1 250
box -6 -8 26 248
use FILL  FILL_2__9276_
timestamp 0
transform -1 0 4230 0 1 250
box -6 -8 26 248
use FILL  FILL_2__9279_
timestamp 0
transform 1 0 4330 0 1 250
box -6 -8 26 248
use FILL  FILL_2__9281_
timestamp 0
transform -1 0 6110 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9284_
timestamp 0
transform 1 0 2910 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__9286_
timestamp 0
transform 1 0 1990 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__9288_
timestamp 0
transform -1 0 570 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__9291_
timestamp 0
transform -1 0 4270 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9293_
timestamp 0
transform -1 0 2390 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9295_
timestamp 0
transform -1 0 2390 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9298_
timestamp 0
transform 1 0 1830 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__9300_
timestamp 0
transform 1 0 2790 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9303_
timestamp 0
transform 1 0 2330 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__9305_
timestamp 0
transform -1 0 3870 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__9307_
timestamp 0
transform 1 0 3270 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__9310_
timestamp 0
transform 1 0 1290 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__9312_
timestamp 0
transform 1 0 1870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__9315_
timestamp 0
transform 1 0 1290 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9317_
timestamp 0
transform -1 0 2450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__9319_
timestamp 0
transform 1 0 1410 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9322_
timestamp 0
transform -1 0 2210 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9324_
timestamp 0
transform -1 0 2230 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9326_
timestamp 0
transform 1 0 2390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__9329_
timestamp 0
transform -1 0 2650 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__9331_
timestamp 0
transform 1 0 3050 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__9334_
timestamp 0
transform 1 0 2510 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__9336_
timestamp 0
transform 1 0 2130 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__9338_
timestamp 0
transform 1 0 2390 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__9341_
timestamp 0
transform -1 0 1830 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9343_
timestamp 0
transform 1 0 1710 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__9346_
timestamp 0
transform 1 0 2050 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9348_
timestamp 0
transform 1 0 2290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9350_
timestamp 0
transform 1 0 2450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9353_
timestamp 0
transform -1 0 3390 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9355_
timestamp 0
transform 1 0 3910 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__9357_
timestamp 0
transform -1 0 2550 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__9360_
timestamp 0
transform -1 0 1110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__9362_
timestamp 0
transform 1 0 2070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9365_
timestamp 0
transform 1 0 1390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__9367_
timestamp 0
transform 1 0 1950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__9369_
timestamp 0
transform 1 0 2250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__9372_
timestamp 0
transform 1 0 2650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__9374_
timestamp 0
transform -1 0 3210 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__9376_
timestamp 0
transform -1 0 5490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9379_
timestamp 0
transform -1 0 850 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__9381_
timestamp 0
transform -1 0 1570 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__9384_
timestamp 0
transform 1 0 1870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__9386_
timestamp 0
transform -1 0 1730 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__9388_
timestamp 0
transform -1 0 1590 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__9391_
timestamp 0
transform 1 0 1990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__9393_
timestamp 0
transform 1 0 2030 0 1 730
box -6 -8 26 248
use FILL  FILL_2__9396_
timestamp 0
transform 1 0 2570 0 1 730
box -6 -8 26 248
use FILL  FILL_2__9398_
timestamp 0
transform -1 0 5670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__9400_
timestamp 0
transform 1 0 2570 0 1 250
box -6 -8 26 248
use FILL  FILL_2__9403_
timestamp 0
transform -1 0 1010 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__9405_
timestamp 0
transform 1 0 1150 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__9407_
timestamp 0
transform 1 0 1930 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__9410_
timestamp 0
transform 1 0 1590 0 1 730
box -6 -8 26 248
use FILL  FILL_2__9412_
timestamp 0
transform -1 0 1870 0 1 250
box -6 -8 26 248
use FILL  FILL_2__9415_
timestamp 0
transform -1 0 2290 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__9417_
timestamp 0
transform 1 0 3150 0 1 250
box -6 -8 26 248
use FILL  FILL_2__9419_
timestamp 0
transform -1 0 3850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__9422_
timestamp 0
transform -1 0 690 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__9424_
timestamp 0
transform -1 0 1050 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__9427_
timestamp 0
transform 1 0 910 0 1 250
box -6 -8 26 248
use FILL  FILL_2__9429_
timestamp 0
transform -1 0 1330 0 1 250
box -6 -8 26 248
use FILL  FILL_2__9431_
timestamp 0
transform 1 0 1570 0 1 250
box -6 -8 26 248
use FILL  FILL_2__9434_
timestamp 0
transform 1 0 2290 0 1 250
box -6 -8 26 248
use FILL  FILL_2__9436_
timestamp 0
transform 1 0 2410 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__9438_
timestamp 0
transform 1 0 2730 0 1 250
box -6 -8 26 248
use FILL  FILL_2__9441_
timestamp 0
transform -1 0 1890 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__9443_
timestamp 0
transform 1 0 2890 0 1 250
box -6 -8 26 248
use FILL  FILL_2__9446_
timestamp 0
transform -1 0 5250 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9448_
timestamp 0
transform 1 0 2670 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__9450_
timestamp 0
transform -1 0 430 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__9453_
timestamp 0
transform -1 0 170 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__9455_
timestamp 0
transform -1 0 1030 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__9458_
timestamp 0
transform 1 0 310 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__9460_
timestamp 0
transform 1 0 850 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__9462_
timestamp 0
transform 1 0 2790 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__9465_
timestamp 0
transform 1 0 3170 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__9467_
timestamp 0
transform -1 0 1310 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__9469_
timestamp 0
transform -1 0 1470 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__9472_
timestamp 0
transform -1 0 1210 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__9474_
timestamp 0
transform 1 0 910 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__9477_
timestamp 0
transform 1 0 630 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__9479_
timestamp 0
transform 1 0 350 0 1 250
box -6 -8 26 248
use FILL  FILL_2__9481_
timestamp 0
transform 1 0 1150 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__9484_
timestamp 0
transform 1 0 2090 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__9486_
timestamp 0
transform -1 0 3190 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__9489_
timestamp 0
transform 1 0 2310 0 1 730
box -6 -8 26 248
use FILL  FILL_2__9491_
timestamp 0
transform -1 0 330 0 1 730
box -6 -8 26 248
use FILL  FILL_2__9493_
timestamp 0
transform -1 0 450 0 1 730
box -6 -8 26 248
use FILL  FILL_2__9496_
timestamp 0
transform -1 0 430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__9498_
timestamp 0
transform 1 0 1310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__9500_
timestamp 0
transform 1 0 2550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__9503_
timestamp 0
transform 1 0 950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__9505_
timestamp 0
transform 1 0 1310 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__9508_
timestamp 0
transform -1 0 350 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__9510_
timestamp 0
transform -1 0 210 0 1 250
box -6 -8 26 248
use FILL  FILL_2__9512_
timestamp 0
transform 1 0 350 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__9515_
timestamp 0
transform 1 0 190 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__9517_
timestamp 0
transform 1 0 170 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__9519_
timestamp 0
transform -1 0 70 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__9522_
timestamp 0
transform -1 0 4970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__9524_
timestamp 0
transform 1 0 50 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__9527_
timestamp 0
transform -1 0 2770 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__9529_
timestamp 0
transform -1 0 2910 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__9531_
timestamp 0
transform 1 0 2990 0 1 730
box -6 -8 26 248
use FILL  FILL_2__9534_
timestamp 0
transform 1 0 1430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9536_
timestamp 0
transform 1 0 1290 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9539_
timestamp 0
transform 1 0 3630 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9541_
timestamp 0
transform 1 0 2090 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9543_
timestamp 0
transform 1 0 1270 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__9546_
timestamp 0
transform 1 0 830 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9548_
timestamp 0
transform 1 0 870 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9550_
timestamp 0
transform -1 0 730 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9553_
timestamp 0
transform -1 0 1330 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9555_
timestamp 0
transform 1 0 1690 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9558_
timestamp 0
transform 1 0 170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__9560_
timestamp 0
transform -1 0 210 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__9562_
timestamp 0
transform -1 0 70 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9565_
timestamp 0
transform 1 0 270 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9567_
timestamp 0
transform -1 0 590 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9570_
timestamp 0
transform -1 0 190 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__9572_
timestamp 0
transform -1 0 930 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__9574_
timestamp 0
transform 1 0 470 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__9577_
timestamp 0
transform 1 0 650 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__9579_
timestamp 0
transform -1 0 730 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9581_
timestamp 0
transform -1 0 430 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__9584_
timestamp 0
transform 1 0 4350 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__9586_
timestamp 0
transform 1 0 990 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9589_
timestamp 0
transform 1 0 3190 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__9591_
timestamp 0
transform 1 0 3470 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__9593_
timestamp 0
transform 1 0 3870 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__9596_
timestamp 0
transform -1 0 3710 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9598_
timestamp 0
transform -1 0 1510 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__9601_
timestamp 0
transform 1 0 1530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__9603_
timestamp 0
transform -1 0 2770 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__9605_
timestamp 0
transform 1 0 3290 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__9608_
timestamp 0
transform -1 0 4690 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9610_
timestamp 0
transform -1 0 4490 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9612_
timestamp 0
transform -1 0 3870 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9615_
timestamp 0
transform 1 0 3990 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9617_
timestamp 0
transform 1 0 370 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__9620_
timestamp 0
transform -1 0 470 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9622_
timestamp 0
transform 1 0 2470 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9624_
timestamp 0
transform 1 0 3010 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9627_
timestamp 0
transform -1 0 4550 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9629_
timestamp 0
transform -1 0 4630 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9631_
timestamp 0
transform -1 0 2310 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__9634_
timestamp 0
transform -1 0 1690 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__9636_
timestamp 0
transform 1 0 2230 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9639_
timestamp 0
transform 1 0 4150 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__9641_
timestamp 0
transform -1 0 4310 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9643_
timestamp 0
transform -1 0 1370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__9646_
timestamp 0
transform 1 0 2830 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__9648_
timestamp 0
transform 1 0 2690 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__9651_
timestamp 0
transform 1 0 3130 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9653_
timestamp 0
transform -1 0 3310 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9655_
timestamp 0
transform -1 0 3290 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__9658_
timestamp 0
transform -1 0 2970 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__9660_
timestamp 0
transform -1 0 2010 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__9662_
timestamp 0
transform -1 0 2870 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__9665_
timestamp 0
transform -1 0 3650 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__9667_
timestamp 0
transform 1 0 2410 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__9670_
timestamp 0
transform 1 0 2690 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__9672_
timestamp 0
transform 1 0 2670 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__9674_
timestamp 0
transform 1 0 3190 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__9677_
timestamp 0
transform -1 0 4190 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__9679_
timestamp 0
transform 1 0 4010 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__9682_
timestamp 0
transform -1 0 2890 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__9684_
timestamp 0
transform -1 0 310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9686_
timestamp 0
transform -1 0 70 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__9689_
timestamp 0
transform 1 0 710 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__9691_
timestamp 0
transform -1 0 70 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__9693_
timestamp 0
transform -1 0 330 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__9696_
timestamp 0
transform -1 0 70 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__9698_
timestamp 0
transform -1 0 310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__9701_
timestamp 0
transform 1 0 1270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__9703_
timestamp 0
transform -1 0 1790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9705_
timestamp 0
transform 1 0 1010 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__9708_
timestamp 0
transform -1 0 1850 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__9710_
timestamp 0
transform -1 0 930 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__9713_
timestamp 0
transform -1 0 2950 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9715_
timestamp 0
transform -1 0 310 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9717_
timestamp 0
transform 1 0 2030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__9720_
timestamp 0
transform 1 0 3610 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__9722_
timestamp 0
transform 1 0 2350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__9724_
timestamp 0
transform -1 0 3050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__9727_
timestamp 0
transform -1 0 3430 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__9729_
timestamp 0
transform -1 0 2470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9732_
timestamp 0
transform -1 0 2850 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__9734_
timestamp 0
transform -1 0 2510 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__9736_
timestamp 0
transform -1 0 850 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__9739_
timestamp 0
transform -1 0 2530 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__9741_
timestamp 0
transform 1 0 1110 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__9743_
timestamp 0
transform 1 0 1670 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__9746_
timestamp 0
transform 1 0 2110 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__9748_
timestamp 0
transform -1 0 2330 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9751_
timestamp 0
transform 1 0 2450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9753_
timestamp 0
transform -1 0 2710 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__9755_
timestamp 0
transform 1 0 2970 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9758_
timestamp 0
transform -1 0 1050 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__9760_
timestamp 0
transform 1 0 1830 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__9763_
timestamp 0
transform -1 0 1010 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__9845_
timestamp 0
transform 1 0 9830 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__9847_
timestamp 0
transform 1 0 9950 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__9850_
timestamp 0
transform -1 0 10810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__9852_
timestamp 0
transform 1 0 10530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__9854_
timestamp 0
transform -1 0 10690 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__9857_
timestamp 0
transform 1 0 9870 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9859_
timestamp 0
transform 1 0 11690 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__9862_
timestamp 0
transform -1 0 10470 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__9864_
timestamp 0
transform -1 0 10410 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__9866_
timestamp 0
transform 1 0 9430 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__9869_
timestamp 0
transform -1 0 12610 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__9871_
timestamp 0
transform -1 0 13650 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9874_
timestamp 0
transform -1 0 12450 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9876_
timestamp 0
transform -1 0 12190 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__9878_
timestamp 0
transform -1 0 12930 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__9881_
timestamp 0
transform -1 0 12910 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__9883_
timestamp 0
transform -1 0 12770 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__9885_
timestamp 0
transform 1 0 12610 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__9888_
timestamp 0
transform -1 0 12190 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__9890_
timestamp 0
transform -1 0 11250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__9893_
timestamp 0
transform -1 0 10910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__9895_
timestamp 0
transform 1 0 11890 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__9897_
timestamp 0
transform -1 0 11730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__9900_
timestamp 0
transform 1 0 10450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__9902_
timestamp 0
transform -1 0 12530 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__9905_
timestamp 0
transform 1 0 15530 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__9907_
timestamp 0
transform -1 0 14770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__9909_
timestamp 0
transform -1 0 13370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__9912_
timestamp 0
transform -1 0 13990 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__9914_
timestamp 0
transform -1 0 13130 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__9916_
timestamp 0
transform -1 0 12590 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__9919_
timestamp 0
transform 1 0 13490 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__9921_
timestamp 0
transform 1 0 12570 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__9924_
timestamp 0
transform 1 0 12650 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__9926_
timestamp 0
transform -1 0 12390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__9928_
timestamp 0
transform 1 0 12710 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9931_
timestamp 0
transform -1 0 13930 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__9933_
timestamp 0
transform 1 0 13710 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__9935_
timestamp 0
transform -1 0 11610 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__9938_
timestamp 0
transform 1 0 12630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__9940_
timestamp 0
transform -1 0 12930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__9943_
timestamp 0
transform 1 0 14850 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__9945_
timestamp 0
transform -1 0 15950 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__9947_
timestamp 0
transform -1 0 13770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__9950_
timestamp 0
transform -1 0 14170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__9952_
timestamp 0
transform 1 0 13830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__9955_
timestamp 0
transform -1 0 13110 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__9957_
timestamp 0
transform -1 0 13550 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__9959_
timestamp 0
transform 1 0 13230 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__9962_
timestamp 0
transform -1 0 14670 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__9964_
timestamp 0
transform 1 0 14150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__9966_
timestamp 0
transform 1 0 14650 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__9969_
timestamp 0
transform -1 0 13630 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__9971_
timestamp 0
transform -1 0 13470 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__9974_
timestamp 0
transform 1 0 13310 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9976_
timestamp 0
transform 1 0 7730 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__9978_
timestamp 0
transform 1 0 7690 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__9981_
timestamp 0
transform -1 0 15370 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__9983_
timestamp 0
transform 1 0 14230 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__9986_
timestamp 0
transform -1 0 14590 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__9988_
timestamp 0
transform 1 0 14170 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__9990_
timestamp 0
transform 1 0 13390 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__9993_
timestamp 0
transform 1 0 14010 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__9995_
timestamp 0
transform -1 0 14170 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__9997_
timestamp 0
transform -1 0 13930 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10001_
timestamp 0
transform -1 0 13630 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10003_
timestamp 0
transform -1 0 13250 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__10005_
timestamp 0
transform 1 0 14450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10008_
timestamp 0
transform 1 0 14330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10010_
timestamp 0
transform 1 0 16450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__10013_
timestamp 0
transform -1 0 15730 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__10015_
timestamp 0
transform 1 0 14470 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10017_
timestamp 0
transform -1 0 15530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__10020_
timestamp 0
transform -1 0 14730 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__10022_
timestamp 0
transform -1 0 14730 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10025_
timestamp 0
transform -1 0 14270 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__10027_
timestamp 0
transform -1 0 13870 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__10029_
timestamp 0
transform 1 0 14490 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__10032_
timestamp 0
transform -1 0 15190 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__10034_
timestamp 0
transform -1 0 16050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__10036_
timestamp 0
transform -1 0 14710 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__10039_
timestamp 0
transform -1 0 14950 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10041_
timestamp 0
transform 1 0 15110 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__10044_
timestamp 0
transform -1 0 14650 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10046_
timestamp 0
transform 1 0 14770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10048_
timestamp 0
transform -1 0 14830 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10051_
timestamp 0
transform 1 0 14970 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10053_
timestamp 0
transform 1 0 14550 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__10056_
timestamp 0
transform 1 0 16010 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__10058_
timestamp 0
transform -1 0 15810 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__10060_
timestamp 0
transform 1 0 15330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10063_
timestamp 0
transform -1 0 15450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10065_
timestamp 0
transform 1 0 15330 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__10067_
timestamp 0
transform -1 0 14890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__10070_
timestamp 0
transform 1 0 13030 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__10072_
timestamp 0
transform -1 0 15610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10075_
timestamp 0
transform -1 0 15970 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__10077_
timestamp 0
transform 1 0 15690 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__10079_
timestamp 0
transform 1 0 15530 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__10082_
timestamp 0
transform 1 0 16070 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__10084_
timestamp 0
transform 1 0 16130 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10087_
timestamp 0
transform -1 0 15070 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__10089_
timestamp 0
transform -1 0 15150 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10091_
timestamp 0
transform -1 0 15150 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__10094_
timestamp 0
transform 1 0 15850 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10096_
timestamp 0
transform 1 0 15450 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__10098_
timestamp 0
transform 1 0 15610 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__10101_
timestamp 0
transform 1 0 15810 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10103_
timestamp 0
transform 1 0 16510 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__10106_
timestamp 0
transform -1 0 16310 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10108_
timestamp 0
transform 1 0 16230 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__10110_
timestamp 0
transform -1 0 16030 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10113_
timestamp 0
transform 1 0 15970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10115_
timestamp 0
transform -1 0 15530 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10117_
timestamp 0
transform 1 0 15570 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__10120_
timestamp 0
transform 1 0 13690 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__10122_
timestamp 0
transform 1 0 13530 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__10125_
timestamp 0
transform 1 0 15730 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__10127_
timestamp 0
transform 1 0 16510 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__10129_
timestamp 0
transform 1 0 16470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__10132_
timestamp 0
transform -1 0 16950 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10134_
timestamp 0
transform 1 0 16630 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__10137_
timestamp 0
transform -1 0 16870 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10139_
timestamp 0
transform -1 0 16470 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__10141_
timestamp 0
transform -1 0 16310 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__10144_
timestamp 0
transform -1 0 16050 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__10146_
timestamp 0
transform 1 0 16010 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10148_
timestamp 0
transform 1 0 16590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10151_
timestamp 0
transform 1 0 16450 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10153_
timestamp 0
transform 1 0 16630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__10156_
timestamp 0
transform 1 0 16790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__10158_
timestamp 0
transform 1 0 16250 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__10160_
timestamp 0
transform 1 0 16830 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10163_
timestamp 0
transform -1 0 16310 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10165_
timestamp 0
transform 1 0 13330 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10168_
timestamp 0
transform -1 0 17070 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__10170_
timestamp 0
transform -1 0 16910 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__10172_
timestamp 0
transform 1 0 16750 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__10175_
timestamp 0
transform -1 0 17110 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__10177_
timestamp 0
transform 1 0 16970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__10179_
timestamp 0
transform 1 0 17050 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__10182_
timestamp 0
transform 1 0 16470 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__10184_
timestamp 0
transform -1 0 17030 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10187_
timestamp 0
transform -1 0 16470 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10189_
timestamp 0
transform 1 0 14490 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10191_
timestamp 0
transform -1 0 16910 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10194_
timestamp 0
transform -1 0 16950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__10196_
timestamp 0
transform 1 0 16750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__10199_
timestamp 0
transform 1 0 16990 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__10201_
timestamp 0
transform -1 0 16890 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__10203_
timestamp 0
transform -1 0 16730 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__10206_
timestamp 0
transform -1 0 11590 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__10208_
timestamp 0
transform 1 0 14550 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__10210_
timestamp 0
transform 1 0 14170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__10213_
timestamp 0
transform -1 0 13070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10215_
timestamp 0
transform 1 0 15770 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10218_
timestamp 0
transform 1 0 15350 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__10220_
timestamp 0
transform 1 0 15390 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__10222_
timestamp 0
transform 1 0 12990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__10225_
timestamp 0
transform 1 0 15370 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__10227_
timestamp 0
transform 1 0 13250 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__10229_
timestamp 0
transform 1 0 10830 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__10232_
timestamp 0
transform 1 0 14710 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10234_
timestamp 0
transform -1 0 14330 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10237_
timestamp 0
transform -1 0 15830 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__10239_
timestamp 0
transform 1 0 15950 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__10241_
timestamp 0
transform 1 0 15630 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__10244_
timestamp 0
transform -1 0 15670 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__10246_
timestamp 0
transform -1 0 15570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__10249_
timestamp 0
transform -1 0 12790 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__10251_
timestamp 0
transform -1 0 12950 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__10253_
timestamp 0
transform 1 0 12690 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__10256_
timestamp 0
transform -1 0 10990 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__10258_
timestamp 0
transform 1 0 12610 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__10260_
timestamp 0
transform 1 0 16330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__10263_
timestamp 0
transform 1 0 16230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__10265_
timestamp 0
transform -1 0 14970 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__10268_
timestamp 0
transform -1 0 14550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__10270_
timestamp 0
transform 1 0 15090 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__10272_
timestamp 0
transform -1 0 13450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__10275_
timestamp 0
transform 1 0 13050 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__10277_
timestamp 0
transform 1 0 12230 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__10280_
timestamp 0
transform 1 0 12890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__10282_
timestamp 0
transform 1 0 16690 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__10284_
timestamp 0
transform 1 0 16070 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__10287_
timestamp 0
transform -1 0 14990 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__10289_
timestamp 0
transform 1 0 14790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__10291_
timestamp 0
transform -1 0 14130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__10294_
timestamp 0
transform -1 0 12810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__10296_
timestamp 0
transform -1 0 12670 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__10299_
timestamp 0
transform -1 0 12490 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__10301_
timestamp 0
transform 1 0 12910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__10303_
timestamp 0
transform 1 0 16790 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__10306_
timestamp 0
transform 1 0 15490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__10308_
timestamp 0
transform -1 0 15370 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__10311_
timestamp 0
transform -1 0 14530 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__10313_
timestamp 0
transform 1 0 15410 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__10315_
timestamp 0
transform -1 0 14690 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__10318_
timestamp 0
transform -1 0 13530 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__10320_
timestamp 0
transform -1 0 13390 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__10322_
timestamp 0
transform 1 0 12430 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__10325_
timestamp 0
transform 1 0 15830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__10327_
timestamp 0
transform 1 0 16150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__10330_
timestamp 0
transform -1 0 16130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__10332_
timestamp 0
transform 1 0 14950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__10334_
timestamp 0
transform 1 0 15690 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__10337_
timestamp 0
transform -1 0 14650 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__10339_
timestamp 0
transform -1 0 13950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__10341_
timestamp 0
transform -1 0 13530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__10344_
timestamp 0
transform 1 0 11370 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__10346_
timestamp 0
transform 1 0 16310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__10349_
timestamp 0
transform 1 0 15170 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__10351_
timestamp 0
transform 1 0 15610 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__10353_
timestamp 0
transform 1 0 15030 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__10356_
timestamp 0
transform -1 0 14510 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__10358_
timestamp 0
transform 1 0 14230 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__10361_
timestamp 0
transform -1 0 14250 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__10363_
timestamp 0
transform -1 0 13670 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__10365_
timestamp 0
transform 1 0 14470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__10368_
timestamp 0
transform -1 0 13870 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__10370_
timestamp 0
transform 1 0 11490 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__10372_
timestamp 0
transform -1 0 14030 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__10375_
timestamp 0
transform 1 0 16470 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__10377_
timestamp 0
transform -1 0 14870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__10380_
timestamp 0
transform -1 0 15030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__10382_
timestamp 0
transform 1 0 15510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__10384_
timestamp 0
transform -1 0 15650 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__10387_
timestamp 0
transform -1 0 13330 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__10389_
timestamp 0
transform -1 0 13070 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__10392_
timestamp 0
transform -1 0 14310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__10394_
timestamp 0
transform 1 0 16150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__10396_
timestamp 0
transform -1 0 16250 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__10399_
timestamp 0
transform -1 0 16570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__10401_
timestamp 0
transform -1 0 16290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__10403_
timestamp 0
transform -1 0 16730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__10406_
timestamp 0
transform -1 0 14150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__10408_
timestamp 0
transform -1 0 15370 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__10411_
timestamp 0
transform 1 0 12790 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__10413_
timestamp 0
transform -1 0 14010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__10415_
timestamp 0
transform 1 0 16930 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__10418_
timestamp 0
transform 1 0 15430 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__10420_
timestamp 0
transform 1 0 16950 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__10423_
timestamp 0
transform -1 0 13350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__10425_
timestamp 0
transform -1 0 13050 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__10427_
timestamp 0
transform 1 0 16830 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__10430_
timestamp 0
transform -1 0 16470 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__10432_
timestamp 0
transform -1 0 16350 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__10434_
timestamp 0
transform 1 0 16590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__10437_
timestamp 0
transform -1 0 16770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__10439_
timestamp 0
transform 1 0 17050 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__10442_
timestamp 0
transform 1 0 16530 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__10444_
timestamp 0
transform -1 0 15870 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__10446_
timestamp 0
transform 1 0 13190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__10449_
timestamp 0
transform 1 0 16130 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__10451_
timestamp 0
transform 1 0 16650 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__10453_
timestamp 0
transform 1 0 16510 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__10456_
timestamp 0
transform -1 0 12510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__10458_
timestamp 0
transform -1 0 9430 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__10461_
timestamp 0
transform 1 0 9570 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__10463_
timestamp 0
transform 1 0 9990 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__10465_
timestamp 0
transform 1 0 9290 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__10468_
timestamp 0
transform -1 0 9990 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10470_
timestamp 0
transform 1 0 9970 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__10473_
timestamp 0
transform -1 0 8670 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__10475_
timestamp 0
transform -1 0 8650 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10477_
timestamp 0
transform -1 0 8890 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10480_
timestamp 0
transform 1 0 8810 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__10482_
timestamp 0
transform -1 0 11130 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__10484_
timestamp 0
transform -1 0 10410 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__10487_
timestamp 0
transform 1 0 9090 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__10489_
timestamp 0
transform -1 0 8750 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__10492_
timestamp 0
transform 1 0 9590 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10494_
timestamp 0
transform 1 0 9890 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10496_
timestamp 0
transform 1 0 10270 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10499_
timestamp 0
transform 1 0 11030 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__10501_
timestamp 0
transform 1 0 10510 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10504_
timestamp 0
transform -1 0 9510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10506_
timestamp 0
transform 1 0 9330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10508_
timestamp 0
transform 1 0 11010 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__10511_
timestamp 0
transform 1 0 10730 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__10513_
timestamp 0
transform 1 0 10510 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10515_
timestamp 0
transform 1 0 10470 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__10518_
timestamp 0
transform 1 0 10990 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__10520_
timestamp 0
transform -1 0 10850 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__10523_
timestamp 0
transform 1 0 13150 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10525_
timestamp 0
transform -1 0 12890 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10527_
timestamp 0
transform -1 0 11110 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10530_
timestamp 0
transform 1 0 10990 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__10532_
timestamp 0
transform 1 0 10730 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__10535_
timestamp 0
transform 1 0 10610 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__10537_
timestamp 0
transform 1 0 10670 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10539_
timestamp 0
transform -1 0 10570 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__10542_
timestamp 0
transform -1 0 10530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10544_
timestamp 0
transform -1 0 10670 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10546_
timestamp 0
transform 1 0 10990 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10549_
timestamp 0
transform -1 0 9890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__10551_
timestamp 0
transform 1 0 9730 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__10554_
timestamp 0
transform -1 0 9850 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10556_
timestamp 0
transform 1 0 10730 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10558_
timestamp 0
transform -1 0 10470 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10561_
timestamp 0
transform 1 0 10310 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10563_
timestamp 0
transform -1 0 9550 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10566_
timestamp 0
transform 1 0 11150 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__10568_
timestamp 0
transform 1 0 11450 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__10570_
timestamp 0
transform -1 0 11150 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__10573_
timestamp 0
transform 1 0 10110 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10575_
timestamp 0
transform 1 0 10110 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__10577_
timestamp 0
transform -1 0 10290 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__10580_
timestamp 0
transform 1 0 11670 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__10582_
timestamp 0
transform 1 0 11390 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__10585_
timestamp 0
transform -1 0 11650 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10587_
timestamp 0
transform 1 0 11670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__10589_
timestamp 0
transform -1 0 11830 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__10592_
timestamp 0
transform -1 0 11270 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__10594_
timestamp 0
transform -1 0 11890 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__10596_
timestamp 0
transform 1 0 11910 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__10599_
timestamp 0
transform -1 0 12350 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__10601_
timestamp 0
transform -1 0 11970 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__10604_
timestamp 0
transform 1 0 10470 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__10606_
timestamp 0
transform 1 0 10610 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__10608_
timestamp 0
transform -1 0 16610 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__10611_
timestamp 0
transform 1 0 11590 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__10613_
timestamp 0
transform 1 0 11290 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__10616_
timestamp 0
transform 1 0 10890 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__10618_
timestamp 0
transform -1 0 10650 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__10620_
timestamp 0
transform 1 0 12610 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__10623_
timestamp 0
transform 1 0 10150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__10625_
timestamp 0
transform 1 0 13450 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__10627_
timestamp 0
transform -1 0 13870 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__10630_
timestamp 0
transform -1 0 12290 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__10632_
timestamp 0
transform 1 0 12470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__10635_
timestamp 0
transform 1 0 13530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__10637_
timestamp 0
transform -1 0 16450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__10639_
timestamp 0
transform -1 0 15890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__10642_
timestamp 0
transform 1 0 11950 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10644_
timestamp 0
transform 1 0 12390 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10647_
timestamp 0
transform 1 0 12010 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10649_
timestamp 0
transform 1 0 12790 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10651_
timestamp 0
transform 1 0 15230 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10654_
timestamp 0
transform -1 0 11730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10656_
timestamp 0
transform 1 0 12230 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__10658_
timestamp 0
transform -1 0 11890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10661_
timestamp 0
transform -1 0 13430 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10663_
timestamp 0
transform -1 0 11930 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__10666_
timestamp 0
transform -1 0 9750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10668_
timestamp 0
transform 1 0 11170 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10670_
timestamp 0
transform -1 0 10970 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__10673_
timestamp 0
transform -1 0 10790 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__10675_
timestamp 0
transform -1 0 10370 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__10678_
timestamp 0
transform 1 0 11150 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10680_
timestamp 0
transform -1 0 9690 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__10682_
timestamp 0
transform -1 0 10090 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__10685_
timestamp 0
transform 1 0 9230 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10687_
timestamp 0
transform -1 0 8730 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__10769_
timestamp 0
transform -1 0 4870 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__10772_
timestamp 0
transform 1 0 5650 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__10774_
timestamp 0
transform 1 0 5570 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__10777_
timestamp 0
transform 1 0 5450 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__10779_
timestamp 0
transform 1 0 5790 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__10781_
timestamp 0
transform -1 0 5830 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__10784_
timestamp 0
transform 1 0 5350 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__10786_
timestamp 0
transform -1 0 6770 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__10788_
timestamp 0
transform -1 0 6130 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__10791_
timestamp 0
transform 1 0 6650 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__10793_
timestamp 0
transform -1 0 5330 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__10796_
timestamp 0
transform 1 0 6170 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__10798_
timestamp 0
transform 1 0 5610 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__10800_
timestamp 0
transform 1 0 6330 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__10803_
timestamp 0
transform 1 0 5770 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__10805_
timestamp 0
transform 1 0 5770 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__10808_
timestamp 0
transform 1 0 5110 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__10810_
timestamp 0
transform 1 0 1110 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__10812_
timestamp 0
transform 1 0 1250 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__10815_
timestamp 0
transform -1 0 1430 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__10817_
timestamp 0
transform 1 0 2790 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__10819_
timestamp 0
transform 1 0 2750 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__10822_
timestamp 0
transform -1 0 1870 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__10824_
timestamp 0
transform -1 0 2810 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__10827_
timestamp 0
transform -1 0 5010 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__10829_
timestamp 0
transform -1 0 470 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__10831_
timestamp 0
transform 1 0 1510 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__10834_
timestamp 0
transform 1 0 2270 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__10836_
timestamp 0
transform 1 0 1890 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__10839_
timestamp 0
transform 1 0 3070 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__10841_
timestamp 0
transform 1 0 3030 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__10843_
timestamp 0
transform -1 0 2810 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__10846_
timestamp 0
transform 1 0 4850 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__10848_
timestamp 0
transform -1 0 3190 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__10850_
timestamp 0
transform -1 0 1350 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__10853_
timestamp 0
transform 1 0 1830 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__10855_
timestamp 0
transform 1 0 3890 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__10858_
timestamp 0
transform 1 0 3410 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__10860_
timestamp 0
transform 1 0 3590 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__10862_
timestamp 0
transform 1 0 2890 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__10865_
timestamp 0
transform 1 0 3590 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__10867_
timestamp 0
transform 1 0 750 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__10870_
timestamp 0
transform 1 0 1850 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__10872_
timestamp 0
transform -1 0 2070 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__10874_
timestamp 0
transform -1 0 2290 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__10877_
timestamp 0
transform 1 0 2210 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__10879_
timestamp 0
transform -1 0 1950 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__10881_
timestamp 0
transform -1 0 2130 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__10884_
timestamp 0
transform -1 0 2350 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__10886_
timestamp 0
transform 1 0 2450 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__10889_
timestamp 0
transform 1 0 3290 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__10891_
timestamp 0
transform -1 0 4510 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__10893_
timestamp 0
transform -1 0 4470 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__10896_
timestamp 0
transform 1 0 4530 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__10898_
timestamp 0
transform -1 0 4710 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__10900_
timestamp 0
transform -1 0 8370 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__10903_
timestamp 0
transform 1 0 5510 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__10905_
timestamp 0
transform -1 0 2490 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__10908_
timestamp 0
transform -1 0 3610 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__10910_
timestamp 0
transform 1 0 3950 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__10912_
timestamp 0
transform 1 0 4790 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__10915_
timestamp 0
transform -1 0 4130 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__10917_
timestamp 0
transform 1 0 5070 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__10920_
timestamp 0
transform 1 0 4850 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__10922_
timestamp 0
transform -1 0 5250 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__10924_
timestamp 0
transform -1 0 1050 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__10927_
timestamp 0
transform 1 0 5650 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__10929_
timestamp 0
transform 1 0 5390 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__10931_
timestamp 0
transform 1 0 3670 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__10934_
timestamp 0
transform 1 0 1630 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__10936_
timestamp 0
transform 1 0 1770 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__10939_
timestamp 0
transform -1 0 3850 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__10941_
timestamp 0
transform 1 0 1850 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__10943_
timestamp 0
transform 1 0 3670 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__10946_
timestamp 0
transform 1 0 4070 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__10948_
timestamp 0
transform -1 0 4550 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__10951_
timestamp 0
transform -1 0 5230 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__10953_
timestamp 0
transform -1 0 4790 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__10955_
timestamp 0
transform -1 0 1790 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__10958_
timestamp 0
transform 1 0 1710 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__10960_
timestamp 0
transform 1 0 3310 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__10962_
timestamp 0
transform 1 0 2770 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__10965_
timestamp 0
transform -1 0 3410 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__10967_
timestamp 0
transform 1 0 4430 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__10970_
timestamp 0
transform 1 0 3890 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__10972_
timestamp 0
transform 1 0 4910 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__10974_
timestamp 0
transform -1 0 5790 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__10977_
timestamp 0
transform 1 0 3810 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__10979_
timestamp 0
transform 1 0 1290 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__10982_
timestamp 0
transform 1 0 2470 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__10984_
timestamp 0
transform 1 0 2890 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__10986_
timestamp 0
transform 1 0 3230 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__10989_
timestamp 0
transform 1 0 4870 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__10991_
timestamp 0
transform 1 0 5150 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__10993_
timestamp 0
transform 1 0 5450 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__10996_
timestamp 0
transform 1 0 1970 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__10998_
timestamp 0
transform -1 0 1290 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__11001_
timestamp 0
transform 1 0 2510 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__11003_
timestamp 0
transform -1 0 3690 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__11005_
timestamp 0
transform 1 0 2910 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__11008_
timestamp 0
transform 1 0 3450 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__11010_
timestamp 0
transform 1 0 4270 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__11012_
timestamp 0
transform -1 0 4610 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__11015_
timestamp 0
transform 1 0 5350 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__11017_
timestamp 0
transform 1 0 5750 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__11020_
timestamp 0
transform -1 0 4950 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__11022_
timestamp 0
transform -1 0 4790 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__11024_
timestamp 0
transform -1 0 1310 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__11027_
timestamp 0
transform -1 0 2170 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__11029_
timestamp 0
transform -1 0 1450 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__11032_
timestamp 0
transform -1 0 2370 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__11034_
timestamp 0
transform 1 0 1410 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__11036_
timestamp 0
transform 1 0 2210 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__11039_
timestamp 0
transform 1 0 4270 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__11041_
timestamp 0
transform -1 0 4590 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__11043_
timestamp 0
transform 1 0 5250 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__11046_
timestamp 0
transform -1 0 5370 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__11048_
timestamp 0
transform -1 0 4170 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__11051_
timestamp 0
transform -1 0 2810 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__11053_
timestamp 0
transform -1 0 1610 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__11055_
timestamp 0
transform -1 0 1990 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__11058_
timestamp 0
transform -1 0 2650 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__11060_
timestamp 0
transform -1 0 2490 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__11063_
timestamp 0
transform 1 0 4930 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__11065_
timestamp 0
transform 1 0 5190 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__11067_
timestamp 0
transform -1 0 3350 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__11070_
timestamp 0
transform 1 0 3610 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__11072_
timestamp 0
transform -1 0 4050 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__11074_
timestamp 0
transform 1 0 3270 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__11077_
timestamp 0
transform -1 0 2330 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__11079_
timestamp 0
transform 1 0 2630 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__11082_
timestamp 0
transform 1 0 3070 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__11084_
timestamp 0
transform 1 0 3230 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__11086_
timestamp 0
transform 1 0 4470 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__11089_
timestamp 0
transform -1 0 5490 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__11091_
timestamp 0
transform 1 0 2150 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__11094_
timestamp 0
transform 1 0 2810 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__11096_
timestamp 0
transform -1 0 3550 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__11098_
timestamp 0
transform -1 0 3970 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__11101_
timestamp 0
transform -1 0 3450 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__11103_
timestamp 0
transform -1 0 4390 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__11105_
timestamp 0
transform 1 0 4110 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__11108_
timestamp 0
transform 1 0 4510 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__11110_
timestamp 0
transform 1 0 4230 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__11113_
timestamp 0
transform -1 0 5750 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__11115_
timestamp 0
transform 1 0 4670 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__11117_
timestamp 0
transform -1 0 2470 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__11120_
timestamp 0
transform -1 0 3050 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__11122_
timestamp 0
transform 1 0 3290 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__11125_
timestamp 0
transform 1 0 4570 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__11127_
timestamp 0
transform 1 0 4810 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__11129_
timestamp 0
transform -1 0 5970 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__11132_
timestamp 0
transform 1 0 3530 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__11134_
timestamp 0
transform 1 0 2350 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__11136_
timestamp 0
transform 1 0 3730 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__11139_
timestamp 0
transform 1 0 1150 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__11141_
timestamp 0
transform -1 0 4110 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__11144_
timestamp 0
transform 1 0 170 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__11146_
timestamp 0
transform -1 0 1390 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__11148_
timestamp 0
transform -1 0 1170 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__11151_
timestamp 0
transform -1 0 1670 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__11153_
timestamp 0
transform -1 0 2570 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__11155_
timestamp 0
transform 1 0 3390 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__11158_
timestamp 0
transform -1 0 3690 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__11160_
timestamp 0
transform 1 0 470 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__11163_
timestamp 0
transform -1 0 70 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__11165_
timestamp 0
transform 1 0 1690 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__11167_
timestamp 0
transform 1 0 170 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__11170_
timestamp 0
transform 1 0 570 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__11172_
timestamp 0
transform -1 0 1630 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__11175_
timestamp 0
transform -1 0 1530 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__11177_
timestamp 0
transform 1 0 1970 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__11179_
timestamp 0
transform 1 0 2110 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__11182_
timestamp 0
transform -1 0 1730 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__11184_
timestamp 0
transform 1 0 1550 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__11186_
timestamp 0
transform 1 0 610 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__11189_
timestamp 0
transform 1 0 1310 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__11191_
timestamp 0
transform 1 0 910 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__11194_
timestamp 0
transform -1 0 1330 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__11196_
timestamp 0
transform -1 0 950 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__11198_
timestamp 0
transform 1 0 1090 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__11201_
timestamp 0
transform -1 0 1310 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__11203_
timestamp 0
transform 1 0 1990 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__11206_
timestamp 0
transform 1 0 2010 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__11208_
timestamp 0
transform -1 0 630 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__11210_
timestamp 0
transform -1 0 1590 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__11213_
timestamp 0
transform -1 0 70 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__11215_
timestamp 0
transform 1 0 330 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__11217_
timestamp 0
transform 1 0 590 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__11220_
timestamp 0
transform -1 0 70 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__11222_
timestamp 0
transform -1 0 70 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__11225_
timestamp 0
transform -1 0 310 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__11227_
timestamp 0
transform -1 0 2710 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__11229_
timestamp 0
transform -1 0 330 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__11232_
timestamp 0
transform 1 0 350 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__11234_
timestamp 0
transform 1 0 170 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__11237_
timestamp 0
transform -1 0 70 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__11239_
timestamp 0
transform 1 0 330 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__11241_
timestamp 0
transform -1 0 70 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__11244_
timestamp 0
transform -1 0 230 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__11246_
timestamp 0
transform -1 0 1170 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__11248_
timestamp 0
transform -1 0 70 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__11251_
timestamp 0
transform -1 0 810 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__11253_
timestamp 0
transform -1 0 190 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__11256_
timestamp 0
transform -1 0 230 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__11258_
timestamp 0
transform -1 0 570 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__11260_
timestamp 0
transform -1 0 370 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__11263_
timestamp 0
transform -1 0 190 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__11265_
timestamp 0
transform 1 0 170 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__11267_
timestamp 0
transform -1 0 70 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__11270_
timestamp 0
transform -1 0 970 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__11272_
timestamp 0
transform 1 0 490 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__11275_
timestamp 0
transform -1 0 610 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__11277_
timestamp 0
transform -1 0 470 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__11279_
timestamp 0
transform 1 0 590 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__11282_
timestamp 0
transform -1 0 170 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__11284_
timestamp 0
transform 1 0 450 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__11287_
timestamp 0
transform 1 0 50 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__11289_
timestamp 0
transform 1 0 290 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__11291_
timestamp 0
transform 1 0 870 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__11294_
timestamp 0
transform -1 0 1370 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__11296_
timestamp 0
transform -1 0 630 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__11298_
timestamp 0
transform -1 0 1210 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__11301_
timestamp 0
transform 1 0 910 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__11303_
timestamp 0
transform 1 0 590 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__11306_
timestamp 0
transform 1 0 830 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__11308_
timestamp 0
transform -1 0 1010 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__11310_
timestamp 0
transform 1 0 170 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__11313_
timestamp 0
transform 1 0 570 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__11315_
timestamp 0
transform 1 0 710 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__11318_
timestamp 0
transform -1 0 890 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__11320_
timestamp 0
transform -1 0 70 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__11322_
timestamp 0
transform -1 0 1130 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__11325_
timestamp 0
transform -1 0 1010 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__11327_
timestamp 0
transform -1 0 1330 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__11329_
timestamp 0
transform 1 0 1150 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__11332_
timestamp 0
transform 1 0 1290 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__11334_
timestamp 0
transform -1 0 570 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__11337_
timestamp 0
transform -1 0 610 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__11339_
timestamp 0
transform 1 0 1390 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__11341_
timestamp 0
transform 1 0 1350 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__11344_
timestamp 0
transform -1 0 1010 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__11346_
timestamp 0
transform 1 0 1150 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__11349_
timestamp 0
transform -1 0 750 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__11351_
timestamp 0
transform -1 0 1110 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__11353_
timestamp 0
transform -1 0 890 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__11356_
timestamp 0
transform 1 0 830 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__11358_
timestamp 0
transform 1 0 1230 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__11360_
timestamp 0
transform -1 0 1550 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__11363_
timestamp 0
transform 1 0 1670 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__11365_
timestamp 0
transform 1 0 1770 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__11368_
timestamp 0
transform -1 0 1510 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__11370_
timestamp 0
transform -1 0 1690 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__11372_
timestamp 0
transform -1 0 1470 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__11375_
timestamp 0
transform -1 0 2390 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__11377_
timestamp 0
transform -1 0 2530 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__11379_
timestamp 0
transform -1 0 1730 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__11382_
timestamp 0
transform 1 0 4250 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__11384_
timestamp 0
transform -1 0 3990 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__11387_
timestamp 0
transform 1 0 5990 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__11389_
timestamp 0
transform -1 0 6130 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__11391_
timestamp 0
transform -1 0 3610 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__11394_
timestamp 0
transform 1 0 3810 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__11396_
timestamp 0
transform -1 0 4910 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__11399_
timestamp 0
transform 1 0 5330 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__11401_
timestamp 0
transform 1 0 4970 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__11403_
timestamp 0
transform 1 0 5950 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__11406_
timestamp 0
transform -1 0 2810 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__11408_
timestamp 0
transform 1 0 3110 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__11410_
timestamp 0
transform 1 0 4230 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__11413_
timestamp 0
transform 1 0 5230 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__11415_
timestamp 0
transform -1 0 5390 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__11418_
timestamp 0
transform 1 0 5330 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__11420_
timestamp 0
transform 1 0 5210 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__11422_
timestamp 0
transform -1 0 3750 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__11425_
timestamp 0
transform 1 0 6670 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__11427_
timestamp 0
transform 1 0 7190 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__11430_
timestamp 0
transform 1 0 6530 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__11432_
timestamp 0
transform 1 0 6130 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__11434_
timestamp 0
transform 1 0 3830 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__11437_
timestamp 0
transform 1 0 6710 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__11439_
timestamp 0
transform 1 0 6870 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__11441_
timestamp 0
transform -1 0 6150 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__11444_
timestamp 0
transform 1 0 7010 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__11446_
timestamp 0
transform -1 0 3950 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__11449_
timestamp 0
transform 1 0 4170 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__11451_
timestamp 0
transform -1 0 6270 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__11453_
timestamp 0
transform 1 0 6910 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__11456_
timestamp 0
transform -1 0 7430 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__11458_
timestamp 0
transform -1 0 6430 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__11461_
timestamp 0
transform -1 0 6770 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__11463_
timestamp 0
transform 1 0 6590 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__11465_
timestamp 0
transform -1 0 4330 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__11468_
timestamp 0
transform 1 0 4710 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__11470_
timestamp 0
transform 1 0 5330 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__11472_
timestamp 0
transform 1 0 6090 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__11475_
timestamp 0
transform 1 0 6790 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__11477_
timestamp 0
transform 1 0 5710 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__11480_
timestamp 0
transform -1 0 3430 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__11482_
timestamp 0
transform 1 0 3690 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__11484_
timestamp 0
transform 1 0 5790 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__11487_
timestamp 0
transform 1 0 6150 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__11489_
timestamp 0
transform 1 0 5830 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__11492_
timestamp 0
transform 1 0 2670 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__11494_
timestamp 0
transform -1 0 3530 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__11496_
timestamp 0
transform 1 0 3370 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__11499_
timestamp 0
transform -1 0 6090 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__11501_
timestamp 0
transform -1 0 5930 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__11503_
timestamp 0
transform -1 0 4970 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__11506_
timestamp 0
transform -1 0 4350 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__11508_
timestamp 0
transform -1 0 3850 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__11511_
timestamp 0
transform 1 0 4630 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__11513_
timestamp 0
transform 1 0 5190 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__11515_
timestamp 0
transform 1 0 4170 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__11518_
timestamp 0
transform 1 0 3310 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__11520_
timestamp 0
transform -1 0 3570 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__11522_
timestamp 0
transform -1 0 4530 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__11525_
timestamp 0
transform 1 0 5290 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__11527_
timestamp 0
transform 1 0 5130 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__11530_
timestamp 0
transform -1 0 3810 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__11532_
timestamp 0
transform 1 0 2070 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__11534_
timestamp 0
transform 1 0 2730 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__11537_
timestamp 0
transform -1 0 2510 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__11539_
timestamp 0
transform -1 0 2790 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__11542_
timestamp 0
transform -1 0 3330 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__11544_
timestamp 0
transform -1 0 2330 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__11546_
timestamp 0
transform -1 0 2470 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__11549_
timestamp 0
transform 1 0 2050 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__11551_
timestamp 0
transform 1 0 2750 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__11553_
timestamp 0
transform 1 0 3270 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__11556_
timestamp 0
transform 1 0 2650 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__11558_
timestamp 0
transform 1 0 2970 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__11561_
timestamp 0
transform 1 0 3970 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__11563_
timestamp 0
transform 1 0 3130 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__11565_
timestamp 0
transform 1 0 3730 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__11568_
timestamp 0
transform -1 0 3310 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__11570_
timestamp 0
transform 1 0 4210 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__11573_
timestamp 0
transform -1 0 3470 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__11575_
timestamp 0
transform 1 0 4870 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__11577_
timestamp 0
transform 1 0 4250 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__11580_
timestamp 0
transform 1 0 3370 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__11582_
timestamp 0
transform 1 0 5130 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__11584_
timestamp 0
transform -1 0 3670 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__11587_
timestamp 0
transform 1 0 3330 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__11589_
timestamp 0
transform -1 0 3150 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__11592_
timestamp 0
transform -1 0 3830 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__11594_
timestamp 0
transform 1 0 3870 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__11596_
timestamp 0
transform -1 0 4850 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__11599_
timestamp 0
transform 1 0 4410 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__11601_
timestamp 0
transform 1 0 6670 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__11604_
timestamp 0
transform 1 0 3970 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__11606_
timestamp 0
transform 1 0 4810 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__11608_
timestamp 0
transform -1 0 3750 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__11611_
timestamp 0
transform -1 0 4270 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__11693_
timestamp 0
transform 1 0 11350 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__11695_
timestamp 0
transform 1 0 13290 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__11698_
timestamp 0
transform -1 0 11790 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__11700_
timestamp 0
transform -1 0 11870 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__11703_
timestamp 0
transform -1 0 10950 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__11705_
timestamp 0
transform -1 0 11910 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__11707_
timestamp 0
transform 1 0 11510 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__11710_
timestamp 0
transform 1 0 9630 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__11712_
timestamp 0
transform -1 0 10950 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__11714_
timestamp 0
transform 1 0 11430 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__11717_
timestamp 0
transform -1 0 13510 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__11719_
timestamp 0
transform -1 0 13570 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__11722_
timestamp 0
transform -1 0 12950 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__11724_
timestamp 0
transform 1 0 12870 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__11726_
timestamp 0
transform 1 0 13190 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__11729_
timestamp 0
transform 1 0 12850 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__11731_
timestamp 0
transform -1 0 12790 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__11734_
timestamp 0
transform -1 0 13230 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__11736_
timestamp 0
transform -1 0 13070 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__11738_
timestamp 0
transform -1 0 12370 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__11741_
timestamp 0
transform 1 0 12990 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__11743_
timestamp 0
transform -1 0 14590 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__11745_
timestamp 0
transform -1 0 12990 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__11748_
timestamp 0
transform -1 0 12610 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__11750_
timestamp 0
transform 1 0 12490 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__11753_
timestamp 0
transform -1 0 16170 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__11755_
timestamp 0
transform 1 0 15010 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__11757_
timestamp 0
transform -1 0 16330 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__11760_
timestamp 0
transform 1 0 14850 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__11762_
timestamp 0
transform 1 0 13330 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__11765_
timestamp 0
transform 1 0 13390 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__11767_
timestamp 0
transform -1 0 12930 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__11769_
timestamp 0
transform 1 0 13150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__11772_
timestamp 0
transform 1 0 14890 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__11774_
timestamp 0
transform -1 0 13310 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__11776_
timestamp 0
transform 1 0 12610 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__11779_
timestamp 0
transform -1 0 13970 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__11781_
timestamp 0
transform 1 0 15310 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__11784_
timestamp 0
transform -1 0 13190 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__11786_
timestamp 0
transform -1 0 12890 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__11788_
timestamp 0
transform 1 0 12850 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__11791_
timestamp 0
transform -1 0 12030 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__11793_
timestamp 0
transform -1 0 15450 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__11796_
timestamp 0
transform -1 0 15170 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__11798_
timestamp 0
transform 1 0 15650 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__11800_
timestamp 0
transform 1 0 15370 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__11803_
timestamp 0
transform -1 0 14930 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__11805_
timestamp 0
transform -1 0 15210 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__11807_
timestamp 0
transform -1 0 13430 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__11810_
timestamp 0
transform -1 0 15570 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__11812_
timestamp 0
transform 1 0 13450 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__11815_
timestamp 0
transform 1 0 13290 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__11817_
timestamp 0
transform -1 0 12390 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__11819_
timestamp 0
transform 1 0 12490 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__11822_
timestamp 0
transform -1 0 12710 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__11824_
timestamp 0
transform 1 0 9370 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__11826_
timestamp 0
transform -1 0 8870 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__11829_
timestamp 0
transform 1 0 15330 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__11831_
timestamp 0
transform 1 0 14710 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__11834_
timestamp 0
transform -1 0 14830 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__11836_
timestamp 0
transform 1 0 13630 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__11838_
timestamp 0
transform 1 0 13570 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__11841_
timestamp 0
transform 1 0 13170 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__11843_
timestamp 0
transform 1 0 13250 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__11846_
timestamp 0
transform -1 0 13010 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__11848_
timestamp 0
transform 1 0 15370 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__11850_
timestamp 0
transform -1 0 12650 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__11853_
timestamp 0
transform 1 0 13410 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__11855_
timestamp 0
transform 1 0 16170 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__11857_
timestamp 0
transform -1 0 14750 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__11860_
timestamp 0
transform -1 0 15650 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__11862_
timestamp 0
transform 1 0 17030 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__11865_
timestamp 0
transform 1 0 15930 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__11867_
timestamp 0
transform 1 0 17090 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__11869_
timestamp 0
transform 1 0 16790 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__11872_
timestamp 0
transform -1 0 14930 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__11874_
timestamp 0
transform -1 0 13670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__11877_
timestamp 0
transform 1 0 15170 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__11879_
timestamp 0
transform 1 0 14430 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__11881_
timestamp 0
transform 1 0 14470 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__11884_
timestamp 0
transform -1 0 15810 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__11886_
timestamp 0
transform -1 0 16830 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__11888_
timestamp 0
transform 1 0 16970 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__11891_
timestamp 0
transform 1 0 16810 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__11893_
timestamp 0
transform -1 0 17030 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__11896_
timestamp 0
transform -1 0 15490 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__11898_
timestamp 0
transform 1 0 14010 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__11900_
timestamp 0
transform -1 0 16950 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__11903_
timestamp 0
transform 1 0 14970 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__11905_
timestamp 0
transform 1 0 15510 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__11908_
timestamp 0
transform -1 0 16570 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__11910_
timestamp 0
transform -1 0 16370 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__11912_
timestamp 0
transform 1 0 16490 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__11915_
timestamp 0
transform -1 0 15190 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__11917_
timestamp 0
transform -1 0 14730 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__11919_
timestamp 0
transform 1 0 14430 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__11922_
timestamp 0
transform -1 0 15230 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__11924_
timestamp 0
transform 1 0 15290 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__11927_
timestamp 0
transform 1 0 16450 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__11929_
timestamp 0
transform -1 0 16210 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__11931_
timestamp 0
transform 1 0 16310 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__11934_
timestamp 0
transform -1 0 16670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__11936_
timestamp 0
transform 1 0 16910 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__11938_
timestamp 0
transform -1 0 15790 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__11941_
timestamp 0
transform 1 0 12870 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__11943_
timestamp 0
transform 1 0 17010 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__11946_
timestamp 0
transform 1 0 16450 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__11948_
timestamp 0
transform -1 0 16310 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__11950_
timestamp 0
transform 1 0 14570 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__11953_
timestamp 0
transform 1 0 15890 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__11955_
timestamp 0
transform 1 0 16590 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__11958_
timestamp 0
transform 1 0 15890 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__11960_
timestamp 0
transform -1 0 16470 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__11962_
timestamp 0
transform 1 0 15850 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__11965_
timestamp 0
transform 1 0 15930 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__11967_
timestamp 0
transform -1 0 13270 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__11969_
timestamp 0
transform -1 0 14370 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__11972_
timestamp 0
transform 1 0 16130 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__11974_
timestamp 0
transform 1 0 16290 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__11977_
timestamp 0
transform -1 0 15750 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__11979_
timestamp 0
transform 1 0 16010 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__11981_
timestamp 0
transform -1 0 15650 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__11984_
timestamp 0
transform -1 0 15870 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__11986_
timestamp 0
transform 1 0 15270 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__11989_
timestamp 0
transform 1 0 14970 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__11991_
timestamp 0
transform -1 0 15770 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__11993_
timestamp 0
transform -1 0 15910 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__11996_
timestamp 0
transform -1 0 15170 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__11998_
timestamp 0
transform 1 0 14690 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__12000_
timestamp 0
transform -1 0 15330 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__12003_
timestamp 0
transform -1 0 15150 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__12005_
timestamp 0
transform 1 0 14810 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__12008_
timestamp 0
transform 1 0 14710 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__12010_
timestamp 0
transform -1 0 14830 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__12012_
timestamp 0
transform -1 0 14530 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__12015_
timestamp 0
transform 1 0 15130 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__12017_
timestamp 0
transform -1 0 14890 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__12020_
timestamp 0
transform 1 0 14530 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__12022_
timestamp 0
transform 1 0 14310 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__12024_
timestamp 0
transform -1 0 14550 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__12027_
timestamp 0
transform -1 0 14370 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__12029_
timestamp 0
transform -1 0 15010 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__12031_
timestamp 0
transform -1 0 14510 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__12034_
timestamp 0
transform -1 0 14570 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__12036_
timestamp 0
transform -1 0 14090 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__12039_
timestamp 0
transform -1 0 14250 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__12041_
timestamp 0
transform 1 0 14810 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__12043_
timestamp 0
transform -1 0 14570 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__12046_
timestamp 0
transform -1 0 14070 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__12048_
timestamp 0
transform 1 0 13830 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__12051_
timestamp 0
transform -1 0 13690 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__12053_
timestamp 0
transform 1 0 13390 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__12055_
timestamp 0
transform -1 0 15850 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__12058_
timestamp 0
transform -1 0 16050 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__12060_
timestamp 0
transform 1 0 12870 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__12062_
timestamp 0
transform 1 0 16170 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__12065_
timestamp 0
transform -1 0 17070 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__12067_
timestamp 0
transform 1 0 16730 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__12070_
timestamp 0
transform 1 0 12870 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__12072_
timestamp 0
transform -1 0 16930 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__12074_
timestamp 0
transform -1 0 16950 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__12077_
timestamp 0
transform -1 0 12590 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__12079_
timestamp 0
transform 1 0 15590 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__12081_
timestamp 0
transform 1 0 13810 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__12084_
timestamp 0
transform 1 0 16590 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__12086_
timestamp 0
transform -1 0 16230 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__12089_
timestamp 0
transform 1 0 16770 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__12091_
timestamp 0
transform 1 0 16810 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__12093_
timestamp 0
transform -1 0 15450 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__12096_
timestamp 0
transform 1 0 16390 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__12098_
timestamp 0
transform -1 0 15190 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__12101_
timestamp 0
transform 1 0 13810 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__12103_
timestamp 0
transform -1 0 13530 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__12105_
timestamp 0
transform -1 0 13190 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12108_
timestamp 0
transform -1 0 15570 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__12110_
timestamp 0
transform 1 0 16590 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__12112_
timestamp 0
transform -1 0 16350 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__12115_
timestamp 0
transform 1 0 16390 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__12117_
timestamp 0
transform -1 0 16810 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12120_
timestamp 0
transform 1 0 16490 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12122_
timestamp 0
transform 1 0 16330 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12124_
timestamp 0
transform -1 0 15710 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12127_
timestamp 0
transform -1 0 13330 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12129_
timestamp 0
transform 1 0 17050 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__12132_
timestamp 0
transform -1 0 16270 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__12134_
timestamp 0
transform 1 0 16890 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__12136_
timestamp 0
transform 1 0 16890 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__12139_
timestamp 0
transform 1 0 17070 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__12141_
timestamp 0
transform -1 0 16570 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__12143_
timestamp 0
transform 1 0 16710 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__12146_
timestamp 0
transform 1 0 16770 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__12148_
timestamp 0
transform 1 0 14390 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__12151_
timestamp 0
transform 1 0 15050 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__12153_
timestamp 0
transform -1 0 15890 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__12155_
timestamp 0
transform 1 0 16670 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__12158_
timestamp 0
transform 1 0 17010 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__12160_
timestamp 0
transform 1 0 16870 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__12163_
timestamp 0
transform 1 0 17010 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__12165_
timestamp 0
transform -1 0 16590 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__12167_
timestamp 0
transform -1 0 15370 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__12170_
timestamp 0
transform 1 0 13810 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__12172_
timestamp 0
transform 1 0 15870 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__12174_
timestamp 0
transform -1 0 15990 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__12177_
timestamp 0
transform 1 0 16310 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__12179_
timestamp 0
transform 1 0 16250 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__12182_
timestamp 0
transform -1 0 16410 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__12184_
timestamp 0
transform -1 0 16290 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__12186_
timestamp 0
transform -1 0 16450 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__12189_
timestamp 0
transform -1 0 14970 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__12191_
timestamp 0
transform 1 0 14090 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__12193_
timestamp 0
transform -1 0 15990 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__12196_
timestamp 0
transform -1 0 16250 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__12198_
timestamp 0
transform -1 0 16310 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__12201_
timestamp 0
transform 1 0 15410 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__12203_
timestamp 0
transform 1 0 15130 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__12205_
timestamp 0
transform -1 0 16430 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__12208_
timestamp 0
transform 1 0 15590 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__12210_
timestamp 0
transform -1 0 15210 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__12213_
timestamp 0
transform -1 0 16130 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__12215_
timestamp 0
transform -1 0 15070 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__12217_
timestamp 0
transform 1 0 13150 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__12220_
timestamp 0
transform -1 0 14810 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__12222_
timestamp 0
transform 1 0 15830 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__12224_
timestamp 0
transform -1 0 15990 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__12227_
timestamp 0
transform -1 0 15830 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__12229_
timestamp 0
transform -1 0 15450 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__12232_
timestamp 0
transform -1 0 15750 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__12234_
timestamp 0
transform -1 0 14530 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__12236_
timestamp 0
transform -1 0 14410 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__12239_
timestamp 0
transform 1 0 14850 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__12241_
timestamp 0
transform -1 0 14590 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__12244_
timestamp 0
transform -1 0 16130 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__12246_
timestamp 0
transform -1 0 15230 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__12248_
timestamp 0
transform -1 0 15350 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__12251_
timestamp 0
transform -1 0 15250 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12253_
timestamp 0
transform -1 0 14690 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__12255_
timestamp 0
transform -1 0 13770 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__12258_
timestamp 0
transform 1 0 13570 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__12260_
timestamp 0
transform -1 0 14030 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__12263_
timestamp 0
transform 1 0 14910 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__12265_
timestamp 0
transform 1 0 14950 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12267_
timestamp 0
transform -1 0 14550 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12270_
timestamp 0
transform 1 0 14290 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__12272_
timestamp 0
transform 1 0 14130 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__12275_
timestamp 0
transform -1 0 14230 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__12277_
timestamp 0
transform -1 0 14450 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__12279_
timestamp 0
transform -1 0 14490 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__12282_
timestamp 0
transform 1 0 15390 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12284_
timestamp 0
transform 1 0 14510 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__12286_
timestamp 0
transform 1 0 14430 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__12289_
timestamp 0
transform -1 0 14110 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__12291_
timestamp 0
transform -1 0 13830 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__12294_
timestamp 0
transform 1 0 13510 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__12296_
timestamp 0
transform -1 0 14430 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12298_
timestamp 0
transform 1 0 14290 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__12301_
timestamp 0
transform -1 0 14170 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__12303_
timestamp 0
transform -1 0 13870 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12305_
timestamp 0
transform -1 0 11910 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__12308_
timestamp 0
transform -1 0 10970 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__12310_
timestamp 0
transform 1 0 11210 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__12313_
timestamp 0
transform -1 0 11290 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__12315_
timestamp 0
transform 1 0 10750 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__12317_
timestamp 0
transform -1 0 10070 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__12320_
timestamp 0
transform 1 0 10270 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__12322_
timestamp 0
transform -1 0 10130 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__12325_
timestamp 0
transform -1 0 10750 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__12327_
timestamp 0
transform 1 0 11110 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__12329_
timestamp 0
transform 1 0 10570 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__12332_
timestamp 0
transform -1 0 11690 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__12334_
timestamp 0
transform -1 0 11110 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__12336_
timestamp 0
transform -1 0 10870 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__12339_
timestamp 0
transform 1 0 10270 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__12341_
timestamp 0
transform 1 0 11170 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__12344_
timestamp 0
transform 1 0 11670 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__12346_
timestamp 0
transform -1 0 12350 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__12348_
timestamp 0
transform -1 0 12050 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__12351_
timestamp 0
transform -1 0 10650 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__12353_
timestamp 0
transform 1 0 11130 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__12356_
timestamp 0
transform 1 0 10670 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__12358_
timestamp 0
transform -1 0 10490 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__12360_
timestamp 0
transform -1 0 10050 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__12363_
timestamp 0
transform -1 0 9790 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12365_
timestamp 0
transform 1 0 9970 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__12367_
timestamp 0
transform 1 0 10270 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__12370_
timestamp 0
transform 1 0 12690 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__12372_
timestamp 0
transform 1 0 12190 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__12375_
timestamp 0
transform -1 0 10250 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__12377_
timestamp 0
transform 1 0 9910 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12379_
timestamp 0
transform -1 0 9430 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__12382_
timestamp 0
transform 1 0 10670 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__12384_
timestamp 0
transform 1 0 9790 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__12387_
timestamp 0
transform -1 0 9770 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__12389_
timestamp 0
transform 1 0 12490 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__12391_
timestamp 0
transform -1 0 12350 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__12394_
timestamp 0
transform -1 0 10890 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__12396_
timestamp 0
transform -1 0 10050 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__12398_
timestamp 0
transform -1 0 9930 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__12401_
timestamp 0
transform 1 0 10390 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__12403_
timestamp 0
transform 1 0 11330 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__12406_
timestamp 0
transform 1 0 10670 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__12408_
timestamp 0
transform -1 0 10630 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__12410_
timestamp 0
transform -1 0 10490 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__12413_
timestamp 0
transform 1 0 10510 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__12415_
timestamp 0
transform 1 0 11890 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__12417_
timestamp 0
transform -1 0 11670 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__12420_
timestamp 0
transform -1 0 11770 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__12422_
timestamp 0
transform -1 0 10350 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12425_
timestamp 0
transform 1 0 10170 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12427_
timestamp 0
transform -1 0 11110 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__12429_
timestamp 0
transform 1 0 10990 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12432_
timestamp 0
transform -1 0 11630 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__12434_
timestamp 0
transform -1 0 11250 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__12437_
timestamp 0
transform -1 0 11810 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12439_
timestamp 0
transform -1 0 11370 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__12441_
timestamp 0
transform 1 0 11490 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12444_
timestamp 0
transform -1 0 12030 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__12446_
timestamp 0
transform -1 0 12110 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12448_
timestamp 0
transform -1 0 11950 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__12451_
timestamp 0
transform 1 0 12050 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__12453_
timestamp 0
transform -1 0 11710 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__12456_
timestamp 0
transform -1 0 14010 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__12458_
timestamp 0
transform -1 0 14090 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__12460_
timestamp 0
transform -1 0 11730 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__12463_
timestamp 0
transform 1 0 14150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__12465_
timestamp 0
transform -1 0 13570 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__12468_
timestamp 0
transform 1 0 14270 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__12470_
timestamp 0
transform 1 0 13950 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__12472_
timestamp 0
transform 1 0 16430 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__12475_
timestamp 0
transform -1 0 15570 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__12477_
timestamp 0
transform -1 0 13730 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__12479_
timestamp 0
transform -1 0 13790 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__12482_
timestamp 0
transform 1 0 13670 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__12484_
timestamp 0
transform -1 0 14030 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__12487_
timestamp 0
transform -1 0 14310 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__12489_
timestamp 0
transform -1 0 13770 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__12491_
timestamp 0
transform -1 0 14070 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__12494_
timestamp 0
transform -1 0 14490 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__12496_
timestamp 0
transform -1 0 14770 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__12499_
timestamp 0
transform -1 0 16630 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__12501_
timestamp 0
transform -1 0 16670 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__12503_
timestamp 0
transform -1 0 13490 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__12506_
timestamp 0
transform -1 0 12110 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__12508_
timestamp 0
transform -1 0 11810 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__12510_
timestamp 0
transform 1 0 12470 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__12513_
timestamp 0
transform -1 0 11970 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__12515_
timestamp 0
transform -1 0 12330 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__12518_
timestamp 0
transform -1 0 12170 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__12520_
timestamp 0
transform 1 0 11010 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__12522_
timestamp 0
transform 1 0 11410 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__12525_
timestamp 0
transform -1 0 9550 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__12527_
timestamp 0
transform -1 0 9790 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__12530_
timestamp 0
transform -1 0 11610 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__12532_
timestamp 0
transform 1 0 11190 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__12534_
timestamp 0
transform 1 0 10810 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__12617_
timestamp 0
transform -1 0 11410 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__12619_
timestamp 0
transform 1 0 11510 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__12621_
timestamp 0
transform -1 0 10850 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__12624_
timestamp 0
transform -1 0 11550 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__12626_
timestamp 0
transform -1 0 11570 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__12629_
timestamp 0
transform 1 0 11350 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__12631_
timestamp 0
transform 1 0 11210 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__12633_
timestamp 0
transform 1 0 11650 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__12636_
timestamp 0
transform -1 0 11650 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__12638_
timestamp 0
transform 1 0 11650 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__12640_
timestamp 0
transform -1 0 11670 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__12643_
timestamp 0
transform -1 0 11330 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__12645_
timestamp 0
transform -1 0 11170 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__12648_
timestamp 0
transform 1 0 11090 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__12650_
timestamp 0
transform -1 0 10950 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__12652_
timestamp 0
transform 1 0 11150 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__12655_
timestamp 0
transform 1 0 11210 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__12657_
timestamp 0
transform 1 0 11350 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__12660_
timestamp 0
transform -1 0 12530 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__12662_
timestamp 0
transform -1 0 12390 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__12664_
timestamp 0
transform -1 0 12110 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__12667_
timestamp 0
transform -1 0 12030 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__12669_
timestamp 0
transform -1 0 17030 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__12671_
timestamp 0
transform 1 0 16710 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__12674_
timestamp 0
transform 1 0 16890 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__12676_
timestamp 0
transform 1 0 16930 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__12679_
timestamp 0
transform -1 0 16190 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__12681_
timestamp 0
transform 1 0 15950 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__12683_
timestamp 0
transform 1 0 16550 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__12686_
timestamp 0
transform -1 0 13130 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__12688_
timestamp 0
transform -1 0 12670 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__12691_
timestamp 0
transform 1 0 12910 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__12693_
timestamp 0
transform 1 0 12070 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__12695_
timestamp 0
transform 1 0 11370 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__12698_
timestamp 0
transform -1 0 16430 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__12700_
timestamp 0
transform 1 0 16190 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__12702_
timestamp 0
transform -1 0 15910 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__12705_
timestamp 0
transform -1 0 16230 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__12707_
timestamp 0
transform 1 0 14490 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__12710_
timestamp 0
transform 1 0 15770 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__12712_
timestamp 0
transform -1 0 16690 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__12714_
timestamp 0
transform 1 0 16670 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__12717_
timestamp 0
transform 1 0 17090 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__12719_
timestamp 0
transform 1 0 16710 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__12722_
timestamp 0
transform 1 0 16950 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__12724_
timestamp 0
transform -1 0 14450 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__12726_
timestamp 0
transform -1 0 16990 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__12729_
timestamp 0
transform 1 0 16750 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__12731_
timestamp 0
transform -1 0 16230 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__12733_
timestamp 0
transform -1 0 13930 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__12736_
timestamp 0
transform -1 0 13670 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__12738_
timestamp 0
transform -1 0 13050 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__12741_
timestamp 0
transform -1 0 9030 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__12743_
timestamp 0
transform 1 0 9130 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__12745_
timestamp 0
transform -1 0 13390 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__12748_
timestamp 0
transform -1 0 15710 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__12750_
timestamp 0
transform 1 0 15510 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__12752_
timestamp 0
transform -1 0 13850 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__12755_
timestamp 0
transform -1 0 14610 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__12757_
timestamp 0
transform -1 0 13470 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__12760_
timestamp 0
transform -1 0 12930 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__12762_
timestamp 0
transform -1 0 12410 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__12764_
timestamp 0
transform -1 0 12250 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__12767_
timestamp 0
transform -1 0 12110 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__12769_
timestamp 0
transform 1 0 12390 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__12772_
timestamp 0
transform 1 0 14990 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__12774_
timestamp 0
transform 1 0 15170 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__12776_
timestamp 0
transform 1 0 15470 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__12779_
timestamp 0
transform 1 0 17030 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__12781_
timestamp 0
transform 1 0 16490 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__12783_
timestamp 0
transform -1 0 13210 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__12786_
timestamp 0
transform 1 0 13090 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__12788_
timestamp 0
transform 1 0 13370 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__12791_
timestamp 0
transform -1 0 12630 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__12793_
timestamp 0
transform 1 0 11930 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__12795_
timestamp 0
transform -1 0 14090 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__12798_
timestamp 0
transform 1 0 15250 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__12800_
timestamp 0
transform -1 0 15410 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__12803_
timestamp 0
transform -1 0 13510 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__12805_
timestamp 0
transform -1 0 13510 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__12807_
timestamp 0
transform 1 0 12810 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__12810_
timestamp 0
transform 1 0 13650 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__12812_
timestamp 0
transform 1 0 12750 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__12814_
timestamp 0
transform 1 0 12710 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__12817_
timestamp 0
transform -1 0 14570 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__12819_
timestamp 0
transform 1 0 15670 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__12822_
timestamp 0
transform 1 0 16410 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__12824_
timestamp 0
transform -1 0 13810 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__12826_
timestamp 0
transform -1 0 14110 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__12829_
timestamp 0
transform -1 0 13130 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__12831_
timestamp 0
transform 1 0 13130 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__12834_
timestamp 0
transform -1 0 12290 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__12836_
timestamp 0
transform 1 0 12170 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__12838_
timestamp 0
transform 1 0 13410 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__12841_
timestamp 0
transform -1 0 15350 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__12843_
timestamp 0
transform -1 0 14130 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__12845_
timestamp 0
transform 1 0 13830 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__12848_
timestamp 0
transform 1 0 13970 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__12850_
timestamp 0
transform -1 0 12770 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__12853_
timestamp 0
transform 1 0 12890 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__12855_
timestamp 0
transform -1 0 12450 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__12857_
timestamp 0
transform 1 0 12290 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__12860_
timestamp 0
transform -1 0 13350 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__12862_
timestamp 0
transform 1 0 13150 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__12864_
timestamp 0
transform -1 0 13150 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__12867_
timestamp 0
transform 1 0 15230 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__12869_
timestamp 0
transform -1 0 15270 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__12872_
timestamp 0
transform -1 0 14350 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__12874_
timestamp 0
transform 1 0 13770 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__12876_
timestamp 0
transform 1 0 14050 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__12879_
timestamp 0
transform -1 0 13030 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__12881_
timestamp 0
transform 1 0 12990 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__12884_
timestamp 0
transform -1 0 12090 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__12886_
timestamp 0
transform -1 0 12150 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__12888_
timestamp 0
transform -1 0 11450 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__12891_
timestamp 0
transform -1 0 12730 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__12893_
timestamp 0
transform -1 0 13870 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__12895_
timestamp 0
transform -1 0 13710 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__12898_
timestamp 0
transform 1 0 14010 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__12900_
timestamp 0
transform -1 0 13870 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__12903_
timestamp 0
transform -1 0 13390 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__12905_
timestamp 0
transform -1 0 12390 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__12907_
timestamp 0
transform 1 0 11790 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__12910_
timestamp 0
transform 1 0 13290 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__12912_
timestamp 0
transform 1 0 13150 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__12915_
timestamp 0
transform 1 0 14270 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__12917_
timestamp 0
transform 1 0 14690 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__12919_
timestamp 0
transform -1 0 14550 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__12922_
timestamp 0
transform 1 0 14410 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__12924_
timestamp 0
transform 1 0 14530 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__12926_
timestamp 0
transform -1 0 13550 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__12929_
timestamp 0
transform -1 0 11950 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__12931_
timestamp 0
transform 1 0 15090 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__12934_
timestamp 0
transform 1 0 14950 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__12936_
timestamp 0
transform -1 0 14010 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__12938_
timestamp 0
transform -1 0 14550 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__12941_
timestamp 0
transform -1 0 13850 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__12943_
timestamp 0
transform -1 0 14270 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__12946_
timestamp 0
transform -1 0 13210 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__12948_
timestamp 0
transform -1 0 12950 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__12950_
timestamp 0
transform -1 0 13050 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__12953_
timestamp 0
transform -1 0 12390 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__12955_
timestamp 0
transform 1 0 11950 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__12957_
timestamp 0
transform 1 0 15110 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__12960_
timestamp 0
transform -1 0 14850 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__12962_
timestamp 0
transform 1 0 13910 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__12965_
timestamp 0
transform 1 0 13190 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__12967_
timestamp 0
transform 1 0 12670 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__12969_
timestamp 0
transform -1 0 12690 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__12972_
timestamp 0
transform 1 0 15730 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__12974_
timestamp 0
transform -1 0 15990 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__12977_
timestamp 0
transform -1 0 14090 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__12979_
timestamp 0
transform -1 0 16150 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__12981_
timestamp 0
transform 1 0 14570 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__12984_
timestamp 0
transform 1 0 16230 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__12986_
timestamp 0
transform 1 0 16650 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__12988_
timestamp 0
transform -1 0 15870 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__12991_
timestamp 0
transform 1 0 16050 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__12993_
timestamp 0
transform -1 0 15650 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__12996_
timestamp 0
transform -1 0 15130 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__12998_
timestamp 0
transform -1 0 15490 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__13000_
timestamp 0
transform -1 0 16490 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__13003_
timestamp 0
transform 1 0 14250 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13005_
timestamp 0
transform -1 0 14230 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__13007_
timestamp 0
transform 1 0 16450 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__13010_
timestamp 0
transform -1 0 17010 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13012_
timestamp 0
transform -1 0 16730 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__13015_
timestamp 0
transform 1 0 15930 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13017_
timestamp 0
transform -1 0 15790 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13019_
timestamp 0
transform -1 0 15510 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13022_
timestamp 0
transform -1 0 12290 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__13024_
timestamp 0
transform 1 0 16650 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13027_
timestamp 0
transform 1 0 16130 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__13029_
timestamp 0
transform -1 0 16210 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13031_
timestamp 0
transform -1 0 16230 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__13034_
timestamp 0
transform -1 0 16810 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13036_
timestamp 0
transform 1 0 16950 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__13038_
timestamp 0
transform 1 0 16850 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13041_
timestamp 0
transform -1 0 16390 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__13043_
timestamp 0
transform -1 0 16230 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__13046_
timestamp 0
transform -1 0 16710 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__13048_
timestamp 0
transform -1 0 15470 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__13050_
timestamp 0
transform 1 0 16050 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13053_
timestamp 0
transform -1 0 16910 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__13055_
timestamp 0
transform 1 0 16950 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13058_
timestamp 0
transform 1 0 17030 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13060_
timestamp 0
transform -1 0 16890 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13062_
timestamp 0
transform -1 0 16610 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13065_
timestamp 0
transform 1 0 12630 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13067_
timestamp 0
transform -1 0 15390 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13069_
timestamp 0
transform -1 0 15730 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__13072_
timestamp 0
transform 1 0 16530 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__13074_
timestamp 0
transform 1 0 16530 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__13077_
timestamp 0
transform -1 0 17070 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__13079_
timestamp 0
transform -1 0 16650 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__13081_
timestamp 0
transform -1 0 16770 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13084_
timestamp 0
transform 1 0 14470 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13086_
timestamp 0
transform -1 0 16190 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13089_
timestamp 0
transform 1 0 16430 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13091_
timestamp 0
transform -1 0 15590 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__13093_
timestamp 0
transform 1 0 16330 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13096_
timestamp 0
transform 1 0 17010 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13098_
timestamp 0
transform 1 0 16690 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__13100_
timestamp 0
transform 1 0 16630 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__13103_
timestamp 0
transform 1 0 16730 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13105_
timestamp 0
transform 1 0 15810 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13108_
timestamp 0
transform 1 0 12610 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13110_
timestamp 0
transform 1 0 16590 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13112_
timestamp 0
transform -1 0 16130 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__13115_
timestamp 0
transform -1 0 16410 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__13117_
timestamp 0
transform 1 0 16230 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13119_
timestamp 0
transform 1 0 15970 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__13122_
timestamp 0
transform 1 0 16850 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13124_
timestamp 0
transform -1 0 14330 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13127_
timestamp 0
transform -1 0 13090 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13129_
timestamp 0
transform -1 0 14650 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13131_
timestamp 0
transform -1 0 14170 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13134_
timestamp 0
transform 1 0 9790 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13136_
timestamp 0
transform 1 0 11310 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13139_
timestamp 0
transform -1 0 15730 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__13141_
timestamp 0
transform 1 0 15550 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__13143_
timestamp 0
transform 1 0 16110 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13146_
timestamp 0
transform -1 0 15390 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13148_
timestamp 0
transform -1 0 16070 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13150_
timestamp 0
transform 1 0 13890 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13153_
timestamp 0
transform -1 0 11770 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13155_
timestamp 0
transform 1 0 11430 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13158_
timestamp 0
transform -1 0 13250 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13160_
timestamp 0
transform -1 0 15850 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13162_
timestamp 0
transform -1 0 15730 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__13165_
timestamp 0
transform -1 0 15490 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13167_
timestamp 0
transform -1 0 15230 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13170_
timestamp 0
transform -1 0 14850 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13172_
timestamp 0
transform -1 0 10970 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13174_
timestamp 0
transform -1 0 12290 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13177_
timestamp 0
transform 1 0 12810 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13179_
timestamp 0
transform -1 0 15270 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__13181_
timestamp 0
transform 1 0 15670 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13184_
timestamp 0
transform -1 0 15050 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13186_
timestamp 0
transform 1 0 14830 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13189_
timestamp 0
transform 1 0 13950 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13191_
timestamp 0
transform -1 0 10190 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13193_
timestamp 0
transform -1 0 14570 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13196_
timestamp 0
transform 1 0 14390 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13198_
timestamp 0
transform -1 0 15630 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__13201_
timestamp 0
transform 1 0 14890 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13203_
timestamp 0
transform -1 0 14610 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13205_
timestamp 0
transform 1 0 14970 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__13208_
timestamp 0
transform -1 0 14130 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13210_
timestamp 0
transform -1 0 13990 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13212_
timestamp 0
transform -1 0 13050 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13215_
timestamp 0
transform -1 0 14470 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13217_
timestamp 0
transform -1 0 14190 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13220_
timestamp 0
transform -1 0 13570 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13222_
timestamp 0
transform -1 0 13370 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13224_
timestamp 0
transform -1 0 12770 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13227_
timestamp 0
transform -1 0 13090 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13229_
timestamp 0
transform -1 0 13670 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__13231_
timestamp 0
transform -1 0 12930 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13234_
timestamp 0
transform -1 0 11490 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__13236_
timestamp 0
transform -1 0 11430 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__13239_
timestamp 0
transform 1 0 11550 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__13241_
timestamp 0
transform 1 0 10970 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13243_
timestamp 0
transform 1 0 11770 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__13246_
timestamp 0
transform -1 0 11150 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13248_
timestamp 0
transform -1 0 10450 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13251_
timestamp 0
transform -1 0 10190 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13253_
timestamp 0
transform -1 0 12110 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__13255_
timestamp 0
transform -1 0 14370 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13258_
timestamp 0
transform -1 0 11190 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13260_
timestamp 0
transform -1 0 10910 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13262_
timestamp 0
transform -1 0 10610 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__13265_
timestamp 0
transform -1 0 12050 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__13267_
timestamp 0
transform -1 0 14030 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__13270_
timestamp 0
transform 1 0 12050 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__13272_
timestamp 0
transform 1 0 11010 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13274_
timestamp 0
transform 1 0 13450 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__13277_
timestamp 0
transform -1 0 13790 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13279_
timestamp 0
transform -1 0 12410 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__13282_
timestamp 0
transform -1 0 11510 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__13284_
timestamp 0
transform -1 0 10750 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__13286_
timestamp 0
transform 1 0 10950 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__13289_
timestamp 0
transform 1 0 11610 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__13291_
timestamp 0
transform 1 0 10990 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__13293_
timestamp 0
transform 1 0 14430 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__13296_
timestamp 0
transform -1 0 14190 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__13298_
timestamp 0
transform -1 0 12310 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__13301_
timestamp 0
transform -1 0 11270 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__13303_
timestamp 0
transform -1 0 12170 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__13305_
timestamp 0
transform -1 0 13230 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__13308_
timestamp 0
transform 1 0 12810 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__13310_
timestamp 0
transform 1 0 12670 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__13313_
timestamp 0
transform -1 0 11870 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__13315_
timestamp 0
transform 1 0 13090 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__13317_
timestamp 0
transform -1 0 12630 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__13320_
timestamp 0
transform -1 0 12350 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__13322_
timestamp 0
transform 1 0 11910 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__13324_
timestamp 0
transform 1 0 11490 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__13327_
timestamp 0
transform -1 0 12110 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__13329_
timestamp 0
transform 1 0 11950 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__13332_
timestamp 0
transform 1 0 11630 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__13334_
timestamp 0
transform 1 0 12010 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__13336_
timestamp 0
transform 1 0 11850 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__13339_
timestamp 0
transform 1 0 12970 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__13341_
timestamp 0
transform -1 0 11650 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__13343_
timestamp 0
transform -1 0 11810 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13346_
timestamp 0
transform 1 0 12090 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__13348_
timestamp 0
transform 1 0 14950 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__13351_
timestamp 0
transform 1 0 15030 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13353_
timestamp 0
transform 1 0 14890 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__13355_
timestamp 0
transform -1 0 15150 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__13358_
timestamp 0
transform -1 0 11670 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13360_
timestamp 0
transform 1 0 15150 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13363_
timestamp 0
transform 1 0 12350 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__13365_
timestamp 0
transform -1 0 16850 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13367_
timestamp 0
transform 1 0 16790 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13370_
timestamp 0
transform 1 0 14830 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13372_
timestamp 0
transform -1 0 15690 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13374_
timestamp 0
transform -1 0 16090 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13377_
timestamp 0
transform -1 0 14270 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13379_
timestamp 0
transform -1 0 14810 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13382_
timestamp 0
transform 1 0 14790 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__13384_
timestamp 0
transform 1 0 14330 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13386_
timestamp 0
transform -1 0 13850 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13389_
timestamp 0
transform -1 0 14270 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__13391_
timestamp 0
transform 1 0 14310 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__13394_
timestamp 0
transform -1 0 13550 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13396_
timestamp 0
transform 1 0 14550 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13398_
timestamp 0
transform 1 0 13010 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13401_
timestamp 0
transform -1 0 14990 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__13403_
timestamp 0
transform -1 0 12090 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13405_
timestamp 0
transform -1 0 13130 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__13408_
timestamp 0
transform 1 0 12550 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__13410_
timestamp 0
transform -1 0 12770 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__13413_
timestamp 0
transform -1 0 11810 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13415_
timestamp 0
transform -1 0 12310 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13417_
timestamp 0
transform 1 0 12450 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__13420_
timestamp 0
transform -1 0 11670 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13422_
timestamp 0
transform -1 0 12230 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__13425_
timestamp 0
transform -1 0 12610 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13427_
timestamp 0
transform -1 0 10830 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13503_
timestamp 0
transform -1 0 7530 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__13506_
timestamp 0
transform 1 0 8370 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__13508_
timestamp 0
transform 1 0 8450 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__13510_
timestamp 0
transform -1 0 7170 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__13513_
timestamp 0
transform 1 0 6390 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__13515_
timestamp 0
transform -1 0 7690 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__13518_
timestamp 0
transform 1 0 7950 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__13520_
timestamp 0
transform 1 0 8090 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__13522_
timestamp 0
transform 1 0 7830 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__13525_
timestamp 0
transform -1 0 7690 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__13527_
timestamp 0
transform 1 0 7590 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__13530_
timestamp 0
transform -1 0 8930 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__13532_
timestamp 0
transform -1 0 8750 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13534_
timestamp 0
transform -1 0 8770 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__13537_
timestamp 0
transform 1 0 8690 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__13539_
timestamp 0
transform -1 0 9230 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__13541_
timestamp 0
transform -1 0 8870 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__13544_
timestamp 0
transform -1 0 7170 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__13546_
timestamp 0
transform -1 0 7910 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13549_
timestamp 0
transform -1 0 9910 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13551_
timestamp 0
transform 1 0 10230 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__13553_
timestamp 0
transform -1 0 10050 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__13556_
timestamp 0
transform -1 0 8190 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__13558_
timestamp 0
transform 1 0 8150 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13560_
timestamp 0
transform 1 0 8310 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__13563_
timestamp 0
transform 1 0 7130 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__13565_
timestamp 0
transform 1 0 7310 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__13568_
timestamp 0
transform 1 0 9930 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__13570_
timestamp 0
transform 1 0 7270 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__13572_
timestamp 0
transform -1 0 6230 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13575_
timestamp 0
transform -1 0 9470 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__13577_
timestamp 0
transform -1 0 7450 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__13580_
timestamp 0
transform 1 0 8150 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__13582_
timestamp 0
transform 1 0 8310 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__13584_
timestamp 0
transform -1 0 7090 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__13587_
timestamp 0
transform -1 0 9410 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13589_
timestamp 0
transform -1 0 9650 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__13591_
timestamp 0
transform 1 0 9270 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__13594_
timestamp 0
transform 1 0 9330 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13596_
timestamp 0
transform 1 0 8910 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__13599_
timestamp 0
transform 1 0 7750 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13601_
timestamp 0
transform 1 0 6310 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13603_
timestamp 0
transform -1 0 9330 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__13606_
timestamp 0
transform 1 0 8830 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__13608_
timestamp 0
transform -1 0 7450 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__13611_
timestamp 0
transform -1 0 6170 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13613_
timestamp 0
transform 1 0 6250 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13615_
timestamp 0
transform 1 0 6310 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__13618_
timestamp 0
transform 1 0 9130 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__13620_
timestamp 0
transform 1 0 9250 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__13622_
timestamp 0
transform -1 0 6110 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13625_
timestamp 0
transform -1 0 8430 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__13627_
timestamp 0
transform 1 0 8230 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__13630_
timestamp 0
transform -1 0 5570 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13632_
timestamp 0
transform -1 0 6170 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13634_
timestamp 0
transform -1 0 5270 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13637_
timestamp 0
transform -1 0 4630 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13639_
timestamp 0
transform 1 0 5410 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13642_
timestamp 0
transform 1 0 6770 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13644_
timestamp 0
transform 1 0 6730 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__13646_
timestamp 0
transform -1 0 6690 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__13649_
timestamp 0
transform -1 0 5830 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13651_
timestamp 0
transform 1 0 9910 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__13653_
timestamp 0
transform 1 0 9970 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__13656_
timestamp 0
transform 1 0 7310 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13658_
timestamp 0
transform -1 0 7590 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13661_
timestamp 0
transform -1 0 5910 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13663_
timestamp 0
transform -1 0 5750 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13665_
timestamp 0
transform 1 0 5790 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13668_
timestamp 0
transform 1 0 4990 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13670_
timestamp 0
transform -1 0 5630 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13672_
timestamp 0
transform -1 0 5630 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13675_
timestamp 0
transform 1 0 9810 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13677_
timestamp 0
transform 1 0 9150 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13680_
timestamp 0
transform -1 0 7090 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__13682_
timestamp 0
transform -1 0 5990 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__13684_
timestamp 0
transform -1 0 6430 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__13687_
timestamp 0
transform -1 0 6030 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__13689_
timestamp 0
transform 1 0 6050 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__13692_
timestamp 0
transform -1 0 5990 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__13694_
timestamp 0
transform -1 0 7010 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13696_
timestamp 0
transform 1 0 9670 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13699_
timestamp 0
transform 1 0 7490 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13701_
timestamp 0
transform 1 0 6290 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13703_
timestamp 0
transform 1 0 6610 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13706_
timestamp 0
transform -1 0 6470 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13708_
timestamp 0
transform 1 0 6870 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__13711_
timestamp 0
transform 1 0 6510 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__13713_
timestamp 0
transform -1 0 5810 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13715_
timestamp 0
transform 1 0 6690 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__13718_
timestamp 0
transform 1 0 8190 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__13720_
timestamp 0
transform 1 0 7430 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__13723_
timestamp 0
transform -1 0 6390 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13725_
timestamp 0
transform 1 0 7030 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__13727_
timestamp 0
transform -1 0 6230 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13730_
timestamp 0
transform 1 0 6590 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__13732_
timestamp 0
transform -1 0 6070 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13734_
timestamp 0
transform 1 0 5910 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13737_
timestamp 0
transform 1 0 6190 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__13739_
timestamp 0
transform -1 0 6010 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13742_
timestamp 0
transform -1 0 7370 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13744_
timestamp 0
transform -1 0 9710 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__13746_
timestamp 0
transform -1 0 9570 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__13749_
timestamp 0
transform -1 0 7110 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13751_
timestamp 0
transform -1 0 6970 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13754_
timestamp 0
transform -1 0 6930 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__13756_
timestamp 0
transform -1 0 6770 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__13758_
timestamp 0
transform -1 0 6930 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__13761_
timestamp 0
transform -1 0 6910 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__13763_
timestamp 0
transform 1 0 6750 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__13765_
timestamp 0
transform -1 0 6970 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13768_
timestamp 0
transform 1 0 6470 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13770_
timestamp 0
transform 1 0 7910 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13773_
timestamp 0
transform -1 0 8090 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13775_
timestamp 0
transform -1 0 8070 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__13777_
timestamp 0
transform -1 0 8230 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__13780_
timestamp 0
transform 1 0 7530 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13782_
timestamp 0
transform -1 0 7150 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13784_
timestamp 0
transform -1 0 6910 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__13787_
timestamp 0
transform 1 0 6310 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__13789_
timestamp 0
transform 1 0 6490 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__13792_
timestamp 0
transform -1 0 8990 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__13794_
timestamp 0
transform -1 0 8570 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13796_
timestamp 0
transform -1 0 8410 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13799_
timestamp 0
transform -1 0 8110 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13801_
timestamp 0
transform -1 0 8770 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__13804_
timestamp 0
transform -1 0 7330 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__13806_
timestamp 0
transform -1 0 7330 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__13808_
timestamp 0
transform -1 0 9830 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13811_
timestamp 0
transform 1 0 9130 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__13813_
timestamp 0
transform 1 0 9230 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13815_
timestamp 0
transform -1 0 8950 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13818_
timestamp 0
transform 1 0 9370 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13820_
timestamp 0
transform 1 0 9090 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__13823_
timestamp 0
transform 1 0 7930 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13825_
timestamp 0
transform 1 0 8250 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__13827_
timestamp 0
transform 1 0 7950 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__13830_
timestamp 0
transform -1 0 7650 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__13832_
timestamp 0
transform -1 0 7370 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13835_
timestamp 0
transform 1 0 10450 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__13837_
timestamp 0
transform -1 0 9990 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__13839_
timestamp 0
transform -1 0 9490 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__13842_
timestamp 0
transform -1 0 8030 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__13844_
timestamp 0
transform 1 0 8190 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__13846_
timestamp 0
transform -1 0 7490 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__13849_
timestamp 0
transform -1 0 5830 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13851_
timestamp 0
transform -1 0 5950 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13854_
timestamp 0
transform 1 0 7010 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13856_
timestamp 0
transform -1 0 6750 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13858_
timestamp 0
transform -1 0 7930 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__13861_
timestamp 0
transform -1 0 7950 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__13863_
timestamp 0
transform 1 0 7830 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13866_
timestamp 0
transform 1 0 7930 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13868_
timestamp 0
transform 1 0 7670 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13870_
timestamp 0
transform 1 0 8670 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__13873_
timestamp 0
transform 1 0 5510 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13875_
timestamp 0
transform -1 0 6290 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13877_
timestamp 0
transform -1 0 6570 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13880_
timestamp 0
transform 1 0 7630 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13882_
timestamp 0
transform 1 0 7550 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__13885_
timestamp 0
transform -1 0 7030 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13887_
timestamp 0
transform -1 0 8130 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13889_
timestamp 0
transform 1 0 7210 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13892_
timestamp 0
transform 1 0 8790 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13894_
timestamp 0
transform -1 0 8650 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13896_
timestamp 0
transform -1 0 8090 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13899_
timestamp 0
transform -1 0 7530 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__13901_
timestamp 0
transform 1 0 8430 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13904_
timestamp 0
transform -1 0 8810 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__13906_
timestamp 0
transform -1 0 6230 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13908_
timestamp 0
transform 1 0 6470 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13911_
timestamp 0
transform 1 0 8670 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13913_
timestamp 0
transform 1 0 8910 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13916_
timestamp 0
transform -1 0 8910 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13918_
timestamp 0
transform -1 0 8490 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__13920_
timestamp 0
transform 1 0 8750 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__13923_
timestamp 0
transform -1 0 7150 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13925_
timestamp 0
transform -1 0 9670 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__13927_
timestamp 0
transform 1 0 9430 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__13930_
timestamp 0
transform 1 0 7790 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13932_
timestamp 0
transform 1 0 8830 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13935_
timestamp 0
transform -1 0 7930 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13937_
timestamp 0
transform -1 0 7770 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13939_
timestamp 0
transform -1 0 6750 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13942_
timestamp 0
transform -1 0 8150 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__13944_
timestamp 0
transform 1 0 10310 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__13947_
timestamp 0
transform 1 0 10450 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__13949_
timestamp 0
transform 1 0 10510 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__13951_
timestamp 0
transform 1 0 8270 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13954_
timestamp 0
transform 1 0 9390 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13956_
timestamp 0
transform -1 0 10150 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13958_
timestamp 0
transform 1 0 10430 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13961_
timestamp 0
transform -1 0 8090 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13963_
timestamp 0
transform -1 0 9150 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13966_
timestamp 0
transform 1 0 9630 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13968_
timestamp 0
transform 1 0 10230 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13970_
timestamp 0
transform -1 0 9150 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__13973_
timestamp 0
transform -1 0 8570 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13975_
timestamp 0
transform 1 0 9210 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__13978_
timestamp 0
transform -1 0 8250 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13980_
timestamp 0
transform 1 0 8390 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2__13982_
timestamp 0
transform -1 0 9630 0 1 16090
box -6 -8 26 248
use FILL  FILL_2__13985_
timestamp 0
transform 1 0 9210 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__13987_
timestamp 0
transform 1 0 10330 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__13989_
timestamp 0
transform 1 0 10510 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__13992_
timestamp 0
transform 1 0 9990 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2__13994_
timestamp 0
transform 1 0 10690 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__13997_
timestamp 0
transform -1 0 10510 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__13999_
timestamp 0
transform -1 0 10470 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__14001_
timestamp 0
transform 1 0 9810 0 1 16570
box -6 -8 26 248
use FILL  FILL_2__14004_
timestamp 0
transform -1 0 10290 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__14006_
timestamp 0
transform -1 0 10170 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2__14009_
timestamp 0
transform -1 0 9970 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__14011_
timestamp 0
transform -1 0 9670 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__14013_
timestamp 0
transform -1 0 8690 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__14016_
timestamp 0
transform 1 0 10730 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__14018_
timestamp 0
transform 1 0 10870 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__14020_
timestamp 0
transform -1 0 10830 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__14023_
timestamp 0
transform -1 0 10570 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__14025_
timestamp 0
transform 1 0 11250 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__14028_
timestamp 0
transform -1 0 9450 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__14030_
timestamp 0
transform 1 0 10210 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__14032_
timestamp 0
transform 1 0 8930 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__14035_
timestamp 0
transform 1 0 10090 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__14037_
timestamp 0
transform -1 0 10670 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__14039_
timestamp 0
transform 1 0 10630 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__14042_
timestamp 0
transform 1 0 11030 0 1 14650
box -6 -8 26 248
use FILL  FILL_2__14044_
timestamp 0
transform -1 0 10910 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__14047_
timestamp 0
transform -1 0 10470 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__14049_
timestamp 0
transform 1 0 9990 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__14051_
timestamp 0
transform -1 0 9550 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__14054_
timestamp 0
transform 1 0 9690 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__14056_
timestamp 0
transform 1 0 10470 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__14059_
timestamp 0
transform -1 0 9950 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__14061_
timestamp 0
transform 1 0 10290 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__14063_
timestamp 0
transform 1 0 10030 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2__14066_
timestamp 0
transform -1 0 10330 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__14068_
timestamp 0
transform 1 0 9370 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__14070_
timestamp 0
transform -1 0 10630 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__14073_
timestamp 0
transform 1 0 10570 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__14075_
timestamp 0
transform 1 0 10490 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__14078_
timestamp 0
transform 1 0 10130 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__14080_
timestamp 0
transform -1 0 9690 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__14082_
timestamp 0
transform -1 0 9270 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__14085_
timestamp 0
transform -1 0 10090 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__14087_
timestamp 0
transform -1 0 9950 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__14090_
timestamp 0
transform 1 0 11090 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2__14092_
timestamp 0
transform 1 0 10070 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__14094_
timestamp 0
transform -1 0 9930 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__14097_
timestamp 0
transform -1 0 9790 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__14099_
timestamp 0
transform 1 0 8790 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__14101_
timestamp 0
transform 1 0 8790 0 1 12730
box -6 -8 26 248
use FILL  FILL_2__14104_
timestamp 0
transform -1 0 9710 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__14106_
timestamp 0
transform -1 0 9590 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__14109_
timestamp 0
transform 1 0 9750 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__14111_
timestamp 0
transform 1 0 9350 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__14113_
timestamp 0
transform 1 0 7610 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__14116_
timestamp 0
transform -1 0 9610 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2__14118_
timestamp 0
transform -1 0 7890 0 1 12250
box -6 -8 26 248
use FILL  FILL_2__14121_
timestamp 0
transform 1 0 9870 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__14123_
timestamp 0
transform -1 0 8450 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__14125_
timestamp 0
transform 1 0 8130 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__14128_
timestamp 0
transform -1 0 8530 0 1 15130
box -6 -8 26 248
use FILL  FILL_2__14130_
timestamp 0
transform 1 0 9030 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2__14132_
timestamp 0
transform 1 0 10170 0 1 13690
box -6 -8 26 248
use FILL  FILL_2__14135_
timestamp 0
transform -1 0 8470 0 1 14170
box -6 -8 26 248
use FILL  FILL_2__14137_
timestamp 0
transform 1 0 9050 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__14140_
timestamp 0
transform 1 0 8910 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2__14142_
timestamp 0
transform 1 0 7650 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__14144_
timestamp 0
transform -1 0 7830 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2__14147_
timestamp 0
transform 1 0 7570 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2__14149_
timestamp 0
transform -1 0 7490 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2__14151_
timestamp 0
transform -1 0 7630 0 1 13210
box -6 -8 26 248
use FILL  FILL_2__14154_
timestamp 0
transform -1 0 6990 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__14156_
timestamp 0
transform 1 0 7270 0 1 15610
box -6 -8 26 248
use FILL  FILL_2__14216_
timestamp 0
transform 1 0 7490 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__14218_
timestamp 0
transform -1 0 7730 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__14220_
timestamp 0
transform 1 0 7670 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__14223_
timestamp 0
transform -1 0 6930 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__14225_
timestamp 0
transform 1 0 6850 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__14228_
timestamp 0
transform -1 0 8550 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__14230_
timestamp 0
transform -1 0 8390 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__14232_
timestamp 0
transform -1 0 9970 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__14235_
timestamp 0
transform 1 0 8550 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__14237_
timestamp 0
transform -1 0 8890 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__14239_
timestamp 0
transform -1 0 8030 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__14242_
timestamp 0
transform -1 0 8310 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__14244_
timestamp 0
transform 1 0 6910 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__14247_
timestamp 0
transform 1 0 8730 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__14249_
timestamp 0
transform 1 0 9830 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__14251_
timestamp 0
transform 1 0 9850 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__14254_
timestamp 0
transform 1 0 7670 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__14256_
timestamp 0
transform 1 0 7170 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__14259_
timestamp 0
transform -1 0 7190 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__14261_
timestamp 0
transform 1 0 7750 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__14263_
timestamp 0
transform -1 0 7830 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__14266_
timestamp 0
transform -1 0 6950 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__14268_
timestamp 0
transform -1 0 6910 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__14270_
timestamp 0
transform 1 0 6930 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__14273_
timestamp 0
transform 1 0 7570 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__14275_
timestamp 0
transform 1 0 7290 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__14278_
timestamp 0
transform -1 0 7990 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__14280_
timestamp 0
transform -1 0 9270 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__14282_
timestamp 0
transform -1 0 9390 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__14285_
timestamp 0
transform -1 0 8430 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__14287_
timestamp 0
transform -1 0 9190 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__14290_
timestamp 0
transform 1 0 7950 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__14292_
timestamp 0
transform -1 0 8210 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__14294_
timestamp 0
transform -1 0 9250 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__14297_
timestamp 0
transform 1 0 9090 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__14299_
timestamp 0
transform -1 0 8850 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__14301_
timestamp 0
transform 1 0 7850 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__14304_
timestamp 0
transform -1 0 9010 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__14306_
timestamp 0
transform -1 0 8850 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__14309_
timestamp 0
transform 1 0 9390 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__14311_
timestamp 0
transform -1 0 8370 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__14313_
timestamp 0
transform -1 0 9670 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__14316_
timestamp 0
transform 1 0 8690 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__14318_
timestamp 0
transform 1 0 8450 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__14320_
timestamp 0
transform -1 0 9730 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__14323_
timestamp 0
transform 1 0 8570 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__14325_
timestamp 0
transform 1 0 8450 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__14328_
timestamp 0
transform 1 0 8870 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__14330_
timestamp 0
transform 1 0 9030 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__14332_
timestamp 0
transform -1 0 9310 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__14335_
timestamp 0
transform -1 0 8670 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__14337_
timestamp 0
transform -1 0 8430 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__14340_
timestamp 0
transform -1 0 9030 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__14342_
timestamp 0
transform 1 0 9150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__14344_
timestamp 0
transform 1 0 8990 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__14347_
timestamp 0
transform -1 0 9590 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__14349_
timestamp 0
transform 1 0 7870 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__14351_
timestamp 0
transform -1 0 7710 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__14354_
timestamp 0
transform -1 0 8030 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__14356_
timestamp 0
transform 1 0 8310 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__14359_
timestamp 0
transform 1 0 8450 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__14361_
timestamp 0
transform 1 0 8470 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__14363_
timestamp 0
transform 1 0 8150 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__14366_
timestamp 0
transform 1 0 8050 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__14368_
timestamp 0
transform -1 0 9430 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__14371_
timestamp 0
transform -1 0 9670 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__14373_
timestamp 0
transform 1 0 8690 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__14375_
timestamp 0
transform 1 0 10390 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__14378_
timestamp 0
transform 1 0 10970 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__14380_
timestamp 0
transform -1 0 11150 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__14382_
timestamp 0
transform 1 0 9530 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__14385_
timestamp 0
transform 1 0 10730 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__14387_
timestamp 0
transform 1 0 10650 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__14390_
timestamp 0
transform -1 0 10350 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__14392_
timestamp 0
transform 1 0 10630 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__14394_
timestamp 0
transform -1 0 10930 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__14397_
timestamp 0
transform 1 0 9790 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__14399_
timestamp 0
transform 1 0 10590 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__14402_
timestamp 0
transform 1 0 10090 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__14404_
timestamp 0
transform -1 0 8970 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__14406_
timestamp 0
transform 1 0 10270 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__14409_
timestamp 0
transform -1 0 9030 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__14411_
timestamp 0
transform -1 0 10450 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__14413_
timestamp 0
transform 1 0 10270 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__14416_
timestamp 0
transform 1 0 9870 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__14418_
timestamp 0
transform -1 0 9270 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__14421_
timestamp 0
transform -1 0 8190 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__14423_
timestamp 0
transform 1 0 8990 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__14425_
timestamp 0
transform 1 0 9610 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__14428_
timestamp 0
transform -1 0 10070 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__14430_
timestamp 0
transform 1 0 9810 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__14433_
timestamp 0
transform 1 0 8050 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__14435_
timestamp 0
transform 1 0 8510 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__14437_
timestamp 0
transform -1 0 8150 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__14440_
timestamp 0
transform 1 0 9150 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__14442_
timestamp 0
transform 1 0 8330 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__14444_
timestamp 0
transform 1 0 9030 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__14447_
timestamp 0
transform 1 0 8670 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__14449_
timestamp 0
transform 1 0 8030 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__14452_
timestamp 0
transform 1 0 8890 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__14454_
timestamp 0
transform 1 0 8150 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__14456_
timestamp 0
transform 1 0 8570 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__14459_
timestamp 0
transform 1 0 8150 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__14461_
timestamp 0
transform 1 0 8190 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__14463_
timestamp 0
transform 1 0 8230 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__14466_
timestamp 0
transform -1 0 7750 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__14468_
timestamp 0
transform 1 0 7910 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__14471_
timestamp 0
transform 1 0 7170 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__14473_
timestamp 0
transform 1 0 9210 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__14475_
timestamp 0
transform -1 0 8030 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__14478_
timestamp 0
transform -1 0 9270 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__14480_
timestamp 0
transform 1 0 9730 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__14483_
timestamp 0
transform 1 0 9830 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__14485_
timestamp 0
transform 1 0 9530 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__14487_
timestamp 0
transform 1 0 9890 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__14490_
timestamp 0
transform 1 0 8410 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__14492_
timestamp 0
transform 1 0 8250 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__14494_
timestamp 0
transform -1 0 7510 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__14497_
timestamp 0
transform -1 0 7350 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__14499_
timestamp 0
transform -1 0 9590 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__14558_
timestamp 0
transform -1 0 14070 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__14560_
timestamp 0
transform -1 0 12170 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__14562_
timestamp 0
transform 1 0 11730 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__14565_
timestamp 0
transform -1 0 12670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__14567_
timestamp 0
transform -1 0 14610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__14570_
timestamp 0
transform 1 0 15070 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__14572_
timestamp 0
transform -1 0 14150 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__14574_
timestamp 0
transform 1 0 11670 0 1 730
box -6 -8 26 248
use FILL  FILL_2__14577_
timestamp 0
transform -1 0 13190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__14579_
timestamp 0
transform -1 0 13430 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__14581_
timestamp 0
transform 1 0 14350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__14584_
timestamp 0
transform -1 0 13950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__14586_
timestamp 0
transform -1 0 9770 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14589_
timestamp 0
transform -1 0 9930 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14591_
timestamp 0
transform -1 0 12010 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__14593_
timestamp 0
transform 1 0 13050 0 1 730
box -6 -8 26 248
use FILL  FILL_2__14596_
timestamp 0
transform 1 0 14290 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__14598_
timestamp 0
transform 1 0 13810 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__14601_
timestamp 0
transform -1 0 11870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__14603_
timestamp 0
transform 1 0 15330 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__14605_
timestamp 0
transform -1 0 15050 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__14608_
timestamp 0
transform -1 0 14870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__14610_
timestamp 0
transform -1 0 15790 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__14612_
timestamp 0
transform 1 0 16190 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__14615_
timestamp 0
transform 1 0 15210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__14617_
timestamp 0
transform -1 0 14710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__14620_
timestamp 0
transform 1 0 14350 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__14622_
timestamp 0
transform 1 0 13930 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__14624_
timestamp 0
transform -1 0 13810 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__14627_
timestamp 0
transform 1 0 14690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__14629_
timestamp 0
transform 1 0 14430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__14631_
timestamp 0
transform -1 0 14170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__14634_
timestamp 0
transform -1 0 13750 0 1 730
box -6 -8 26 248
use FILL  FILL_2__14636_
timestamp 0
transform 1 0 14630 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__14639_
timestamp 0
transform 1 0 15530 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__14641_
timestamp 0
transform -1 0 15710 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__14643_
timestamp 0
transform 1 0 15850 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__14646_
timestamp 0
transform -1 0 15630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__14648_
timestamp 0
transform 1 0 16150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__14651_
timestamp 0
transform 1 0 16970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__14653_
timestamp 0
transform 1 0 16430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__14655_
timestamp 0
transform -1 0 16830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__14658_
timestamp 0
transform 1 0 16690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__14660_
timestamp 0
transform 1 0 16110 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__14662_
timestamp 0
transform -1 0 16910 0 1 730
box -6 -8 26 248
use FILL  FILL_2__14665_
timestamp 0
transform 1 0 17050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__14667_
timestamp 0
transform 1 0 17030 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14670_
timestamp 0
transform -1 0 16650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__14672_
timestamp 0
transform -1 0 16750 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14674_
timestamp 0
transform -1 0 16370 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14677_
timestamp 0
transform -1 0 15990 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14679_
timestamp 0
transform 1 0 16270 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14682_
timestamp 0
transform -1 0 15970 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14684_
timestamp 0
transform -1 0 16590 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14686_
timestamp 0
transform -1 0 16810 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__14689_
timestamp 0
transform 1 0 16370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__14691_
timestamp 0
transform -1 0 15830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__14693_
timestamp 0
transform 1 0 14470 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14696_
timestamp 0
transform 1 0 14690 0 1 730
box -6 -8 26 248
use FILL  FILL_2__14698_
timestamp 0
transform -1 0 14870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__14701_
timestamp 0
transform 1 0 14850 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14703_
timestamp 0
transform -1 0 14330 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14705_
timestamp 0
transform 1 0 14990 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14708_
timestamp 0
transform -1 0 13990 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14710_
timestamp 0
transform 1 0 14170 0 1 730
box -6 -8 26 248
use FILL  FILL_2__14713_
timestamp 0
transform 1 0 15270 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14715_
timestamp 0
transform 1 0 15150 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14717_
timestamp 0
transform 1 0 15690 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14720_
timestamp 0
transform 1 0 15550 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14722_
timestamp 0
transform 1 0 15470 0 1 730
box -6 -8 26 248
use FILL  FILL_2__14724_
timestamp 0
transform -1 0 15850 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14727_
timestamp 0
transform 1 0 15810 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14729_
timestamp 0
transform 1 0 16110 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14732_
timestamp 0
transform 1 0 16010 0 1 730
box -6 -8 26 248
use FILL  FILL_2__14734_
timestamp 0
transform 1 0 12770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__14736_
timestamp 0
transform -1 0 15410 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14739_
timestamp 0
transform -1 0 15190 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14741_
timestamp 0
transform 1 0 14690 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14743_
timestamp 0
transform -1 0 12050 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14746_
timestamp 0
transform -1 0 12590 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14748_
timestamp 0
transform -1 0 12630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__14751_
timestamp 0
transform -1 0 11270 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14753_
timestamp 0
transform 1 0 12310 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14755_
timestamp 0
transform 1 0 12250 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14758_
timestamp 0
transform 1 0 12730 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14760_
timestamp 0
transform -1 0 11530 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14763_
timestamp 0
transform -1 0 12330 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14765_
timestamp 0
transform 1 0 13430 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14767_
timestamp 0
transform 1 0 13010 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14770_
timestamp 0
transform 1 0 12870 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14772_
timestamp 0
transform 1 0 13490 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14774_
timestamp 0
transform -1 0 13750 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14777_
timestamp 0
transform 1 0 13990 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14779_
timestamp 0
transform -1 0 13230 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14782_
timestamp 0
transform 1 0 13010 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14784_
timestamp 0
transform -1 0 14410 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14786_
timestamp 0
transform 1 0 13590 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14789_
timestamp 0
transform 1 0 13430 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14791_
timestamp 0
transform 1 0 13990 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14794_
timestamp 0
transform 1 0 11110 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14796_
timestamp 0
transform 1 0 11630 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14798_
timestamp 0
transform 1 0 16090 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__14801_
timestamp 0
transform 1 0 14550 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14803_
timestamp 0
transform -1 0 14170 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14805_
timestamp 0
transform 1 0 11890 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14808_
timestamp 0
transform -1 0 11690 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14810_
timestamp 0
transform 1 0 10810 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14813_
timestamp 0
transform 1 0 11350 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14815_
timestamp 0
transform -1 0 11110 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14817_
timestamp 0
transform -1 0 11090 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14820_
timestamp 0
transform -1 0 10290 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14822_
timestamp 0
transform 1 0 10390 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14825_
timestamp 0
transform -1 0 10230 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14827_
timestamp 0
transform -1 0 10070 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14829_
timestamp 0
transform -1 0 10130 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14832_
timestamp 0
transform -1 0 10930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__14834_
timestamp 0
transform -1 0 9550 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14836_
timestamp 0
transform -1 0 9150 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__14839_
timestamp 0
transform 1 0 10530 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14841_
timestamp 0
transform 1 0 10250 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14844_
timestamp 0
transform -1 0 12270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__14846_
timestamp 0
transform 1 0 12390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__14848_
timestamp 0
transform -1 0 13490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__14851_
timestamp 0
transform 1 0 15470 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__14853_
timestamp 0
transform -1 0 13350 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__14855_
timestamp 0
transform 1 0 14410 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__14858_
timestamp 0
transform 1 0 13050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__14860_
timestamp 0
transform -1 0 13510 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__14863_
timestamp 0
transform 1 0 12170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__14865_
timestamp 0
transform -1 0 10950 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__14867_
timestamp 0
transform 1 0 11030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__14909_
timestamp 0
transform -1 0 70 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__14911_
timestamp 0
transform -1 0 9790 0 1 250
box -6 -8 26 248
use FILL  FILL_2__14914_
timestamp 0
transform 1 0 8250 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__14916_
timestamp 0
transform 1 0 8450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__14918_
timestamp 0
transform -1 0 8130 0 1 6010
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert1
timestamp 0
transform 1 0 9510 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert3
timestamp 0
transform 1 0 9470 0 1 8410
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert5
timestamp 0
transform 1 0 5430 0 1 9370
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert8
timestamp 0
transform -1 0 1190 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert10
timestamp 0
transform 1 0 4150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert13
timestamp 0
transform -1 0 4450 0 1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert15
timestamp 0
transform 1 0 6870 0 1 7930
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert17
timestamp 0
transform -1 0 3250 0 1 7450
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert20
timestamp 0
transform -1 0 16290 0 1 7930
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert22
timestamp 0
transform -1 0 12130 0 1 7930
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert25
timestamp 0
transform 1 0 1070 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert27
timestamp 0
transform -1 0 1210 0 1 10810
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert108
timestamp 0
transform -1 0 7830 0 1 7450
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert110
timestamp 0
transform -1 0 9050 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert113
timestamp 0
transform -1 0 13870 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert115
timestamp 0
transform -1 0 14370 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert117
timestamp 0
transform -1 0 6990 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert120
timestamp 0
transform 1 0 7110 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert122
timestamp 0
transform -1 0 7610 0 1 6010
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert125
timestamp 0
transform -1 0 6030 0 1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert127
timestamp 0
transform -1 0 4110 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert129
timestamp 0
transform -1 0 4210 0 1 7450
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert132
timestamp 0
transform 1 0 2690 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert134
timestamp 0
transform -1 0 450 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert137
timestamp 0
transform -1 0 11930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert139
timestamp 0
transform 1 0 15530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert141
timestamp 0
transform -1 0 10990 0 1 11290
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert144
timestamp 0
transform 1 0 12210 0 1 11290
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert146
timestamp 0
transform -1 0 10550 0 1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert148
timestamp 0
transform 1 0 8510 0 1 250
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert151
timestamp 0
transform -1 0 16090 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert153
timestamp 0
transform -1 0 15950 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert156
timestamp 0
transform -1 0 15750 0 1 9370
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert158
timestamp 0
transform 1 0 16970 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert160
timestamp 0
transform 1 0 16430 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert163
timestamp 0
transform 1 0 12750 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert165
timestamp 0
transform -1 0 11710 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert167
timestamp 0
transform -1 0 1170 0 1 9370
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert170
timestamp 0
transform 1 0 1530 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert172
timestamp 0
transform 1 0 12870 0 1 12730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert175
timestamp 0
transform 1 0 14770 0 1 12250
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert177
timestamp 0
transform 1 0 15870 0 1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert179
timestamp 0
transform 1 0 15850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert182
timestamp 0
transform -1 0 10070 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert184
timestamp 0
transform 1 0 11830 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert187
timestamp 0
transform 1 0 8250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert189
timestamp 0
transform -1 0 5990 0 1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert191
timestamp 0
transform 1 0 12530 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert194
timestamp 0
transform -1 0 11450 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert196
timestamp 0
transform -1 0 1410 0 1 5050
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert198
timestamp 0
transform -1 0 750 0 1 5050
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert201
timestamp 0
transform -1 0 11910 0 1 10810
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert203
timestamp 0
transform -1 0 12630 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert206
timestamp 0
transform 1 0 14050 0 1 5050
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert208
timestamp 0
transform 1 0 15510 0 1 5050
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert210
timestamp 0
transform 1 0 1150 0 1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert213
timestamp 0
transform -1 0 70 0 1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert215
timestamp 0
transform -1 0 5750 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert218
timestamp 0
transform 1 0 6710 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert220
timestamp 0
transform 1 0 11770 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert222
timestamp 0
transform -1 0 9990 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert225
timestamp 0
transform 1 0 6970 0 -1 16570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert227
timestamp 0
transform -1 0 6870 0 1 15130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert229
timestamp 0
transform 1 0 8990 0 -1 15130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert232
timestamp 0
transform -1 0 8950 0 1 15130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert234
timestamp 0
transform 1 0 15390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert237
timestamp 0
transform -1 0 13250 0 1 730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert239
timestamp 0
transform -1 0 4690 0 1 13210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert241
timestamp 0
transform 1 0 5650 0 -1 14170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert244
timestamp 0
transform -1 0 1430 0 1 4570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert246
timestamp 0
transform 1 0 2450 0 1 4570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert249
timestamp 0
transform 1 0 3270 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert251
timestamp 0
transform -1 0 1930 0 -1 15610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert253
timestamp 0
transform 1 0 8650 0 1 6010
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert256
timestamp 0
transform 1 0 11130 0 1 4570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert258
timestamp 0
transform -1 0 14010 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert260
timestamp 0
transform 1 0 16490 0 1 15610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert263
timestamp 0
transform -1 0 13370 0 1 13690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert265
timestamp 0
transform 1 0 5450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert268
timestamp 0
transform -1 0 4390 0 1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert270
timestamp 0
transform -1 0 7210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert272
timestamp 0
transform 1 0 8090 0 1 1690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert275
timestamp 0
transform 1 0 9890 0 1 730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert277
timestamp 0
transform -1 0 7050 0 1 730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert279
timestamp 0
transform 1 0 9930 0 1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert282
timestamp 0
transform 1 0 15930 0 1 13690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert284
timestamp 0
transform 1 0 16110 0 -1 13210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert287
timestamp 0
transform 1 0 16390 0 1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert289
timestamp 0
transform -1 0 13030 0 1 9370
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert291
timestamp 0
transform 1 0 6610 0 1 12730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert294
timestamp 0
transform -1 0 11890 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert296
timestamp 0
transform 1 0 15250 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert299
timestamp 0
transform 1 0 16930 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert301
timestamp 0
transform -1 0 8010 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert303
timestamp 0
transform -1 0 8070 0 1 12730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert306
timestamp 0
transform -1 0 9710 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert308
timestamp 0
transform 1 0 10230 0 1 7930
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert310
timestamp 0
transform 1 0 13770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert313
timestamp 0
transform -1 0 15110 0 1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert315
timestamp 0
transform 1 0 16410 0 1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert318
timestamp 0
transform -1 0 11710 0 1 5530
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert320
timestamp 0
transform 1 0 8590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert322
timestamp 0
transform 1 0 7050 0 1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert325
timestamp 0
transform 1 0 2990 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert327
timestamp 0
transform -1 0 2910 0 1 15130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert330
timestamp 0
transform -1 0 2870 0 1 15610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert332
timestamp 0
transform -1 0 2850 0 1 12730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert334
timestamp 0
transform 1 0 2830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert337
timestamp 0
transform -1 0 1190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert339
timestamp 0
transform -1 0 830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert341
timestamp 0
transform -1 0 570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert344
timestamp 0
transform -1 0 70 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert346
timestamp 0
transform -1 0 11090 0 -1 13690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert349
timestamp 0
transform 1 0 8110 0 -1 16090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert351
timestamp 0
transform -1 0 7650 0 1 15130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert353
timestamp 0
transform 1 0 10750 0 -1 14650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert356
timestamp 0
transform 1 0 9470 0 1 16090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert358
timestamp 0
transform 1 0 10790 0 1 13690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert361
timestamp 0
transform -1 0 6330 0 1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert363
timestamp 0
transform 1 0 6690 0 1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert365
timestamp 0
transform -1 0 4830 0 1 13210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert368
timestamp 0
transform -1 0 4770 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert370
timestamp 0
transform -1 0 12930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert372
timestamp 0
transform 1 0 13210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert375
timestamp 0
transform 1 0 3010 0 1 9370
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert377
timestamp 0
transform -1 0 2010 0 1 9370
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert380
timestamp 0
transform 1 0 4950 0 1 13210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert382
timestamp 0
transform 1 0 5770 0 1 11290
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert29
timestamp 0
transform -1 0 9430 0 1 4570
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert32
timestamp 0
transform -1 0 6230 0 1 12250
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert34
timestamp 0
transform -1 0 10070 0 1 7450
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert36
timestamp 0
transform 1 0 3530 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert39
timestamp 0
transform -1 0 5890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert41
timestamp 0
transform -1 0 11330 0 1 3130
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert44
timestamp 0
transform 1 0 2770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert46
timestamp 0
transform 1 0 3510 0 1 6490
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert48
timestamp 0
transform -1 0 2110 0 -1 12730
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert51
timestamp 0
transform 1 0 14730 0 1 13690
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert53
timestamp 0
transform -1 0 4270 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert55
timestamp 0
transform 1 0 14170 0 1 12730
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert58
timestamp 0
transform 1 0 7170 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert60
timestamp 0
transform -1 0 8870 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert63
timestamp 0
transform 1 0 10350 0 1 12250
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert65
timestamp 0
transform 1 0 6950 0 1 2170
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert67
timestamp 0
transform -1 0 15230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert70
timestamp 0
transform 1 0 3050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert72
timestamp 0
transform 1 0 9430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert75
timestamp 0
transform 1 0 10350 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert77
timestamp 0
transform 1 0 11430 0 1 7930
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert79
timestamp 0
transform 1 0 11390 0 1 4570
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert82
timestamp 0
transform 1 0 11970 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert84
timestamp 0
transform 1 0 8470 0 1 11290
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert86
timestamp 0
transform 1 0 12610 0 1 3130
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert89
timestamp 0
transform 1 0 6530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert91
timestamp 0
transform -1 0 2150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert94
timestamp 0
transform -1 0 4130 0 1 4090
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert96
timestamp 0
transform -1 0 9010 0 1 5050
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert98
timestamp 0
transform -1 0 8130 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert101
timestamp 0
transform -1 0 14950 0 -1 12250
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert103
timestamp 0
transform -1 0 10150 0 1 6970
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert106
timestamp 0
transform -1 0 2210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert384
timestamp 0
transform 1 0 8930 0 -1 17050
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert387
timestamp 0
transform 1 0 10790 0 1 7450
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert389
timestamp 0
transform 1 0 8390 0 1 6010
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert391
timestamp 0
transform -1 0 7050 0 1 10810
box -6 -8 26 248
<< labels >>
flabel metal1 s 17202 2 17262 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -62 2 -2 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 9817 -23 9823 -17 7 FreeSans 16 270 0 0 Dout[11]
port 2 nsew
flabel metal2 s 8537 -23 8543 -17 7 FreeSans 16 270 0 0 Dout[10]
port 3 nsew
flabel metal3 s -24 7556 -16 7564 7 FreeSans 16 0 0 0 Dout[9]
port 4 nsew
flabel metal2 s 8117 -23 8123 -17 7 FreeSans 16 270 0 0 Dout[8]
port 5 nsew
flabel metal2 s 7997 -23 8003 -17 7 FreeSans 16 270 0 0 Dout[7]
port 6 nsew
flabel metal2 s 8497 -23 8503 -17 7 FreeSans 16 270 0 0 Dout[6]
port 7 nsew
flabel metal3 s 17236 116 17244 124 3 FreeSans 16 0 0 0 Dout[5]
port 8 nsew
flabel metal2 s 8297 -23 8303 -17 7 FreeSans 16 270 0 0 Dout[4]
port 9 nsew
flabel metal3 s -24 7056 -16 7064 7 FreeSans 16 0 0 0 Dout[3]
port 10 nsew
flabel metal3 s -24 7096 -16 7104 7 FreeSans 16 0 0 0 Dout[2]
port 11 nsew
flabel metal3 s -24 8036 -16 8044 7 FreeSans 16 0 0 0 Dout[1]
port 12 nsew
flabel metal2 s 7637 -23 7643 -17 7 FreeSans 16 270 0 0 Dout[0]
port 13 nsew
flabel metal2 s 12097 -23 12103 -17 7 FreeSans 16 270 0 0 En
port 14 nsew
flabel metal2 s 9177 -23 9183 -17 7 FreeSans 16 270 0 0 FCW[19]
port 15 nsew
flabel metal2 s 10317 -23 10323 -17 7 FreeSans 16 270 0 0 FCW[18]
port 16 nsew
flabel metal2 s 10717 -23 10723 -17 7 FreeSans 16 270 0 0 FCW[17]
port 17 nsew
flabel metal2 s 11137 -23 11143 -17 7 FreeSans 16 270 0 0 FCW[16]
port 18 nsew
flabel metal2 s 13897 -23 13903 -17 7 FreeSans 16 270 0 0 FCW[15]
port 19 nsew
flabel metal2 s 12357 -23 12363 -17 7 FreeSans 16 270 0 0 FCW[14]
port 20 nsew
flabel metal2 s 11317 -23 11323 -17 7 FreeSans 16 270 0 0 FCW[13]
port 21 nsew
flabel metal2 s 12177 -23 12183 -17 7 FreeSans 16 270 0 0 FCW[12]
port 22 nsew
flabel metal2 s 15837 -23 15843 -17 7 FreeSans 16 270 0 0 FCW[11]
port 23 nsew
flabel metal2 s 15677 -23 15683 -17 7 FreeSans 16 270 0 0 FCW[10]
port 24 nsew
flabel metal2 s 14717 -23 14723 -17 7 FreeSans 16 270 0 0 FCW[9]
port 25 nsew
flabel metal2 s 14417 -23 14423 -17 7 FreeSans 16 270 0 0 FCW[8]
port 26 nsew
flabel metal2 s 16137 -23 16143 -17 7 FreeSans 16 270 0 0 FCW[7]
port 27 nsew
flabel metal2 s 16977 -23 16983 -17 7 FreeSans 16 270 0 0 FCW[6]
port 28 nsew
flabel metal3 s 17236 1796 17244 1804 3 FreeSans 16 0 0 0 FCW[5]
port 29 nsew
flabel metal2 s 15457 -23 15463 -17 7 FreeSans 16 270 0 0 FCW[4]
port 30 nsew
flabel metal2 s 14637 -23 14643 -17 7 FreeSans 16 270 0 0 FCW[3]
port 31 nsew
flabel metal2 s 13657 -23 13663 -17 7 FreeSans 16 270 0 0 FCW[2]
port 32 nsew
flabel metal2 s 15017 -23 15023 -17 7 FreeSans 16 270 0 0 FCW[1]
port 33 nsew
flabel metal2 s 14677 -23 14683 -17 7 FreeSans 16 270 0 0 FCW[0]
port 34 nsew
flabel metal2 s 9037 -23 9043 -17 7 FreeSans 16 270 0 0 Vld
port 35 nsew
flabel metal2 s 8957 17097 8963 17103 3 FreeSans 16 90 0 0 clk
port 36 nsew
flabel metal2 s 8317 17097 8323 17103 3 FreeSans 16 90 0 0 selSign
port 37 nsew
flabel metal2 s 8157 -23 8163 -17 7 FreeSans 16 270 0 0 selXY
port 38 nsew
<< properties >>
string FIXED_BBOX -40 -40 17240 17100
<< end >>
