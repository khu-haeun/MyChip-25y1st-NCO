* NGSPICE file created from nco.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL vdd gnd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 D CLK Q vdd gnd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A Y vdd gnd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S Y vdd gnd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A Y vdd gnd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A Y vdd gnd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A Y vdd gnd
.ends

.subckt nco gnd vdd Dout[11] Dout[10] Dout[9] Dout[8] Dout[7] Dout[6] Dout[5] Dout[4]
+ Dout[3] Dout[2] Dout[1] Dout[0] En FCW[19] FCW[18] FCW[17] FCW[16] FCW[15] FCW[14]
+ FCW[13] FCW[12] FCW[11] FCW[10] FCW[9] FCW[8] FCW[7] FCW[6] FCW[5] FCW[4] FCW[3]
+ FCW[2] FCW[1] FCW[0] Vld clk selSign selXY
XFILL_1__13156_ vdd gnd FILL
XFILL_0__12906_ vdd gnd FILL
XFILL_2__9369_ vdd gnd FILL
XFILL_1__10368_ vdd gnd FILL
XFILL_0__13886_ vdd gnd FILL
XFILL_0__7404_ vdd gnd FILL
XFILL_0__8384_ vdd gnd FILL
XFILL_1__12107_ vdd gnd FILL
XFILL_1__13087_ vdd gnd FILL
XFILL_0__12837_ vdd gnd FILL
XFILL_1__10299_ vdd gnd FILL
XFILL_0__7335_ vdd gnd FILL
X_7963_ _7963_/D _7963_/CLK _7963_/Q vdd gnd DFFPOSX1
XFILL_1__12038_ vdd gnd FILL
XFILL_2__11589_ vdd gnd FILL
XFILL_0__12768_ vdd gnd FILL
X_9702_ _9702_/A _9702_/B _9702_/Y vdd gnd NAND2X1
XFILL_0__7266_ vdd gnd FILL
X_7894_ _7894_/A _7894_/Y vdd gnd INVX1
XFILL_0__11719_ vdd gnd FILL
XFILL_0__9005_ vdd gnd FILL
XFILL_0__12699_ vdd gnd FILL
XFILL_0__7197_ vdd gnd FILL
X_9633_ _9633_/A _9633_/B _9633_/Y vdd gnd OR2X2
XFILL_0__14438_ vdd gnd FILL
XFILL_1__13989_ vdd gnd FILL
X_9564_ _9564_/A _9564_/Y vdd gnd INVX1
XFILL_0__14369_ vdd gnd FILL
X_8515_ _8515_/A _8515_/B _8515_/Y vdd gnd AND2X2
X_9495_ _9495_/A _9495_/B _9495_/C _9495_/Y vdd gnd NAND3X1
XFILL_0__9907_ vdd gnd FILL
XFILL_1__8700_ vdd gnd FILL
X_8446_ _8446_/A _8446_/Y vdd gnd INVX1
XFILL_1__9680_ vdd gnd FILL
XFILL_1__8631_ vdd gnd FILL
X_8377_ _8377_/A _8377_/B _8377_/Y vdd gnd NAND2X1
X_7328_ _7328_/A _7328_/Y vdd gnd INVX1
XFILL_1__8562_ vdd gnd FILL
XFILL_1__7513_ vdd gnd FILL
X_7259_ _7259_/A _7259_/Y vdd gnd INVX1
XFILL_1__8493_ vdd gnd FILL
XFILL_1__7444_ vdd gnd FILL
XFILL_2_BUFX2_insert315 vdd gnd FILL
XFILL_1__7375_ vdd gnd FILL
XFILL_2_BUFX2_insert337 vdd gnd FILL
X_11900_ _11900_/A _11900_/Y vdd gnd INVX1
XFILL_1__9114_ vdd gnd FILL
X_12880_ _12880_/A _12880_/Y vdd gnd INVX1
X_11831_ _11831_/A _11831_/B _11831_/S _11831_/Y vdd gnd MUX2X1
XFILL257550x28950 vdd gnd FILL
XFILL_1__9045_ vdd gnd FILL
X_14550_ _14550_/D _14550_/CLK _14550_/Q vdd gnd DFFPOSX1
X_11762_ _11762_/A _11762_/B _11762_/Y vdd gnd NAND2X1
X_13501_ _13501_/D _13501_/CLK _13501_/Q vdd gnd DFFPOSX1
X_10713_ _10713_/D _10713_/CLK _10713_/Q vdd gnd DFFPOSX1
XBUFX2_insert303 BUFX2_insert303/A BUFX2_insert303/Y vdd gnd BUFX2
X_14481_ _14481_/A _14481_/B _14481_/C _14481_/Y vdd gnd OAI21X1
XBUFX2_insert314 BUFX2_insert314/A BUFX2_insert314/Y vdd gnd BUFX2
X_11693_ _11693_/A _11693_/Y vdd gnd INVX2
XBUFX2_insert325 BUFX2_insert325/A BUFX2_insert325/Y vdd gnd BUFX2
XBUFX2_insert336 BUFX2_insert336/A BUFX2_insert336/Y vdd gnd BUFX2
X_13432_ _13432_/D _13432_/CLK _13432_/Q vdd gnd DFFPOSX1
XBUFX2_insert347 BUFX2_insert347/A BUFX2_insert347/Y vdd gnd BUFX2
X_10644_ _10644_/A _10644_/B _10644_/C _10644_/Y vdd gnd OAI21X1
XBUFX2_insert358 BUFX2_insert358/A BUFX2_insert358/Y vdd gnd BUFX2
XFILL_1__9947_ vdd gnd FILL
XBUFX2_insert369 BUFX2_insert369/A BUFX2_insert369/Y vdd gnd BUFX2
X_10575_ _10575_/A _10575_/B _10575_/C _10575_/Y vdd gnd AOI21X1
X_13363_ _13363_/A _13363_/B _13363_/Y vdd gnd AND2X2
XFILL_1__9878_ vdd gnd FILL
X_12314_ _12314_/A _12314_/Y vdd gnd INVX1
XFILL_2__7622_ vdd gnd FILL
XFILL_1__8829_ vdd gnd FILL
X_13294_ _13294_/A _13294_/B _13294_/Y vdd gnd NAND2X1
XFILL_0__10050_ vdd gnd FILL
XFILL_2__10960_ vdd gnd FILL
X_12245_ _12245_/A _12245_/B _12245_/C _12245_/Y vdd gnd OAI21X1
XFILL_2__7553_ vdd gnd FILL
XFILL_1__11340_ vdd gnd FILL
XFILL_2__10891_ vdd gnd FILL
X_12176_ _12176_/A _12176_/B _12176_/Y vdd gnd NAND2X1
XFILL_1__11271_ vdd gnd FILL
XFILL_2__7484_ vdd gnd FILL
X_11127_ _11127_/A _11127_/B _11127_/C _11127_/Y vdd gnd OAI21X1
XFILL_1__13010_ vdd gnd FILL
XFILL_1__10222_ vdd gnd FILL
XFILL_0__13740_ vdd gnd FILL
XFILL_0__10952_ vdd gnd FILL
X_11058_ _11058_/A _11058_/B _11058_/C _11058_/Y vdd gnd NAND3X1
XFILL_1__10153_ vdd gnd FILL
XFILL_0__13671_ vdd gnd FILL
X_10009_ _10009_/A _10009_/Y vdd gnd INVX1
XFILL_0__10883_ vdd gnd FILL
XFILL_2__8105_ vdd gnd FILL
XFILL_0__12622_ vdd gnd FILL
XFILL_0__7120_ vdd gnd FILL
XFILL_1__10084_ vdd gnd FILL
X_14817_ _14817_/A _14817_/B _14817_/Y vdd gnd NAND2X1
XFILL_2__8036_ vdd gnd FILL
XFILL_1__13912_ vdd gnd FILL
X_14748_ _14748_/A _14748_/B _14748_/C _14748_/Y vdd gnd AOI21X1
XFILL_2__10325_ vdd gnd FILL
XFILL_0__11504_ vdd gnd FILL
XFILL_1__13843_ vdd gnd FILL
XFILL_0__12484_ vdd gnd FILL
X_14679_ _14679_/A _14679_/B _14679_/C _14679_/Y vdd gnd AOI21X1
XFILL_2__10256_ vdd gnd FILL
XFILL_0__14223_ vdd gnd FILL
XFILL_0__11435_ vdd gnd FILL
XFILL_1__10986_ vdd gnd FILL
XFILL_1__13774_ vdd gnd FILL
XFILL_2__8938_ vdd gnd FILL
XFILL_2__10187_ vdd gnd FILL
XFILL_1__12725_ vdd gnd FILL
XFILL_0__14154_ vdd gnd FILL
X_8300_ _8300_/A _8300_/Y vdd gnd INVX1
XFILL_0__11366_ vdd gnd FILL
X_9280_ _9280_/A _9280_/B _9280_/C _9280_/Y vdd gnd OAI21X1
XFILL_0__13105_ vdd gnd FILL
XFILL_1__12656_ vdd gnd FILL
XFILL_0__10317_ vdd gnd FILL
XFILL_0__14085_ vdd gnd FILL
X_8231_ _8231_/A _8231_/B _8231_/C _8231_/Y vdd gnd OAI21X1
XFILL_0__11297_ vdd gnd FILL
XFILL_0__7884_ vdd gnd FILL
XFILL_1__11607_ vdd gnd FILL
XFILL_0__13036_ vdd gnd FILL
XFILL_0__10248_ vdd gnd FILL
XFILL_0__9623_ vdd gnd FILL
X_8162_ _8162_/A _8162_/B _8162_/Y vdd gnd NAND2X1
XFILL_1__14326_ vdd gnd FILL
XFILL_1__11538_ vdd gnd FILL
XFILL_2__13877_ vdd gnd FILL
X_7113_ _7113_/A _7113_/B _7113_/Y vdd gnd NAND2X1
XFILL_0__10179_ vdd gnd FILL
XFILL_0__9554_ vdd gnd FILL
X_8093_ _8093_/A _8093_/B _8093_/C _8093_/D _8093_/Y vdd gnd OAI22X1
XFILL_1__14257_ vdd gnd FILL
XFILL_1__11469_ vdd gnd FILL
XFILL_0__8505_ vdd gnd FILL
XFILL_0__9485_ vdd gnd FILL
XFILL_1__13208_ vdd gnd FILL
XFILL_0__13938_ vdd gnd FILL
XFILL_0__8436_ vdd gnd FILL
XFILL_1__13139_ vdd gnd FILL
XFILL_1__7160_ vdd gnd FILL
XFILL_0__13869_ vdd gnd FILL
XFILL_0__8367_ vdd gnd FILL
X_8995_ _8995_/A _8995_/B _8995_/S _8995_/Y vdd gnd MUX2X1
XFILL_0__7318_ vdd gnd FILL
XFILL_1__7091_ vdd gnd FILL
X_7946_ _7946_/D _7946_/CLK _7946_/Q vdd gnd DFFPOSX1
XFILL_0__8298_ vdd gnd FILL
XFILL_0__7249_ vdd gnd FILL
X_7877_ _7877_/A _7877_/B _7877_/C _7877_/Y vdd gnd OAI21X1
X_9616_ _9616_/A _9616_/B _9616_/C _9616_/Y vdd gnd OAI21X1
X_9547_ _9547_/A _9547_/B _9547_/Y vdd gnd AND2X2
XFILL_1__9732_ vdd gnd FILL
X_9478_ _9478_/A _9478_/B _9478_/C _9478_/Y vdd gnd AOI21X1
X_10360_ _10360_/A _10360_/B _10360_/Y vdd gnd NAND2X1
XFILL_1__9663_ vdd gnd FILL
X_8429_ _8429_/A _8429_/B _8429_/Y vdd gnd NOR2X1
X_10291_ _10291_/A _10291_/B _10291_/Y vdd gnd OR2X2
XFILL_1__8614_ vdd gnd FILL
XFILL_1__9594_ vdd gnd FILL
X_12030_ _12030_/A _12030_/B _12030_/C _12030_/Y vdd gnd NAND3X1
XFILL_1__8545_ vdd gnd FILL
XFILL_1__8476_ vdd gnd FILL
X_13981_ _13981_/A _13981_/B _13981_/Y vdd gnd NAND2X1
XFILL_1__7427_ vdd gnd FILL
XFILL_2_BUFX2_insert134 vdd gnd FILL
X_12932_ _12932_/A _12932_/B _12932_/C _12932_/Y vdd gnd OAI21X1
XFILL_1__7358_ vdd gnd FILL
XFILL_2_BUFX2_insert156 vdd gnd FILL
XFILL_2_BUFX2_insert167 vdd gnd FILL
XFILL_2_BUFX2_insert189 vdd gnd FILL
X_12863_ _12863_/A _12863_/B _12863_/C _12863_/Y vdd gnd OAI21X1
XFILL_1__7289_ vdd gnd FILL
X_14602_ _14602_/A _14602_/Y vdd gnd INVX1
X_11814_ _11814_/A _11814_/B _11814_/S _11814_/Y vdd gnd MUX2X1
XFILL_1__9028_ vdd gnd FILL
X_12794_ _12794_/A _12794_/B _12794_/C _12794_/Y vdd gnd AOI21X1
X_14533_ _14533_/D _14533_/CLK _14533_/Q vdd gnd DFFPOSX1
XFILL_2__10110_ vdd gnd FILL
X_11745_ _11745_/A _11745_/B _11745_/C _11745_/Y vdd gnd OAI21X1
XBUFX2_insert111 BUFX2_insert111/A BUFX2_insert111/Y vdd gnd BUFX2
XFILL_1__10840_ vdd gnd FILL
XBUFX2_insert122 BUFX2_insert122/A BUFX2_insert122/Y vdd gnd BUFX2
XBUFX2_insert133 BUFX2_insert133/A BUFX2_insert133/Y vdd gnd BUFX2
X_14464_ _14464_/A _14464_/B _14464_/C _14464_/Y vdd gnd OAI21X1
XFILL_2__10041_ vdd gnd FILL
XBUFX2_insert144 BUFX2_insert144/A BUFX2_insert144/Y vdd gnd BUFX2
X_11676_ _11676_/D _11676_/CLK _11676_/Q vdd gnd DFFPOSX1
XBUFX2_insert155 BUFX2_insert155/A BUFX2_insert155/Y vdd gnd BUFX2
XFILL_0__11220_ vdd gnd FILL
XBUFX2_insert166 BUFX2_insert166/A BUFX2_insert166/Y vdd gnd BUFX2
XFILL_1__10771_ vdd gnd FILL
XBUFX2_insert177 BUFX2_insert177/A BUFX2_insert177/Y vdd gnd BUFX2
X_13415_ _13415_/A _13415_/B _13415_/C _13415_/Y vdd gnd OAI21X1
X_10627_ _10627_/A _10627_/B _10627_/C _10627_/Y vdd gnd OAI21X1
XBUFX2_insert188 BUFX2_insert188/A BUFX2_insert188/Y vdd gnd BUFX2
X_14395_ _14395_/A _14395_/B _14395_/C _14395_/Y vdd gnd NAND3X1
XFILL_1__12510_ vdd gnd FILL
XBUFX2_insert199 BUFX2_insert199/A BUFX2_insert199/Y vdd gnd BUFX2
XFILL_0__11151_ vdd gnd FILL
X_13346_ _13346_/A _13346_/B _13346_/Y vdd gnd NOR2X1
X_10558_ _10558_/A _10558_/B _10558_/Y vdd gnd NAND2X1
XFILL_0__10102_ vdd gnd FILL
XFILL_1__12441_ vdd gnd FILL
XFILL_0__11082_ vdd gnd FILL
X_13277_ _13277_/A _13277_/B _13277_/Y vdd gnd OR2X2
X_10489_ _10489_/A _10489_/B _10489_/Y vdd gnd NOR2X1
XFILL_0__10033_ vdd gnd FILL
XFILL_0__14910_ vdd gnd FILL
XFILL_1__12372_ vdd gnd FILL
XFILL_2__10943_ vdd gnd FILL
X_12228_ _12228_/A _12228_/B _12228_/Y vdd gnd NAND2X1
XFILL_2__7536_ vdd gnd FILL
XFILL_1__14111_ vdd gnd FILL
XFILL_1__11323_ vdd gnd FILL
XFILL_0__14841_ vdd gnd FILL
XFILL_2__10874_ vdd gnd FILL
X_12159_ _12159_/A _12159_/B _12159_/Y vdd gnd OR2X2
XFILL_1__14042_ vdd gnd FILL
XFILL_2__7467_ vdd gnd FILL
XFILL_1__11254_ vdd gnd FILL
XFILL_0__14772_ vdd gnd FILL
XFILL_0__11984_ vdd gnd FILL
XFILL_0__9270_ vdd gnd FILL
XFILL_1__10205_ vdd gnd FILL
XFILL_1__11185_ vdd gnd FILL
XFILL_2__7398_ vdd gnd FILL
XFILL_0__10935_ vdd gnd FILL
XFILL_0__13723_ vdd gnd FILL
XFILL_0__8221_ vdd gnd FILL
XFILL_1__10136_ vdd gnd FILL
XFILL_2__12475_ vdd gnd FILL
XFILL_0__13654_ vdd gnd FILL
XFILL_0__10866_ vdd gnd FILL
X_7800_ _7800_/A _7800_/B _7800_/Y vdd gnd NOR2X1
XFILL_0__8152_ vdd gnd FILL
X_8780_ _8780_/A _8780_/B _8780_/C _8780_/Y vdd gnd OAI21X1
XFILL_1__10067_ vdd gnd FILL
XFILL_0__13585_ vdd gnd FILL
XFILL_0__7103_ vdd gnd FILL
X_7731_ _7731_/A _7731_/Y vdd gnd INVX1
XFILL_0__8083_ vdd gnd FILL
XFILL_0__10797_ vdd gnd FILL
XFILL_2__8019_ vdd gnd FILL
X_7662_ _7662_/A _7662_/B _7662_/Y vdd gnd OR2X2
XFILL_2__10308_ vdd gnd FILL
XFILL_1__13826_ vdd gnd FILL
XFILL_0__12467_ vdd gnd FILL
X_9401_ _9401_/A _9401_/B _9401_/Y vdd gnd NAND2X1
X_7593_ _7593_/A _7593_/B _7593_/C _7593_/Y vdd gnd AOI21X1
XFILL_2__10239_ vdd gnd FILL
XFILL_2__13027_ vdd gnd FILL
XFILL_0__11418_ vdd gnd FILL
XFILL_1__13757_ vdd gnd FILL
XFILL_1__10969_ vdd gnd FILL
XFILL_0__12398_ vdd gnd FILL
X_9332_ _9332_/A _9332_/B _9332_/C _9332_/Y vdd gnd OAI21X1
XFILL_0__8985_ vdd gnd FILL
XFILL_0__14137_ vdd gnd FILL
XFILL_1__12708_ vdd gnd FILL
XFILL_0__11349_ vdd gnd FILL
XFILL_1__13688_ vdd gnd FILL
X_9263_ _9263_/A _9263_/B _9263_/C _9263_/Y vdd gnd OAI21X1
XFILL_0__14068_ vdd gnd FILL
XFILL_1__12639_ vdd gnd FILL
X_8214_ _8214_/A _8214_/B _8214_/C _8214_/Y vdd gnd OAI21X1
X_9194_ _9194_/A _9194_/B _9194_/C _9194_/Y vdd gnd OAI21X1
XFILL_0__7867_ vdd gnd FILL
XFILL_0__13019_ vdd gnd FILL
XFILL_0__9606_ vdd gnd FILL
X_8145_ _8145_/A _8145_/B _8145_/C _8145_/Y vdd gnd NAND3X1
XFILL_0__7798_ vdd gnd FILL
XFILL_1__14309_ vdd gnd FILL
XFILL_0__9537_ vdd gnd FILL
XFILL_1__8330_ vdd gnd FILL
X_8076_ _8076_/A _8076_/B _8076_/Y vdd gnd NAND2X1
XFILL_0__9468_ vdd gnd FILL
XFILL_1__8261_ vdd gnd FILL
XFILL_1__7212_ vdd gnd FILL
XFILL_0__8419_ vdd gnd FILL
XFILL_0__9399_ vdd gnd FILL
XFILL_1__8192_ vdd gnd FILL
XFILL_1__7143_ vdd gnd FILL
X_8978_ _8978_/A _8978_/Y vdd gnd INVX1
XFILL_1_BUFX2_insert108 vdd gnd FILL
XFILL_1_BUFX2_insert119 vdd gnd FILL
XFILL_1__7074_ vdd gnd FILL
X_7929_ _7929_/D _7929_/CLK _7929_/Q vdd gnd DFFPOSX1
X_11530_ _11530_/A _11530_/B _11530_/Y vdd gnd NOR2X1
X_11461_ _11461_/A _11461_/B _11461_/C _11461_/Y vdd gnd OAI21X1
X_13200_ _13200_/A _13200_/B _13200_/C _13200_/Y vdd gnd OAI21X1
X_10412_ _10412_/A _10412_/B _10412_/Y vdd gnd NOR2X1
XFILL_1__9715_ vdd gnd FILL
X_11392_ _11392_/A _11392_/B _11392_/C _11392_/Y vdd gnd AOI21X1
X_14180_ _14180_/D _14180_/CLK _14180_/Q vdd gnd DFFPOSX1
X_13131_ _13131_/A _13131_/B _13131_/C _13131_/Y vdd gnd OAI21X1
X_10343_ _10343_/A _10343_/B _10343_/C _10343_/Y vdd gnd OAI21X1
XFILL_1__9646_ vdd gnd FILL
X_10274_ _10274_/A _10274_/B _10274_/C _10274_/Y vdd gnd AOI21X1
X_13062_ _13062_/A _13062_/B _13062_/Y vdd gnd OR2X2
XFILL_1__9577_ vdd gnd FILL
X_12013_ _12013_/A _12013_/B _12013_/C _12013_/Y vdd gnd OAI21X1
XFILL_1__8528_ vdd gnd FILL
XFILL_1__8459_ vdd gnd FILL
X_13964_ _13964_/A _13964_/B _13964_/C _13964_/D _13964_/Y vdd gnd AOI22X1
X_12915_ _12915_/A _12915_/Y vdd gnd INVX1
X_13895_ _13895_/A _13895_/B _13895_/Y vdd gnd NAND2X1
XFILL257250x93750 vdd gnd FILL
XFILL_2__12260_ vdd gnd FILL
XFILL_0__10651_ vdd gnd FILL
XFILL_1__12990_ vdd gnd FILL
X_12846_ _12846_/A _12846_/B _12846_/C _12846_/Y vdd gnd NAND3X1
XFILL_2__12191_ vdd gnd FILL
XFILL_1__11941_ vdd gnd FILL
XFILL_0__13370_ vdd gnd FILL
XFILL_0__10582_ vdd gnd FILL
X_12777_ _12777_/A _12777_/B _12777_/Y vdd gnd NAND2X1
XFILL_0__12321_ vdd gnd FILL
XFILL_1__14660_ vdd gnd FILL
XFILL_1__11872_ vdd gnd FILL
X_14516_ _14516_/D _14516_/CLK _14516_/Q vdd gnd DFFPOSX1
X_11728_ _11728_/A _11728_/Y vdd gnd INVX1
XFILL_1__13611_ vdd gnd FILL
XFILL_0__12252_ vdd gnd FILL
XFILL_1__10823_ vdd gnd FILL
XFILL_1__14591_ vdd gnd FILL
X_14447_ _14447_/A _14447_/B _14447_/Y vdd gnd NAND2X1
X_11659_ _11659_/D _11659_/CLK _11659_/Q vdd gnd DFFPOSX1
XFILL_2__9755_ vdd gnd FILL
XFILL_0__11203_ vdd gnd FILL
XFILL_1__13542_ vdd gnd FILL
XFILL_0__12183_ vdd gnd FILL
X_14378_ _14378_/A _14378_/B _14378_/C _14378_/Y vdd gnd OAI21X1
XFILL_0__8770_ vdd gnd FILL
XFILL_2__14832_ vdd gnd FILL
XFILL_2__9686_ vdd gnd FILL
XFILL_0__11134_ vdd gnd FILL
XFILL_1__10685_ vdd gnd FILL
XFILL_0__7721_ vdd gnd FILL
X_13329_ _13329_/A _13329_/B _13329_/Y vdd gnd NAND2X1
XFILL_2__14763_ vdd gnd FILL
XFILL_1__12424_ vdd gnd FILL
XFILL_0__11065_ vdd gnd FILL
XFILL_0__7652_ vdd gnd FILL
XFILL_0__10016_ vdd gnd FILL
XFILL_1__12355_ vdd gnd FILL
XFILL256950x216150 vdd gnd FILL
XFILL_0__7583_ vdd gnd FILL
XFILL_1__11306_ vdd gnd FILL
XFILL_0__14824_ vdd gnd FILL
XFILL_1__12286_ vdd gnd FILL
XFILL_0__9322_ vdd gnd FILL
X_9950_ _9950_/A _9950_/B _9950_/S _9950_/Y vdd gnd MUX2X1
XFILL_1__11237_ vdd gnd FILL
XFILL_1__14025_ vdd gnd FILL
XFILL_0__14755_ vdd gnd FILL
XFILL_0__11967_ vdd gnd FILL
XFILL_2__10788_ vdd gnd FILL
XFILL_0__9253_ vdd gnd FILL
X_8901_ _8901_/D _8901_/CLK _8901_/Q vdd gnd DFFPOSX1
X_9881_ _9881_/A _9881_/B _9881_/Y vdd gnd NAND2X1
XFILL_2__12527_ vdd gnd FILL
XFILL_1__11168_ vdd gnd FILL
XFILL_0__10918_ vdd gnd FILL
XFILL_0__13706_ vdd gnd FILL
XFILL_0__8204_ vdd gnd FILL
XFILL_0__14686_ vdd gnd FILL
XFILL_0__11898_ vdd gnd FILL
XFILL_0__9184_ vdd gnd FILL
X_8832_ _8832_/A _8832_/B _8832_/C _8832_/Y vdd gnd OAI21X1
XBUFX2_insert0 BUFX2_insert0/A BUFX2_insert0/Y vdd gnd BUFX2
XFILL_1__10119_ vdd gnd FILL
XFILL_2__12458_ vdd gnd FILL
XFILL_0__13637_ vdd gnd FILL
XFILL257550x244950 vdd gnd FILL
XFILL_0__10849_ vdd gnd FILL
XFILL_1__11099_ vdd gnd FILL
XFILL_0__8135_ vdd gnd FILL
X_8763_ _8763_/A _8763_/Y vdd gnd INVX1
XFILL_2__12389_ vdd gnd FILL
XFILL_0__13568_ vdd gnd FILL
X_7714_ _7714_/A _7714_/B _7714_/Y vdd gnd OR2X2
XFILL_0__8066_ vdd gnd FILL
XFILL_2__14128_ vdd gnd FILL
XFILL_0__12519_ vdd gnd FILL
X_8694_ _8694_/A _8694_/B _8694_/Y vdd gnd NAND2X1
XFILL_1__14858_ vdd gnd FILL
X_7645_ _7645_/A _7645_/B _7645_/Y vdd gnd NAND2X1
XFILL_2__14059_ vdd gnd FILL
XFILL_1__13809_ vdd gnd FILL
XFILL_1__14789_ vdd gnd FILL
XFILL257550x7350 vdd gnd FILL
XFILL_1__7830_ vdd gnd FILL
X_7576_ _7576_/A _7576_/B _7576_/C _7576_/Y vdd gnd OAI21X1
X_9315_ _9315_/A _9315_/Y vdd gnd INVX1
XFILL_0__8968_ vdd gnd FILL
XFILL_1__7761_ vdd gnd FILL
XFILL_1__9500_ vdd gnd FILL
X_9246_ _9246_/A _9246_/B _9246_/C _9246_/Y vdd gnd NAND3X1
XFILL_1__7692_ vdd gnd FILL
XFILL_1__9431_ vdd gnd FILL
X_9177_ _9177_/A _9177_/B _9177_/C _9177_/Y vdd gnd NAND3X1
XFILL256950x126150 vdd gnd FILL
X_8128_ _8128_/A _8128_/Y vdd gnd INVX1
XFILL_1__9362_ vdd gnd FILL
XFILL_1__8313_ vdd gnd FILL
X_8059_ _8059_/A _8059_/B _8059_/Y vdd gnd NAND2X1
XFILL_1__9293_ vdd gnd FILL
XFILL_1__8244_ vdd gnd FILL
X_10961_ _10961_/A _10961_/B _10961_/C _10961_/Y vdd gnd OAI21X1
XFILL_1__8175_ vdd gnd FILL
XFILL257550x154950 vdd gnd FILL
X_12700_ _12700_/A _12700_/Y vdd gnd INVX2
XFILL_1__7126_ vdd gnd FILL
X_13680_ _13680_/A _13680_/Y vdd gnd INVX2
X_10892_ _10892_/A _10892_/B _10892_/C _10892_/Y vdd gnd AOI21X1
X_12631_ _12631_/A _12631_/B _12631_/C _12631_/D _12631_/Y vdd gnd AOI22X1
XFILL257250x25350 vdd gnd FILL
XFILL_1_CLKBUF1_insert60 vdd gnd FILL
X_12562_ _12562_/D _12562_/CLK _12562_/Q vdd gnd DFFPOSX1
XFILL_1_CLKBUF1_insert71 vdd gnd FILL
XFILL_1_CLKBUF1_insert82 vdd gnd FILL
XFILL_2__7870_ vdd gnd FILL
XFILL_1_CLKBUF1_insert93 vdd gnd FILL
X_14301_ _14301_/A _14301_/Y vdd gnd INVX1
X_11513_ _11513_/A _11513_/B _11513_/Y vdd gnd NAND2X1
X_12493_ _12493_/A _12493_/B _12493_/C _12493_/Y vdd gnd OAI21X1
X_14232_ _14232_/A _14232_/B _14232_/Y vdd gnd NAND2X1
X_11444_ _11444_/A _11444_/B _11444_/C _11444_/Y vdd gnd OAI21X1
X_14163_ _14163_/D _14163_/CLK _14163_/Q vdd gnd DFFPOSX1
X_11375_ _11375_/A _11375_/B _11375_/Y vdd gnd NOR2X1
XFILL_1__10470_ vdd gnd FILL
X_13114_ _13114_/A _13114_/B _13114_/C _13114_/Y vdd gnd NAND3X1
X_10326_ _10326_/A _10326_/B _10326_/Y vdd gnd NOR2X1
XFILL_1__9629_ vdd gnd FILL
XFILL_2__8422_ vdd gnd FILL
X_14094_ _14094_/A _14094_/B _14094_/C _14094_/Y vdd gnd AOI21X1
XFILL_2__11760_ vdd gnd FILL
X_13045_ _13045_/A _13045_/B _13045_/C _13045_/Y vdd gnd OAI21X1
X_10257_ _10257_/A _10257_/B _10257_/Y vdd gnd NAND2X1
XFILL_2__8353_ vdd gnd FILL
XFILL_1__12140_ vdd gnd FILL
XFILL_0__12870_ vdd gnd FILL
X_10188_ _10188_/A _10188_/B _10188_/Y vdd gnd OR2X2
XFILL_2__10642_ vdd gnd FILL
XFILL_0__11821_ vdd gnd FILL
XFILL_2__8284_ vdd gnd FILL
XFILL_1__12071_ vdd gnd FILL
XFILL_1__11022_ vdd gnd FILL
XFILL_2__10573_ vdd gnd FILL
XFILL_0__11752_ vdd gnd FILL
X_13947_ _13947_/A _13947_/B _13947_/C _13947_/Y vdd gnd OAI21X1
XFILL_0__14471_ vdd gnd FILL
X_13878_ _13878_/A _13878_/B _13878_/Y vdd gnd NAND2X1
XFILL_0__13422_ vdd gnd FILL
XFILL_0__10634_ vdd gnd FILL
XFILL_1__12973_ vdd gnd FILL
X_12829_ _12829_/A _12829_/B _12829_/C _12829_/Y vdd gnd AOI21X1
XFILL_1__14712_ vdd gnd FILL
XFILL_1__11924_ vdd gnd FILL
XFILL_2__12174_ vdd gnd FILL
XFILL_0__13353_ vdd gnd FILL
XFILL_0__10565_ vdd gnd FILL
XFILL_0__9940_ vdd gnd FILL
XFILL_0__12304_ vdd gnd FILL
XFILL_2__11125_ vdd gnd FILL
XFILL_1__14643_ vdd gnd FILL
XFILL_1__11855_ vdd gnd FILL
XFILL_0__13284_ vdd gnd FILL
X_7430_ _7430_/A _7430_/B _7430_/C _7430_/Y vdd gnd AOI21X1
XFILL_0__10496_ vdd gnd FILL
XFILL_0__9871_ vdd gnd FILL
XFILL_0__12235_ vdd gnd FILL
XFILL_1__10806_ vdd gnd FILL
XFILL_1__14574_ vdd gnd FILL
XFILL_0__8822_ vdd gnd FILL
XFILL_1__11786_ vdd gnd FILL
X_7361_ _7361_/A _7361_/B _7361_/C _7361_/Y vdd gnd OAI21X1
XFILL_1__13525_ vdd gnd FILL
XFILL_0__12166_ vdd gnd FILL
X_9100_ _9100_/A _9100_/Y vdd gnd INVX1
XFILL_0__8753_ vdd gnd FILL
X_7292_ _7292_/A _7292_/B _7292_/C _7292_/Y vdd gnd AOI21X1
XFILL_2__14815_ vdd gnd FILL
XFILL_0__11117_ vdd gnd FILL
XFILL_1__10668_ vdd gnd FILL
X_9031_ _9031_/A _9031_/B _9031_/Y vdd gnd NAND2X1
XFILL_0__7704_ vdd gnd FILL
XFILL_0__12097_ vdd gnd FILL
XFILL_0__8684_ vdd gnd FILL
XFILL_2__14746_ vdd gnd FILL
XFILL_1__12407_ vdd gnd FILL
XFILL_0__11048_ vdd gnd FILL
XFILL_2__11958_ vdd gnd FILL
XFILL_1__10599_ vdd gnd FILL
XFILL_1__13387_ vdd gnd FILL
XFILL_0__7635_ vdd gnd FILL
XFILL_2__14677_ vdd gnd FILL
XFILL_1__12338_ vdd gnd FILL
XFILL_0__7566_ vdd gnd FILL
XFILL_0__14807_ vdd gnd FILL
XFILL_1__12269_ vdd gnd FILL
XFILL_0__9305_ vdd gnd FILL
X_9933_ _9933_/A _9933_/B _9933_/S _9933_/Y vdd gnd MUX2X1
XFILL_0__12999_ vdd gnd FILL
XFILL_1__14008_ vdd gnd FILL
XFILL_0__7497_ vdd gnd FILL
XFILL_0__14738_ vdd gnd FILL
XFILL_0__9236_ vdd gnd FILL
X_9864_ _9864_/A _9864_/B _9864_/C _9864_/Y vdd gnd OAI21X1
XFILL_0__14669_ vdd gnd FILL
XFILL_0__9167_ vdd gnd FILL
X_8815_ _8815_/A _8815_/B _8815_/C _8815_/Y vdd gnd OAI21X1
X_9795_ _9795_/D _9795_/CLK _9795_/Q vdd gnd DFFPOSX1
XFILL_0__8118_ vdd gnd FILL
XFILL_0__9098_ vdd gnd FILL
XFILL_1__9980_ vdd gnd FILL
X_8746_ _8746_/A _8746_/Y vdd gnd INVX1
XFILL_1__8931_ vdd gnd FILL
XFILL_0__8049_ vdd gnd FILL
X_8677_ _8677_/A _8677_/B _8677_/Y vdd gnd NAND2X1
X_7628_ _7628_/A _7628_/B _7628_/C _7628_/Y vdd gnd OAI21X1
XFILL_1_CLKBUF1_insert104 vdd gnd FILL
XFILL_1__7813_ vdd gnd FILL
X_7559_ _7559_/A _7559_/B _7559_/C _7559_/Y vdd gnd NAND3X1
XFILL_1__8793_ vdd gnd FILL
XFILL_1__7744_ vdd gnd FILL
X_11160_ _11160_/A _11160_/B _11160_/Y vdd gnd NAND2X1
X_9229_ _9229_/A _9229_/B _9229_/C _9229_/Y vdd gnd OAI21X1
XFILL_1__7675_ vdd gnd FILL
X_10111_ _10111_/A _10111_/B _10111_/C _10111_/Y vdd gnd NAND3X1
X_11091_ _11091_/A _11091_/B _11091_/C _11091_/Y vdd gnd OAI21X1
XFILL_1__9414_ vdd gnd FILL
X_10042_ _10042_/A _10042_/B _10042_/C _10042_/Y vdd gnd OAI21X1
XFILL_1__9345_ vdd gnd FILL
X_14850_ _14850_/A _14850_/B _14850_/C _14850_/Y vdd gnd OAI21X1
XFILL_1__9276_ vdd gnd FILL
X_13801_ _13801_/A _13801_/B _13801_/C _13801_/Y vdd gnd OAI21X1
X_14781_ _14781_/A _14781_/B _14781_/C _14781_/Y vdd gnd AOI21X1
XFILL_1__8227_ vdd gnd FILL
X_11993_ _11993_/A _11993_/B _11993_/Y vdd gnd AND2X2
X_13732_ _13732_/A _13732_/B _13732_/C _13732_/Y vdd gnd AOI21X1
X_10944_ _10944_/A _10944_/Y vdd gnd INVX1
XFILL_1__8158_ vdd gnd FILL
X_13663_ _13663_/A _13663_/B _13663_/C _13663_/Y vdd gnd OAI21X1
XFILL_1__7109_ vdd gnd FILL
X_10875_ _10875_/A _10875_/Y vdd gnd INVX1
XFILL_2__8971_ vdd gnd FILL
XFILL_1__8089_ vdd gnd FILL
X_12614_ _12614_/D _12614_/CLK _12614_/Q vdd gnd DFFPOSX1
X_13594_ _13594_/A _13594_/B _13594_/Y vdd gnd NAND2X1
XFILL_0__10350_ vdd gnd FILL
X_12545_ _12545_/D _12545_/CLK _12545_/Q vdd gnd DFFPOSX1
XFILL_2__7853_ vdd gnd FILL
XFILL_0__10281_ vdd gnd FILL
X_12476_ _12476_/A _12476_/B _12476_/C _12476_/Y vdd gnd OAI21X1
XFILL_0__12020_ vdd gnd FILL
XFILL_2__7784_ vdd gnd FILL
XFILL_1__11571_ vdd gnd FILL
X_14215_ _14215_/D _14215_/CLK _14215_/Q vdd gnd DFFPOSX1
X_11427_ _11427_/A _11427_/Y vdd gnd INVX1
XFILL_1__10522_ vdd gnd FILL
XFILL_1__13310_ vdd gnd FILL
XFILL_1__14290_ vdd gnd FILL
X_14146_ _14146_/A _14146_/B _14146_/C _14146_/Y vdd gnd OAI21X1
X_11358_ _11358_/A _11358_/B _11358_/Y vdd gnd OR2X2
XFILL_2__11812_ vdd gnd FILL
XFILL_1__10453_ vdd gnd FILL
XCLKBUF1_insert103 CLKBUF1_insert103/A CLKBUF1_insert103/Y vdd gnd CLKBUF1
XFILL_1__13241_ vdd gnd FILL
XFILL_0__13971_ vdd gnd FILL
X_10309_ _10309_/A _10309_/B _10309_/C _10309_/Y vdd gnd NAND3X1
XFILL_2__8405_ vdd gnd FILL
X_14077_ _14077_/A _14077_/B _14077_/C _14077_/Y vdd gnd OAI21X1
X_11289_ _11289_/A _11289_/B _11289_/C _11289_/Y vdd gnd AOI21X1
XFILL_1__13172_ vdd gnd FILL
XFILL_2__11743_ vdd gnd FILL
XFILL_0__12922_ vdd gnd FILL
XFILL_1__10384_ vdd gnd FILL
XFILL_0__7420_ vdd gnd FILL
X_13028_ _13028_/A _13028_/B _13028_/C _13028_/Y vdd gnd OAI21X1
XFILL_2__8336_ vdd gnd FILL
XFILL_1__12123_ vdd gnd FILL
XFILL_0__12853_ vdd gnd FILL
XFILL_0__7351_ vdd gnd FILL
XFILL_2__13413_ vdd gnd FILL
XFILL_2__10625_ vdd gnd FILL
XFILL_2__8267_ vdd gnd FILL
XFILL_1__12054_ vdd gnd FILL
XFILL_0__11804_ vdd gnd FILL
XFILL_0__12784_ vdd gnd FILL
XFILL_1__11005_ vdd gnd FILL
XFILL_0__7282_ vdd gnd FILL
XFILL_2__10556_ vdd gnd FILL
XFILL_0__11735_ vdd gnd FILL
XFILL_2__8198_ vdd gnd FILL
XFILL_0__9021_ vdd gnd FILL
XFILL_2__10487_ vdd gnd FILL
XFILL_0__14454_ vdd gnd FILL
X_8600_ _8600_/A _8600_/Y vdd gnd INVX1
X_9580_ _9580_/A _9580_/B _9580_/Y vdd gnd NOR2X1
XFILL_0__10617_ vdd gnd FILL
XFILL_0__13405_ vdd gnd FILL
XFILL_1__12956_ vdd gnd FILL
XFILL_0__14385_ vdd gnd FILL
XFILL_0__11597_ vdd gnd FILL
XFILL_1_BUFX2_insert280 vdd gnd FILL
XCLKBUF1_insert40 CLKBUF1_insert40/A CLKBUF1_insert40/Y vdd gnd CLKBUF1
X_8531_ _8531_/A _8531_/B _8531_/C _8531_/Y vdd gnd OAI21X1
XFILL_1_BUFX2_insert291 vdd gnd FILL
XCLKBUF1_insert51 CLKBUF1_insert51/A CLKBUF1_insert51/Y vdd gnd CLKBUF1
XFILL_1__11907_ vdd gnd FILL
XFILL_0__10548_ vdd gnd FILL
XCLKBUF1_insert62 CLKBUF1_insert62/A CLKBUF1_insert62/Y vdd gnd CLKBUF1
XFILL_0__13336_ vdd gnd FILL
XCLKBUF1_insert73 CLKBUF1_insert73/A CLKBUF1_insert73/Y vdd gnd CLKBUF1
XFILL_0__9923_ vdd gnd FILL
XFILL_1__12887_ vdd gnd FILL
XCLKBUF1_insert84 CLKBUF1_insert84/A CLKBUF1_insert84/Y vdd gnd CLKBUF1
X_8462_ _8462_/A _8462_/B _8462_/C _8462_/Y vdd gnd OAI21X1
XCLKBUF1_insert95 CLKBUF1_insert95/A CLKBUF1_insert95/Y vdd gnd CLKBUF1
XFILL_2__11108_ vdd gnd FILL
XFILL_1__14626_ vdd gnd FILL
XFILL_1__11838_ vdd gnd FILL
XFILL_0__13267_ vdd gnd FILL
XFILL_0__10479_ vdd gnd FILL
X_7413_ _7413_/A _7413_/B _7413_/C _7413_/Y vdd gnd NAND3X1
XFILL_0__9854_ vdd gnd FILL
X_8393_ _8393_/A _8393_/B _8393_/C _8393_/Y vdd gnd OAI21X1
XFILL_2__11039_ vdd gnd FILL
XFILL_0__12218_ vdd gnd FILL
XFILL_1__14557_ vdd gnd FILL
XFILL_0__13198_ vdd gnd FILL
XFILL_1__11769_ vdd gnd FILL
XFILL_0__8805_ vdd gnd FILL
X_7344_ _7344_/A _7344_/B _7344_/Y vdd gnd NOR2X1
XFILL_1__13508_ vdd gnd FILL
XFILL_0__12149_ vdd gnd FILL
XFILL_1__14488_ vdd gnd FILL
XFILL_0__8736_ vdd gnd FILL
X_7275_ _7275_/A _7275_/B _7275_/Y vdd gnd NAND2X1
X_9014_ _9014_/A _9014_/B _9014_/C _9014_/Y vdd gnd NAND3X1
XFILL_1__7460_ vdd gnd FILL
XFILL_0__8667_ vdd gnd FILL
XFILL_2__14729_ vdd gnd FILL
XFILL_0__7618_ vdd gnd FILL
XFILL_1__7391_ vdd gnd FILL
XFILL_0__8598_ vdd gnd FILL
XFILL_1__9130_ vdd gnd FILL
XFILL_0__7549_ vdd gnd FILL
XFILL_1__9061_ vdd gnd FILL
X_9916_ _9916_/A _9916_/Y vdd gnd INVX1
XFILL_0__9219_ vdd gnd FILL
XFILL_1__8012_ vdd gnd FILL
X_9847_ _9847_/A _9847_/Y vdd gnd INVX2
X_9778_ _9778_/D _9778_/CLK _9778_/Q vdd gnd DFFPOSX1
X_10660_ _10660_/A _10660_/B _10660_/Y vdd gnd NAND2X1
XFILL_1__9963_ vdd gnd FILL
X_8729_ _8729_/A _8729_/B _8729_/C _8729_/Y vdd gnd OAI21X1
X_10591_ _10591_/A _10591_/B _10591_/C _10591_/Y vdd gnd NAND3X1
XFILL_1__9894_ vdd gnd FILL
X_12330_ _12330_/A _12330_/B _12330_/C _12330_/Y vdd gnd OAI21X1
X_12261_ _12261_/A _12261_/B _12261_/Y vdd gnd NOR2X1
XFILL_1__8776_ vdd gnd FILL
X_14000_ _14000_/A _14000_/B _14000_/Y vdd gnd NOR2X1
X_11212_ _11212_/A _11212_/B _11212_/Y vdd gnd NAND2X1
XFILL_1__7727_ vdd gnd FILL
X_12192_ _12192_/A _12192_/Y vdd gnd INVX1
X_11143_ _11143_/A _11143_/B _11143_/S _11143_/Y vdd gnd MUX2X1
XFILL_1__7658_ vdd gnd FILL
X_11074_ _11074_/A _11074_/Y vdd gnd INVX1
XFILL_1__7589_ vdd gnd FILL
X_14902_ _14902_/D _14902_/CLK _14902_/Q vdd gnd DFFPOSX1
X_10025_ _10025_/A _10025_/B _10025_/Y vdd gnd NAND2X1
XFILL_1__9328_ vdd gnd FILL
X_14833_ _14833_/A _14833_/B _14833_/Y vdd gnd NAND2X1
XFILL_1__9259_ vdd gnd FILL
X_14764_ _14764_/A _14764_/B _14764_/Y vdd gnd OR2X2
X_11976_ _11976_/A _11976_/B _11976_/Y vdd gnd OR2X2
XFILL_2__10341_ vdd gnd FILL
XFILL_0__11520_ vdd gnd FILL
X_13715_ _13715_/A _13715_/B _13715_/C _13715_/Y vdd gnd NAND3X1
X_10927_ _10927_/A _10927_/Y vdd gnd INVX1
X_14695_ _14695_/A _14695_/B _14695_/Y vdd gnd OR2X2
XFILL_2__10272_ vdd gnd FILL
XFILL_1__12810_ vdd gnd FILL
XFILL_2__13060_ vdd gnd FILL
XFILL_0__11451_ vdd gnd FILL
XFILL_1__13790_ vdd gnd FILL
X_13646_ _13646_/A _13646_/Y vdd gnd INVX2
X_10858_ _10858_/A _10858_/B _10858_/S _10858_/Y vdd gnd MUX2X1
XFILL_0__10402_ vdd gnd FILL
XFILL_0_BUFX2_insert210 vdd gnd FILL
XFILL_1__12741_ vdd gnd FILL
XFILL_0_BUFX2_insert221 vdd gnd FILL
XFILL_0__11382_ vdd gnd FILL
XFILL_0_BUFX2_insert232 vdd gnd FILL
X_13577_ _13577_/A _13577_/Y vdd gnd INVX1
XFILL_0__13121_ vdd gnd FILL
XFILL_0_BUFX2_insert243 vdd gnd FILL
X_10789_ _10789_/A _10789_/B _10789_/C _10789_/Y vdd gnd OAI21X1
XFILL_0__10333_ vdd gnd FILL
XFILL_0_BUFX2_insert254 vdd gnd FILL
XFILL_0_BUFX2_insert265 vdd gnd FILL
XFILL_1__12672_ vdd gnd FILL
XFILL_0_BUFX2_insert276 vdd gnd FILL
X_12528_ _12528_/A _12528_/B _12528_/C _12528_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert287 vdd gnd FILL
XFILL_1__14411_ vdd gnd FILL
XFILL_0_BUFX2_insert298 vdd gnd FILL
XFILL_0__13052_ vdd gnd FILL
XFILL_0__10264_ vdd gnd FILL
X_12459_ _12459_/A _12459_/Y vdd gnd INVX1
XFILL_0__12003_ vdd gnd FILL
XFILL_1__14342_ vdd gnd FILL
XFILL_1__11554_ vdd gnd FILL
XFILL_0__10195_ vdd gnd FILL
XFILL_0__9570_ vdd gnd FILL
XFILL_1__10505_ vdd gnd FILL
XFILL_2_BUFX2_insert25 vdd gnd FILL
XFILL_2__7698_ vdd gnd FILL
XFILL_1__14273_ vdd gnd FILL
XFILL_0__8521_ vdd gnd FILL
XFILL_1__11485_ vdd gnd FILL
X_14129_ _14129_/A _14129_/B _14129_/Y vdd gnd NAND2X1
XFILL_1__13224_ vdd gnd FILL
XFILL_1__10436_ vdd gnd FILL
XFILL_0__13954_ vdd gnd FILL
XFILL_0__8452_ vdd gnd FILL
XFILL_2__11726_ vdd gnd FILL
XFILL_1__13155_ vdd gnd FILL
XFILL_0__12905_ vdd gnd FILL
XFILL_1__10367_ vdd gnd FILL
XFILL_0__7403_ vdd gnd FILL
XFILL_0__13885_ vdd gnd FILL
XFILL_2__8319_ vdd gnd FILL
XFILL_0__8383_ vdd gnd FILL
XFILL_1__12106_ vdd gnd FILL
XFILL_1__13086_ vdd gnd FILL
XFILL_1__10298_ vdd gnd FILL
XFILL_0__12836_ vdd gnd FILL
XFILL_0__7334_ vdd gnd FILL
X_7962_ _7962_/D _7962_/CLK _7962_/Q vdd gnd DFFPOSX1
XFILL_2__10608_ vdd gnd FILL
XFILL_1__12037_ vdd gnd FILL
X_9701_ _9701_/A _9701_/B _9701_/C _9701_/Y vdd gnd OAI21X1
XFILL_0__12767_ vdd gnd FILL
XFILL_0__7265_ vdd gnd FILL
XFILL_2__13327_ vdd gnd FILL
X_7893_ _7893_/A _7893_/B _7893_/C _7893_/Y vdd gnd OAI21X1
XFILL_2__10539_ vdd gnd FILL
XFILL_0__9004_ vdd gnd FILL
XFILL_0__11718_ vdd gnd FILL
X_9632_ _9632_/A _9632_/B _9632_/Y vdd gnd NAND2X1
XFILL_0__12698_ vdd gnd FILL
XFILL_0__7196_ vdd gnd FILL
XFILL_2__13258_ vdd gnd FILL
XFILL_0__14437_ vdd gnd FILL
XFILL_1__13988_ vdd gnd FILL
X_9563_ _9563_/A _9563_/B _9563_/Y vdd gnd NAND2X1
XFILL_2__13189_ vdd gnd FILL
XFILL_1__12939_ vdd gnd FILL
XFILL_0__14368_ vdd gnd FILL
X_8514_ _8514_/A _8514_/B _8514_/Y vdd gnd AND2X2
X_9494_ _9494_/A _9494_/B _9494_/Y vdd gnd OR2X2
XFILL_0__13319_ vdd gnd FILL
XFILL_0__9906_ vdd gnd FILL
XFILL_0__14299_ vdd gnd FILL
X_8445_ _8445_/A _8445_/B _8445_/C _8445_/Y vdd gnd AOI21X1
XFILL_1__14609_ vdd gnd FILL
XFILL_1__8630_ vdd gnd FILL
X_8376_ _8376_/A _8376_/B _8376_/Y vdd gnd NAND2X1
X_7327_ _7327_/A _7327_/B _7327_/C _7327_/Y vdd gnd AOI21X1
XFILL_1__8561_ vdd gnd FILL
XFILL_1__7512_ vdd gnd FILL
XFILL_0__8719_ vdd gnd FILL
X_7258_ _7258_/A _7258_/Y vdd gnd INVX1
XFILL_0__9699_ vdd gnd FILL
XFILL_1__8492_ vdd gnd FILL
XFILL_1__7443_ vdd gnd FILL
X_7189_ _7189_/A _7189_/B _7189_/S _7189_/Y vdd gnd MUX2X1
XFILL_1__7374_ vdd gnd FILL
XFILL_1_BUFX2_insert0 vdd gnd FILL
XFILL_2_BUFX2_insert327 vdd gnd FILL
XFILL_1__9113_ vdd gnd FILL
XFILL_2_BUFX2_insert349 vdd gnd FILL
X_11830_ _11830_/A _11830_/B _11830_/S _11830_/Y vdd gnd MUX2X1
XFILL_1__9044_ vdd gnd FILL
X_11761_ _11761_/A _11761_/Y vdd gnd INVX1
X_13500_ _13500_/D _13500_/CLK _13500_/Q vdd gnd DFFPOSX1
X_10712_ _10712_/D _10712_/CLK _10712_/Q vdd gnd DFFPOSX1
X_14480_ _14480_/A _14480_/B _14480_/Y vdd gnd NAND2X1
XBUFX2_insert304 BUFX2_insert304/A BUFX2_insert304/Y vdd gnd BUFX2
X_11692_ _11692_/A _11692_/Y vdd gnd INVX1
XBUFX2_insert315 BUFX2_insert315/A BUFX2_insert315/Y vdd gnd BUFX2
XBUFX2_insert326 BUFX2_insert326/A BUFX2_insert326/Y vdd gnd BUFX2
X_13431_ _13431_/D _13431_/CLK _13431_/Q vdd gnd DFFPOSX1
XBUFX2_insert337 BUFX2_insert337/A BUFX2_insert337/Y vdd gnd BUFX2
X_10643_ _10643_/A _10643_/Y vdd gnd INVX1
XBUFX2_insert348 BUFX2_insert348/A BUFX2_insert348/Y vdd gnd BUFX2
XBUFX2_insert359 BUFX2_insert359/A BUFX2_insert359/Y vdd gnd BUFX2
XFILL_1__9946_ vdd gnd FILL
X_13362_ _13362_/A _13362_/B _13362_/C _13362_/Y vdd gnd OAI21X1
X_10574_ _10574_/A _10574_/B _10574_/Y vdd gnd NOR2X1
XFILL_2__8670_ vdd gnd FILL
XFILL_1__9877_ vdd gnd FILL
X_12313_ _12313_/A _12313_/B _12313_/Y vdd gnd NAND2X1
X_13293_ _13293_/A _13293_/B _13293_/Y vdd gnd NOR2X1
XFILL_1__8828_ vdd gnd FILL
X_12244_ _12244_/A _12244_/Y vdd gnd INVX1
XFILL_1__8759_ vdd gnd FILL
X_12175_ _12175_/A _12175_/B _12175_/C _12175_/Y vdd gnd AOI21X1
XFILL_1__11270_ vdd gnd FILL
X_11126_ _11126_/A _11126_/B _11126_/C _11126_/Y vdd gnd AOI21X1
XFILL_2__9222_ vdd gnd FILL
XFILL_1__10221_ vdd gnd FILL
XFILL_0__10951_ vdd gnd FILL
X_11057_ _11057_/A _11057_/B _11057_/C _11057_/Y vdd gnd OAI21X1
XFILL_2__11511_ vdd gnd FILL
XFILL_1__10152_ vdd gnd FILL
XFILL_2__12491_ vdd gnd FILL
X_10008_ _10008_/A _10008_/B _10008_/C _10008_/Y vdd gnd NAND3X1
XFILL_0__13670_ vdd gnd FILL
XFILL_0__10882_ vdd gnd FILL
XFILL_2__14230_ vdd gnd FILL
XFILL_0__12621_ vdd gnd FILL
XFILL_1__10083_ vdd gnd FILL
X_14816_ _14816_/A _14816_/B _14816_/C _14816_/Y vdd gnd AOI21X1
XFILL_1__13911_ vdd gnd FILL
XFILL_2__13112_ vdd gnd FILL
X_14747_ _14747_/A _14747_/B _14747_/C _14747_/Y vdd gnd OAI21X1
X_11959_ _11959_/A _11959_/B _11959_/C _11959_/Y vdd gnd NAND3X1
XFILL_0__11503_ vdd gnd FILL
XFILL_1__13842_ vdd gnd FILL
XFILL_2__14092_ vdd gnd FILL
XFILL_0__12483_ vdd gnd FILL
X_14678_ _14678_/A _14678_/B _14678_/C _14678_/Y vdd gnd OAI21X1
XFILL_2__13043_ vdd gnd FILL
XFILL_0__14222_ vdd gnd FILL
XFILL_0__11434_ vdd gnd FILL
XFILL_2__9986_ vdd gnd FILL
XFILL_1__13773_ vdd gnd FILL
X_13629_ _13629_/A _13629_/B _13629_/C _13629_/Y vdd gnd AOI21X1
XFILL_1__10985_ vdd gnd FILL
XFILL_1__12724_ vdd gnd FILL
XFILL_0__11365_ vdd gnd FILL
XFILL_0__14153_ vdd gnd FILL
XFILL_0__13104_ vdd gnd FILL
XFILL_0__10316_ vdd gnd FILL
XFILL_1__12655_ vdd gnd FILL
XFILL_0__14084_ vdd gnd FILL
XFILL_0__11296_ vdd gnd FILL
X_8230_ _8230_/A _8230_/Y vdd gnd INVX1
XFILL_0__7883_ vdd gnd FILL
XFILL_1__11606_ vdd gnd FILL
XFILL_0__13035_ vdd gnd FILL
XFILL_0__10247_ vdd gnd FILL
XFILL_0__9622_ vdd gnd FILL
X_8161_ _8161_/A _8161_/Y vdd gnd INVX1
XFILL_1__14325_ vdd gnd FILL
XFILL_1__11537_ vdd gnd FILL
XFILL_0__10178_ vdd gnd FILL
X_7112_ _7112_/A _7112_/B _7112_/C _7112_/D _7112_/Y vdd gnd AOI22X1
XFILL_0__9553_ vdd gnd FILL
X_8092_ _8092_/A _8092_/B _8092_/C _8092_/Y vdd gnd NAND3X1
XFILL_1__14256_ vdd gnd FILL
XFILL_0__8504_ vdd gnd FILL
XFILL_1__11468_ vdd gnd FILL
XFILL_0__9484_ vdd gnd FILL
XFILL_1__13207_ vdd gnd FILL
XFILL_1__10419_ vdd gnd FILL
XFILL_0__13937_ vdd gnd FILL
XFILL_0__8435_ vdd gnd FILL
XFILL_1__11399_ vdd gnd FILL
XFILL_1__13138_ vdd gnd FILL
XFILL_0__13868_ vdd gnd FILL
XFILL_0__8366_ vdd gnd FILL
XFILL_2__14428_ vdd gnd FILL
X_8994_ _8994_/A _8994_/B _8994_/C _8994_/Y vdd gnd OAI21X1
XFILL_0__12819_ vdd gnd FILL
XFILL_1__13069_ vdd gnd FILL
XFILL_0__7317_ vdd gnd FILL
XFILL_0__13799_ vdd gnd FILL
XFILL_1__7090_ vdd gnd FILL
X_7945_ _7945_/D _7945_/CLK _7945_/Q vdd gnd DFFPOSX1
XFILL_0__8297_ vdd gnd FILL
XFILL_2__14359_ vdd gnd FILL
XFILL_0__7248_ vdd gnd FILL
X_7876_ _7876_/A _7876_/B _7876_/Y vdd gnd NAND2X1
X_9615_ _9615_/A _9615_/B _9615_/C _9615_/Y vdd gnd OAI21X1
XFILL_0__7179_ vdd gnd FILL
X_9546_ _9546_/A _9546_/B _9546_/C _9546_/Y vdd gnd OAI21X1
XFILL_1__9731_ vdd gnd FILL
X_9477_ _9477_/A _9477_/B _9477_/Y vdd gnd NAND2X1
XFILL_1__9662_ vdd gnd FILL
X_8428_ _8428_/A _8428_/B _8428_/Y vdd gnd AND2X2
XFILL_1__8613_ vdd gnd FILL
X_10290_ _10290_/A _10290_/B _10290_/C _10290_/Y vdd gnd OAI21X1
XFILL_1__9593_ vdd gnd FILL
X_8359_ _8359_/A _8359_/Y vdd gnd INVX1
XFILL_1__8544_ vdd gnd FILL
XFILL_1__8475_ vdd gnd FILL
X_13980_ _13980_/A _13980_/B _13980_/C _13980_/Y vdd gnd NAND3X1
XFILL_1__7426_ vdd gnd FILL
XFILL257250x165750 vdd gnd FILL
XFILL_2_BUFX2_insert113 vdd gnd FILL
X_12931_ _12931_/A _12931_/Y vdd gnd INVX1
XFILL_1__7357_ vdd gnd FILL
XFILL_2_BUFX2_insert146 vdd gnd FILL
X_12862_ _12862_/A _12862_/B _12862_/C _12862_/Y vdd gnd AOI21X1
XFILL_2_BUFX2_insert179 vdd gnd FILL
XFILL_1__7288_ vdd gnd FILL
X_14601_ _14601_/A _14601_/B _14601_/Y vdd gnd NOR2X1
X_11813_ _11813_/A _11813_/B _11813_/S _11813_/Y vdd gnd MUX2X1
XFILL_1__9027_ vdd gnd FILL
X_12793_ _12793_/A _12793_/B _12793_/C _12793_/D _12793_/Y vdd gnd AOI22X1
X_14532_ _14532_/D _14532_/CLK _14532_/Q vdd gnd DFFPOSX1
X_11744_ _11744_/A _11744_/B _11744_/Y vdd gnd NOR2X1
XBUFX2_insert112 BUFX2_insert112/A BUFX2_insert112/Y vdd gnd BUFX2
XBUFX2_insert123 BUFX2_insert123/A BUFX2_insert123/Y vdd gnd BUFX2
X_14463_ _14463_/A _14463_/B _14463_/Y vdd gnd NAND2X1
XBUFX2_insert134 BUFX2_insert134/A BUFX2_insert134/Y vdd gnd BUFX2
X_11675_ _11675_/D _11675_/CLK _11675_/Q vdd gnd DFFPOSX1
XBUFX2_insert145 BUFX2_insert145/A BUFX2_insert145/Y vdd gnd BUFX2
XBUFX2_insert156 BUFX2_insert156/A BUFX2_insert156/Y vdd gnd BUFX2
X_13414_ _13414_/A _13414_/B _13414_/Y vdd gnd NAND2X1
XFILL_1__10770_ vdd gnd FILL
X_10626_ _10626_/A _10626_/B _10626_/Y vdd gnd NAND2X1
XBUFX2_insert167 BUFX2_insert167/A BUFX2_insert167/Y vdd gnd BUFX2
XBUFX2_insert178 BUFX2_insert178/A BUFX2_insert178/Y vdd gnd BUFX2
X_14394_ _14394_/A _14394_/B _14394_/C _14394_/Y vdd gnd NAND3X1
XBUFX2_insert189 BUFX2_insert189/A BUFX2_insert189/Y vdd gnd BUFX2
XFILL_1__9929_ vdd gnd FILL
XFILL_2__8722_ vdd gnd FILL
XFILL_0__11150_ vdd gnd FILL
X_13345_ _13345_/A _13345_/B _13345_/Y vdd gnd NAND2X1
X_10557_ _10557_/A _10557_/B _10557_/Y vdd gnd OR2X2
XFILL_0__10101_ vdd gnd FILL
XFILL_2__8653_ vdd gnd FILL
XFILL_1__12440_ vdd gnd FILL
XFILL_0__11081_ vdd gnd FILL
XFILL_2__11991_ vdd gnd FILL
X_13276_ _13276_/A _13276_/B _13276_/C _13276_/Y vdd gnd OAI21X1
X_10488_ _10488_/A _10488_/Y vdd gnd INVX1
XFILL_2__13730_ vdd gnd FILL
XFILL_0__10032_ vdd gnd FILL
XFILL_2__8584_ vdd gnd FILL
XFILL_1__12371_ vdd gnd FILL
X_12227_ _12227_/A _12227_/B _12227_/C _12227_/Y vdd gnd OAI21X1
XFILL_1__14110_ vdd gnd FILL
XFILL_2__13661_ vdd gnd FILL
XFILL_1__11322_ vdd gnd FILL
XFILL_0__14840_ vdd gnd FILL
X_12158_ _12158_/A _12158_/B _12158_/C _12158_/Y vdd gnd OAI21X1
XFILL_1__14041_ vdd gnd FILL
XFILL_1__11253_ vdd gnd FILL
X_11109_ _11109_/A _11109_/B _11109_/C _11109_/Y vdd gnd NAND3X1
XFILL_0__14771_ vdd gnd FILL
XFILL_2__9205_ vdd gnd FILL
XFILL_0__11983_ vdd gnd FILL
X_12089_ _12089_/A _12089_/B _12089_/C _12089_/Y vdd gnd OAI21X1
XFILL_1__10204_ vdd gnd FILL
XFILL_1__11184_ vdd gnd FILL
XFILL_0__13722_ vdd gnd FILL
XFILL_0__8220_ vdd gnd FILL
XFILL_0__10934_ vdd gnd FILL
XFILL_2__9136_ vdd gnd FILL
XFILL_1__10135_ vdd gnd FILL
XFILL_0__13653_ vdd gnd FILL
XFILL_0__8151_ vdd gnd FILL
XFILL_0__10865_ vdd gnd FILL
XFILL_2__9067_ vdd gnd FILL
XFILL_2__11425_ vdd gnd FILL
XFILL_1__10066_ vdd gnd FILL
XFILL_0__7102_ vdd gnd FILL
XFILL_0__13584_ vdd gnd FILL
XFILL_0__10796_ vdd gnd FILL
X_7730_ _7730_/A _7730_/B _7730_/Y vdd gnd NAND2X1
XFILL_0__8082_ vdd gnd FILL
XFILL_2__14144_ vdd gnd FILL
XFILL_2__11356_ vdd gnd FILL
XFILL_0__12535_ vdd gnd FILL
X_7661_ _7661_/A _7661_/Y vdd gnd INVX1
XFILL_1__13825_ vdd gnd FILL
XFILL_2__14075_ vdd gnd FILL
XFILL_2__11287_ vdd gnd FILL
X_9400_ _9400_/A _9400_/B _9400_/C _9400_/Y vdd gnd OAI21X1
XFILL_0__12466_ vdd gnd FILL
X_7592_ _7592_/A _7592_/B _7592_/C _7592_/Y vdd gnd NAND3X1
XFILL_2__9969_ vdd gnd FILL
XFILL_0__11417_ vdd gnd FILL
XFILL_1__13756_ vdd gnd FILL
XFILL_1__10968_ vdd gnd FILL
XFILL_0__12397_ vdd gnd FILL
X_9331_ _9331_/A _9331_/B _9331_/C _9331_/Y vdd gnd AOI21X1
XFILL257250x230550 vdd gnd FILL
XFILL_0__8984_ vdd gnd FILL
XFILL_1__12707_ vdd gnd FILL
XFILL_0__14136_ vdd gnd FILL
XFILL_0__11348_ vdd gnd FILL
XFILL_1__13687_ vdd gnd FILL
XFILL_1__10899_ vdd gnd FILL
X_9262_ _9262_/A _9262_/B _9262_/C _9262_/Y vdd gnd OAI21X1
XFILL_1__12638_ vdd gnd FILL
XFILL_0__14067_ vdd gnd FILL
XFILL_0__11279_ vdd gnd FILL
X_8213_ _8213_/A _8213_/Y vdd gnd INVX1
XFILL_0__7866_ vdd gnd FILL
X_9193_ _9193_/A _9193_/B _9193_/C _9193_/Y vdd gnd OAI21X1
XFILL_0__13018_ vdd gnd FILL
XFILL_0__9605_ vdd gnd FILL
X_8144_ _8144_/A _8144_/B _8144_/C _8144_/Y vdd gnd AOI21X1
XFILL_0__7797_ vdd gnd FILL
XFILL_1__14308_ vdd gnd FILL
XFILL_0__9536_ vdd gnd FILL
X_8075_ _8075_/A _8075_/Y vdd gnd INVX1
XFILL_1__14239_ vdd gnd FILL
XFILL_0__9467_ vdd gnd FILL
XFILL_1__8260_ vdd gnd FILL
XFILL_1__7211_ vdd gnd FILL
XFILL_0__8418_ vdd gnd FILL
XFILL_0__9398_ vdd gnd FILL
XFILL_1__8191_ vdd gnd FILL
XFILL_1__7142_ vdd gnd FILL
XFILL_0__8349_ vdd gnd FILL
X_8977_ _8977_/A _8977_/B _8977_/C _8977_/Y vdd gnd OAI21X1
XFILL_1_BUFX2_insert109 vdd gnd FILL
X_7928_ _7928_/D _7928_/CLK _7928_/Q vdd gnd DFFPOSX1
XFILL_1__7073_ vdd gnd FILL
X_7859_ _7859_/A _7859_/B _7859_/C _7859_/Y vdd gnd OAI21X1
XFILL257250x140550 vdd gnd FILL
X_11460_ _11460_/A _11460_/B _11460_/Y vdd gnd NAND2X1
X_9529_ _9529_/A _9529_/B _9529_/Y vdd gnd NOR2X1
X_10411_ _10411_/A _10411_/B _10411_/Y vdd gnd NAND2X1
XFILL_1__9714_ vdd gnd FILL
X_11391_ _11391_/A _11391_/B _11391_/Y vdd gnd NOR2X1
X_13130_ _13130_/A _13130_/B _13130_/C _13130_/Y vdd gnd AOI21X1
X_10342_ _10342_/A _10342_/B _10342_/C _10342_/Y vdd gnd OAI21X1
XFILL_1__9645_ vdd gnd FILL
X_13061_ _13061_/A _13061_/B _13061_/Y vdd gnd NAND2X1
X_10273_ _10273_/A _10273_/Y vdd gnd INVX1
XFILL_1__9576_ vdd gnd FILL
X_12012_ _12012_/A _12012_/B _12012_/C _12012_/Y vdd gnd OAI21X1
XFILL_2__7320_ vdd gnd FILL
XFILL_1__8527_ vdd gnd FILL
XFILL_1__8458_ vdd gnd FILL
XFILL_1__7409_ vdd gnd FILL
X_13963_ _13963_/A _13963_/B _13963_/Y vdd gnd NAND2X1
XFILL_1__8389_ vdd gnd FILL
X_12914_ _12914_/A _12914_/B _12914_/C _12914_/Y vdd gnd AOI21X1
X_13894_ _13894_/A _13894_/B _13894_/Y vdd gnd AND2X2
XFILL_0__10650_ vdd gnd FILL
X_12845_ _12845_/A _12845_/B _12845_/Y vdd gnd NAND2X1
XFILL_2__11210_ vdd gnd FILL
XFILL_1__11940_ vdd gnd FILL
XFILL_0__10581_ vdd gnd FILL
X_12776_ _12776_/A _12776_/B _12776_/C _12776_/Y vdd gnd OAI21X1
XFILL_2__11141_ vdd gnd FILL
XFILL_0__12320_ vdd gnd FILL
XFILL_1__11871_ vdd gnd FILL
X_14515_ _14515_/D _14515_/CLK _14515_/Q vdd gnd DFFPOSX1
X_11727_ _11727_/A _11727_/B _11727_/C _11727_/Y vdd gnd AOI21X1
XFILL_1__13610_ vdd gnd FILL
XFILL_2__11072_ vdd gnd FILL
XFILL_0__12251_ vdd gnd FILL
XFILL_1__10822_ vdd gnd FILL
XFILL_1__14590_ vdd gnd FILL
X_14446_ _14446_/A _14446_/B _14446_/Y vdd gnd NAND2X1
X_11658_ _11658_/D _11658_/CLK _11658_/Q vdd gnd DFFPOSX1
XFILL_1__13541_ vdd gnd FILL
XFILL_0__11202_ vdd gnd FILL
XFILL_0__12182_ vdd gnd FILL
X_10609_ _10609_/A _10609_/B _10609_/Y vdd gnd NAND2X1
X_14377_ _14377_/A _14377_/Y vdd gnd INVX1
XFILL_2__8705_ vdd gnd FILL
X_11589_ _11589_/A _11589_/B _11589_/C _11589_/Y vdd gnd OAI21X1
XFILL_0__11133_ vdd gnd FILL
XFILL_1__10684_ vdd gnd FILL
XFILL_0__7720_ vdd gnd FILL
X_13328_ _13328_/A _13328_/B _13328_/Y vdd gnd NAND2X1
XFILL_2__8636_ vdd gnd FILL
XFILL_1__12423_ vdd gnd FILL
XFILL_2__11974_ vdd gnd FILL
XFILL_0__11064_ vdd gnd FILL
XFILL_0__7651_ vdd gnd FILL
X_13259_ _13259_/A _13259_/B _13259_/Y vdd gnd NAND2X1
XFILL_0__10015_ vdd gnd FILL
XFILL_2__8567_ vdd gnd FILL
XFILL_2__13713_ vdd gnd FILL
XFILL_2__14693_ vdd gnd FILL
XFILL_1__12354_ vdd gnd FILL
XFILL_0__7582_ vdd gnd FILL
XFILL_2__13644_ vdd gnd FILL
XFILL_1__11305_ vdd gnd FILL
XFILL_0__14823_ vdd gnd FILL
XFILL_2__8498_ vdd gnd FILL
XFILL_0__9321_ vdd gnd FILL
XFILL_1__12285_ vdd gnd FILL
XFILL_1__14024_ vdd gnd FILL
XFILL_1__11236_ vdd gnd FILL
XFILL_2__13575_ vdd gnd FILL
XFILL_0__14754_ vdd gnd FILL
XFILL_0__9252_ vdd gnd FILL
XFILL_0__11966_ vdd gnd FILL
X_8900_ _8900_/D _8900_/CLK _8900_/Q vdd gnd DFFPOSX1
X_9880_ _9880_/A _9880_/Y vdd gnd INVX1
XFILL_0__13705_ vdd gnd FILL
XFILL_1__11167_ vdd gnd FILL
XFILL_0__8203_ vdd gnd FILL
XFILL_0__10917_ vdd gnd FILL
XFILL_0__14685_ vdd gnd FILL
XFILL_0__9183_ vdd gnd FILL
XFILL_0__11897_ vdd gnd FILL
X_8831_ _8831_/A _8831_/B _8831_/C _8831_/Y vdd gnd OAI21X1
XFILL_2__9119_ vdd gnd FILL
XFILL_1__10118_ vdd gnd FILL
XBUFX2_insert1 BUFX2_insert1/A BUFX2_insert1/Y vdd gnd BUFX2
XFILL_0__13636_ vdd gnd FILL
XFILL_0__8134_ vdd gnd FILL
XFILL_0__10848_ vdd gnd FILL
XFILL_1__11098_ vdd gnd FILL
X_8762_ _8762_/A _8762_/B _8762_/C _8762_/Y vdd gnd OAI21X1
XFILL_2__11408_ vdd gnd FILL
XFILL_1__10049_ vdd gnd FILL
XFILL_0__13567_ vdd gnd FILL
X_7713_ _7713_/A _7713_/B _7713_/Y vdd gnd NAND2X1
XFILL_0__8065_ vdd gnd FILL
XFILL_0__10779_ vdd gnd FILL
X_8693_ _8693_/A _8693_/B _8693_/Y vdd gnd NOR2X1
XFILL_2__11339_ vdd gnd FILL
XFILL_1__14857_ vdd gnd FILL
XFILL_0__12518_ vdd gnd FILL
X_7644_ _7644_/A _7644_/B _7644_/C _7644_/Y vdd gnd OAI21X1
XFILL_1__13808_ vdd gnd FILL
XFILL_1__14788_ vdd gnd FILL
XFILL_0__12449_ vdd gnd FILL
X_7575_ _7575_/A _7575_/B _7575_/Y vdd gnd NAND2X1
XFILL_1__13739_ vdd gnd FILL
X_9314_ _9314_/A _9314_/B _9314_/C _9314_/Y vdd gnd OAI21X1
XFILL_1__7760_ vdd gnd FILL
XFILL_0__8967_ vdd gnd FILL
XFILL_0__14119_ vdd gnd FILL
X_9245_ _9245_/A _9245_/B _9245_/C _9245_/Y vdd gnd AOI21X1
XFILL_1__7691_ vdd gnd FILL
XFILL_1__9430_ vdd gnd FILL
XFILL_0__7849_ vdd gnd FILL
X_9176_ _9176_/A _9176_/Y vdd gnd INVX1
XFILL_1__9361_ vdd gnd FILL
X_8127_ _8127_/A _8127_/B _8127_/C _8127_/Y vdd gnd OAI21X1
XFILL_1__8312_ vdd gnd FILL
XFILL_0__9519_ vdd gnd FILL
XFILL_1__9292_ vdd gnd FILL
X_8058_ _8058_/A _8058_/Y vdd gnd INVX1
XFILL_1__8243_ vdd gnd FILL
X_10960_ _10960_/A _10960_/B _10960_/Y vdd gnd NAND2X1
XFILL_1__8174_ vdd gnd FILL
XFILL_1__7125_ vdd gnd FILL
X_10891_ _10891_/A _10891_/B _10891_/C _10891_/Y vdd gnd OAI21X1
X_12630_ _12630_/A _12630_/B _12630_/C _12630_/Y vdd gnd OAI21X1
XFILL_1_CLKBUF1_insert50 vdd gnd FILL
XFILL_1_CLKBUF1_insert61 vdd gnd FILL
X_12561_ _12561_/D _12561_/CLK _12561_/Q vdd gnd DFFPOSX1
XFILL_1_CLKBUF1_insert72 vdd gnd FILL
XFILL_1_CLKBUF1_insert83 vdd gnd FILL
XFILL_1_CLKBUF1_insert94 vdd gnd FILL
X_14300_ _14300_/A _14300_/B _14300_/C _14300_/Y vdd gnd OAI21X1
X_11512_ _11512_/A _11512_/B _11512_/C _11512_/D _11512_/Y vdd gnd OAI22X1
X_12492_ _12492_/A _12492_/B _12492_/C _12492_/Y vdd gnd OAI21X1
X_14231_ _14231_/A _14231_/Y vdd gnd INVX1
X_11443_ _11443_/A _11443_/B _11443_/C _11443_/Y vdd gnd OAI21X1
X_14162_ _14162_/D _14162_/CLK _14162_/Q vdd gnd DFFPOSX1
X_11374_ _11374_/A _11374_/B _11374_/Y vdd gnd NAND2X1
XFILL_1__7889_ vdd gnd FILL
X_13113_ _13113_/A _13113_/B _13113_/C _13113_/Y vdd gnd OAI21X1
X_10325_ _10325_/A _10325_/B _10325_/Y vdd gnd NAND2X1
X_14093_ _14093_/A _14093_/B _14093_/Y vdd gnd NOR2X1
XFILL_1__9628_ vdd gnd FILL
X_13044_ _13044_/A _13044_/B _13044_/C _13044_/Y vdd gnd OAI21X1
X_10256_ _10256_/A _10256_/B _10256_/C _10256_/Y vdd gnd OAI21X1
XFILL_1__9559_ vdd gnd FILL
XFILL_2__7303_ vdd gnd FILL
X_10187_ _10187_/A _10187_/B _10187_/C _10187_/Y vdd gnd OAI21X1
XFILL_0__11820_ vdd gnd FILL
XFILL_1__12070_ vdd gnd FILL
XFILL_2__7234_ vdd gnd FILL
XFILL_1__11021_ vdd gnd FILL
XFILL_2__13360_ vdd gnd FILL
XFILL_0__11751_ vdd gnd FILL
X_13946_ _13946_/A _13946_/B _13946_/Y vdd gnd NAND2X1
XFILL_2__7165_ vdd gnd FILL
XFILL_2__13291_ vdd gnd FILL
XFILL_0__14470_ vdd gnd FILL
XFILL256650x28950 vdd gnd FILL
X_13877_ _13877_/A _13877_/B _13877_/S _13877_/Y vdd gnd MUX2X1
XFILL_2__7096_ vdd gnd FILL
XFILL_0__13421_ vdd gnd FILL
XFILL_0__10633_ vdd gnd FILL
XFILL_1__12972_ vdd gnd FILL
X_12828_ _12828_/A _12828_/B _12828_/C _12828_/Y vdd gnd NAND3X1
XFILL_1__14711_ vdd gnd FILL
XFILL_1__11923_ vdd gnd FILL
XFILL_0__13352_ vdd gnd FILL
XFILL_0__10564_ vdd gnd FILL
X_12759_ _12759_/A _12759_/Y vdd gnd INVX1
XFILL_1__14642_ vdd gnd FILL
XFILL_0__12303_ vdd gnd FILL
XFILL_1__11854_ vdd gnd FILL
XFILL_0__10495_ vdd gnd FILL
XFILL_0__13283_ vdd gnd FILL
XFILL_0__9870_ vdd gnd FILL
XFILL_2__11055_ vdd gnd FILL
XFILL_1__10805_ vdd gnd FILL
XFILL_1__14573_ vdd gnd FILL
XFILL_0__12234_ vdd gnd FILL
XFILL_2__7998_ vdd gnd FILL
XFILL_1__11785_ vdd gnd FILL
X_14429_ _14429_/A _14429_/B _14429_/C _14429_/Y vdd gnd NAND3X1
XFILL_0__8821_ vdd gnd FILL
X_7360_ _7360_/A _7360_/Y vdd gnd INVX1
XFILL_1__13524_ vdd gnd FILL
XFILL_0__12165_ vdd gnd FILL
XFILL_0__8752_ vdd gnd FILL
X_7291_ _7291_/A _7291_/B _7291_/C _7291_/Y vdd gnd NAND3X1
XFILL_0__11116_ vdd gnd FILL
XFILL_1__10667_ vdd gnd FILL
XFILL_0__7703_ vdd gnd FILL
XFILL_0__12096_ vdd gnd FILL
X_9030_ _9030_/A _9030_/Y vdd gnd INVX1
XFILL_0__8683_ vdd gnd FILL
XFILL_1__12406_ vdd gnd FILL
XFILL_0__11047_ vdd gnd FILL
XFILL_1__13386_ vdd gnd FILL
XFILL_0__7634_ vdd gnd FILL
XFILL_1__10598_ vdd gnd FILL
XFILL_2__10908_ vdd gnd FILL
XFILL_1__12337_ vdd gnd FILL
XFILL_2__11888_ vdd gnd FILL
XFILL_0__7565_ vdd gnd FILL
XFILL_0__14806_ vdd gnd FILL
XFILL_2__10839_ vdd gnd FILL
XFILL_2__13627_ vdd gnd FILL
XFILL_1__12268_ vdd gnd FILL
XFILL_0__9304_ vdd gnd FILL
X_9932_ _9932_/A _9932_/B _9932_/S _9932_/Y vdd gnd MUX2X1
XFILL_0__12998_ vdd gnd FILL
XFILL_1__14007_ vdd gnd FILL
XFILL_0__7496_ vdd gnd FILL
XFILL_1__11219_ vdd gnd FILL
XFILL_2__13558_ vdd gnd FILL
XFILL_0__14737_ vdd gnd FILL
XFILL_0__9235_ vdd gnd FILL
XFILL_0__11949_ vdd gnd FILL
XFILL_1__12199_ vdd gnd FILL
X_9863_ _9863_/A _9863_/B _9863_/Y vdd gnd NAND2X1
XFILL_0__14668_ vdd gnd FILL
XFILL_0__9166_ vdd gnd FILL
X_8814_ _8814_/A _8814_/B _8814_/Y vdd gnd NAND2X1
X_9794_ _9794_/D _9794_/CLK _9794_/Q vdd gnd DFFPOSX1
XFILL_0__13619_ vdd gnd FILL
XFILL_0__8117_ vdd gnd FILL
XFILL_0__14599_ vdd gnd FILL
XFILL_0__9097_ vdd gnd FILL
X_8745_ _8745_/A _8745_/B _8745_/C _8745_/Y vdd gnd AOI21X1
XFILL_1__14909_ vdd gnd FILL
XFILL_0__8048_ vdd gnd FILL
XFILL_1__8930_ vdd gnd FILL
X_8676_ _8676_/A _8676_/B _8676_/Y vdd gnd OR2X2
X_7627_ _7627_/A _7627_/B _7627_/C _7627_/Y vdd gnd NAND3X1
XFILL_1_CLKBUF1_insert105 vdd gnd FILL
XFILL_1__7812_ vdd gnd FILL
X_7558_ _7558_/A _7558_/Y vdd gnd INVX1
XFILL_1__8792_ vdd gnd FILL
XFILL_0__9999_ vdd gnd FILL
XFILL_1__7743_ vdd gnd FILL
X_7489_ _7489_/A _7489_/B _7489_/C _7489_/Y vdd gnd OAI21X1
X_9228_ _9228_/A _9228_/Y vdd gnd INVX1
XFILL_1__7674_ vdd gnd FILL
X_10110_ _10110_/A _10110_/B _10110_/C _10110_/Y vdd gnd NAND3X1
XFILL_1__9413_ vdd gnd FILL
X_11090_ _11090_/A _11090_/Y vdd gnd INVX1
X_9159_ _9159_/A _9159_/B _9159_/Y vdd gnd NAND2X1
X_10041_ _10041_/A _10041_/B _10041_/Y vdd gnd NOR2X1
XFILL_1__9344_ vdd gnd FILL
XFILL_1__9275_ vdd gnd FILL
X_13800_ _13800_/A _13800_/B _13800_/C _13800_/Y vdd gnd NAND3X1
XFILL_1__8226_ vdd gnd FILL
X_14780_ _14780_/A _14780_/B _14780_/C _14780_/Y vdd gnd OAI21X1
X_11992_ _11992_/A _11992_/B _11992_/Y vdd gnd AND2X2
X_13731_ _13731_/A _13731_/B _13731_/Y vdd gnd NAND2X1
X_10943_ _10943_/A _10943_/Y vdd gnd INVX1
XFILL_1__8157_ vdd gnd FILL
XFILL_1__7108_ vdd gnd FILL
X_13662_ _13662_/A _13662_/Y vdd gnd INVX1
X_10874_ _10874_/A _10874_/B _10874_/S _10874_/Y vdd gnd MUX2X1
XFILL_1__8088_ vdd gnd FILL
X_12613_ _12613_/D _12613_/CLK _12613_/Q vdd gnd DFFPOSX1
X_13593_ _13593_/A _13593_/Y vdd gnd INVX1
X_12544_ _12544_/D _12544_/CLK _12544_/Q vdd gnd DFFPOSX1
XFILL_0__10280_ vdd gnd FILL
X_12475_ _12475_/A _12475_/B _12475_/C _12475_/Y vdd gnd OAI21X1
XFILL_1__11570_ vdd gnd FILL
X_14214_ _14214_/D _14214_/CLK _14214_/Q vdd gnd DFFPOSX1
X_11426_ _11426_/A _11426_/B _11426_/Y vdd gnd NAND2X1
XFILL_2__9522_ vdd gnd FILL
XFILL_1__10521_ vdd gnd FILL
XFILL_2__12860_ vdd gnd FILL
X_14145_ _14145_/A _14145_/B _14145_/Y vdd gnd NAND2X1
X_11357_ _11357_/A _11357_/Y vdd gnd INVX1
XFILL_2__9453_ vdd gnd FILL
XFILL_1__13240_ vdd gnd FILL
XFILL_1__10452_ vdd gnd FILL
XCLKBUF1_insert104 CLKBUF1_insert104/A CLKBUF1_insert104/Y vdd gnd CLKBUF1
XFILL_2__12791_ vdd gnd FILL
XFILL_0__13970_ vdd gnd FILL
X_10308_ _10308_/A _10308_/Y vdd gnd INVX1
X_14076_ _14076_/A _14076_/B _14076_/Y vdd gnd OR2X2
X_11288_ _11288_/A _11288_/B _11288_/C _11288_/Y vdd gnd NAND3X1
XFILL_1__13171_ vdd gnd FILL
XFILL_0__12921_ vdd gnd FILL
XFILL_2__9384_ vdd gnd FILL
XFILL_1__10383_ vdd gnd FILL
X_13027_ _13027_/A _13027_/B _13027_/Y vdd gnd NAND2X1
X_10239_ _10239_/A _10239_/Y vdd gnd INVX1
XFILL_2__14461_ vdd gnd FILL
XFILL_1__12122_ vdd gnd FILL
XFILL_0__12852_ vdd gnd FILL
XFILL_0__7350_ vdd gnd FILL
XFILL_1__12053_ vdd gnd FILL
XFILL_2__14392_ vdd gnd FILL
XFILL_0__11803_ vdd gnd FILL
XFILL_0__12783_ vdd gnd FILL
XFILL_2__7217_ vdd gnd FILL
XFILL_0__7281_ vdd gnd FILL
XFILL_1__11004_ vdd gnd FILL
XFILL_2__13343_ vdd gnd FILL
XFILL_0__9020_ vdd gnd FILL
XFILL_0__11734_ vdd gnd FILL
X_13929_ _13929_/A _13929_/B _13929_/Y vdd gnd NAND2X1
XFILL_2__7148_ vdd gnd FILL
XFILL_2__13274_ vdd gnd FILL
XFILL_0__14453_ vdd gnd FILL
XFILL_2__7079_ vdd gnd FILL
XFILL_0__13404_ vdd gnd FILL
XFILL_1__12955_ vdd gnd FILL
XFILL_0__10616_ vdd gnd FILL
XFILL_0__14384_ vdd gnd FILL
XFILL_1_BUFX2_insert270 vdd gnd FILL
X_8530_ _8530_/A _8530_/Y vdd gnd INVX1
XFILL_0__11596_ vdd gnd FILL
XCLKBUF1_insert30 CLKBUF1_insert30/A CLKBUF1_insert30/Y vdd gnd CLKBUF1
XFILL_1_BUFX2_insert281 vdd gnd FILL
XCLKBUF1_insert41 CLKBUF1_insert41/A CLKBUF1_insert41/Y vdd gnd CLKBUF1
XFILL_1__11906_ vdd gnd FILL
XFILL_1_BUFX2_insert292 vdd gnd FILL
XCLKBUF1_insert52 CLKBUF1_insert52/A CLKBUF1_insert52/Y vdd gnd CLKBUF1
XFILL_0__13335_ vdd gnd FILL
XFILL_0__10547_ vdd gnd FILL
XCLKBUF1_insert63 CLKBUF1_insert63/A CLKBUF1_insert63/Y vdd gnd CLKBUF1
XFILL_1__12886_ vdd gnd FILL
XFILL_0__9922_ vdd gnd FILL
XCLKBUF1_insert74 CLKBUF1_insert74/A CLKBUF1_insert74/Y vdd gnd CLKBUF1
X_8461_ _8461_/A _8461_/B _8461_/C _8461_/Y vdd gnd NAND3X1
XFILL_1__14625_ vdd gnd FILL
XCLKBUF1_insert85 CLKBUF1_insert85/A CLKBUF1_insert85/Y vdd gnd CLKBUF1
XCLKBUF1_insert96 CLKBUF1_insert96/A CLKBUF1_insert96/Y vdd gnd CLKBUF1
XFILL_1__11837_ vdd gnd FILL
XFILL_0__13266_ vdd gnd FILL
X_7412_ _7412_/A _7412_/B _7412_/Y vdd gnd AND2X2
XFILL_0__10478_ vdd gnd FILL
XFILL_0__9853_ vdd gnd FILL
X_8392_ _8392_/A _8392_/B _8392_/Y vdd gnd NAND2X1
XFILL_1__14556_ vdd gnd FILL
XFILL_0__12217_ vdd gnd FILL
XFILL_1__11768_ vdd gnd FILL
XFILL_0__13197_ vdd gnd FILL
XFILL_0__8804_ vdd gnd FILL
X_7343_ _7343_/A _7343_/Y vdd gnd INVX1
XFILL_1__13507_ vdd gnd FILL
XFILL_1__14487_ vdd gnd FILL
XFILL_0__12148_ vdd gnd FILL
XFILL_1__11699_ vdd gnd FILL
XFILL_0__8735_ vdd gnd FILL
X_7274_ _7274_/A _7274_/B _7274_/C _7274_/Y vdd gnd OAI21X1
XFILL_0__12079_ vdd gnd FILL
X_9013_ _9013_/A _9013_/B _9013_/C _9013_/Y vdd gnd AOI21X1
XFILL_0__8666_ vdd gnd FILL
XFILL_1__13369_ vdd gnd FILL
XFILL_0__7617_ vdd gnd FILL
XFILL_1__7390_ vdd gnd FILL
XFILL_0__8597_ vdd gnd FILL
XFILL_0__7548_ vdd gnd FILL
XFILL_1__9060_ vdd gnd FILL
XFILL_0__7479_ vdd gnd FILL
X_9915_ _9915_/A _9915_/B _9915_/C _9915_/Y vdd gnd OAI21X1
XFILL_1__8011_ vdd gnd FILL
XFILL_0__9218_ vdd gnd FILL
X_9846_ _9846_/A _9846_/B _9846_/Y vdd gnd NOR2X1
XFILL_0__9149_ vdd gnd FILL
X_9777_ _9777_/D _9777_/CLK _9777_/Q vdd gnd DFFPOSX1
X_8728_ _8728_/A _8728_/B _8728_/C _8728_/Y vdd gnd NAND3X1
XFILL_1__9962_ vdd gnd FILL
X_10590_ _10590_/A _10590_/B _10590_/C _10590_/Y vdd gnd OAI21X1
X_8659_ _8659_/A _8659_/B _8659_/Y vdd gnd NOR2X1
XFILL_1__9893_ vdd gnd FILL
X_12260_ _12260_/A _12260_/B _12260_/Y vdd gnd NOR2X1
XFILL_1__8775_ vdd gnd FILL
X_11211_ _11211_/A _11211_/B _11211_/Y vdd gnd NAND2X1
X_12191_ _12191_/A _12191_/B _12191_/C _12191_/Y vdd gnd OAI21X1
XFILL_1__7726_ vdd gnd FILL
X_11142_ _11142_/A _11142_/B _11142_/C _11142_/Y vdd gnd OAI21X1
XFILL_1__7657_ vdd gnd FILL
X_11073_ _11073_/A _11073_/B _11073_/C _11073_/Y vdd gnd AOI21X1
XFILL_1__7588_ vdd gnd FILL
X_14901_ _14901_/D _14901_/CLK _14901_/Q vdd gnd DFFPOSX1
X_10024_ _10024_/A _10024_/Y vdd gnd INVX1
XFILL_1__9327_ vdd gnd FILL
X_14832_ _14832_/A _14832_/Y vdd gnd INVX1
XFILL_1__9258_ vdd gnd FILL
X_14763_ _14763_/A _14763_/B _14763_/Y vdd gnd NOR2X1
XFILL_1__8209_ vdd gnd FILL
XFILL_1__9189_ vdd gnd FILL
X_11975_ _11975_/A _11975_/Y vdd gnd INVX1
X_13714_ _13714_/A _13714_/Y vdd gnd INVX1
X_10926_ _10926_/A _10926_/B _10926_/C _10926_/Y vdd gnd OAI21X1
X_14694_ _14694_/A _14694_/B _14694_/Y vdd gnd NAND2X1
XFILL_0__11450_ vdd gnd FILL
XFILL_2__12010_ vdd gnd FILL
X_13645_ _13645_/A _13645_/Y vdd gnd INVX1
X_10857_ _10857_/A _10857_/B _10857_/S _10857_/Y vdd gnd MUX2X1
XFILL_0__10401_ vdd gnd FILL
XFILL_0_BUFX2_insert200 vdd gnd FILL
XFILL_1__12740_ vdd gnd FILL
XFILL_0_BUFX2_insert211 vdd gnd FILL
XFILL_0__11381_ vdd gnd FILL
XFILL_0_BUFX2_insert222 vdd gnd FILL
XFILL_0_BUFX2_insert233 vdd gnd FILL
X_10788_ _10788_/A _10788_/B _10788_/C _10788_/Y vdd gnd OAI21X1
X_13576_ _13576_/A _13576_/B _13576_/S _13576_/Y vdd gnd MUX2X1
XFILL_0__13120_ vdd gnd FILL
XFILL_0_BUFX2_insert244 vdd gnd FILL
XFILL_0__10332_ vdd gnd FILL
XFILL_0_BUFX2_insert255 vdd gnd FILL
XFILL_1__12671_ vdd gnd FILL
XFILL_0_BUFX2_insert266 vdd gnd FILL
X_12527_ _12527_/A _12527_/B _12527_/C _12527_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert277 vdd gnd FILL
XFILL_1__14410_ vdd gnd FILL
XFILL_0_BUFX2_insert288 vdd gnd FILL
XFILL_2__13961_ vdd gnd FILL
XFILL_0__10263_ vdd gnd FILL
XFILL_0_BUFX2_insert299 vdd gnd FILL
XFILL_0__13051_ vdd gnd FILL
X_12458_ _12458_/A _12458_/B _12458_/C _12458_/Y vdd gnd OAI21X1
XFILL_0__12002_ vdd gnd FILL
XFILL_1__14341_ vdd gnd FILL
XFILL_2__12912_ vdd gnd FILL
XFILL_1__11553_ vdd gnd FILL
XFILL_2__13892_ vdd gnd FILL
XFILL_0__10194_ vdd gnd FILL
X_11409_ _11409_/A _11409_/B _11409_/Y vdd gnd NAND2X1
XFILL_2__9505_ vdd gnd FILL
X_12389_ _12389_/A _12389_/B _12389_/Y vdd gnd NOR2X1
XFILL_1__10504_ vdd gnd FILL
XFILL_2_BUFX2_insert15 vdd gnd FILL
XFILL_1__14272_ vdd gnd FILL
XFILL_2__12843_ vdd gnd FILL
XFILL_1__11484_ vdd gnd FILL
XFILL_0__8520_ vdd gnd FILL
X_14128_ _14128_/A _14128_/B _14128_/C _14128_/Y vdd gnd OAI21X1
XFILL_2__9436_ vdd gnd FILL
XFILL_1__13223_ vdd gnd FILL
XFILL_1__10435_ vdd gnd FILL
XFILL_2__12774_ vdd gnd FILL
XFILL_0__13953_ vdd gnd FILL
XFILL_0__8451_ vdd gnd FILL
X_14059_ _14059_/A _14059_/B _14059_/Y vdd gnd NAND2X1
XFILL_1__13154_ vdd gnd FILL
XFILL_0__12904_ vdd gnd FILL
XFILL_2__9367_ vdd gnd FILL
XFILL_1__10366_ vdd gnd FILL
XFILL_0__7402_ vdd gnd FILL
XFILL_0__13884_ vdd gnd FILL
XFILL_0__8382_ vdd gnd FILL
XFILL_1__12105_ vdd gnd FILL
XFILL_2__14444_ vdd gnd FILL
XFILL_1__13085_ vdd gnd FILL
XFILL_2__9298_ vdd gnd FILL
XFILL_0__12835_ vdd gnd FILL
XFILL_0__7333_ vdd gnd FILL
XFILL_1__10297_ vdd gnd FILL
X_7961_ _7961_/D _7961_/CLK _7961_/Q vdd gnd DFFPOSX1
XFILL_1__12036_ vdd gnd FILL
XFILL_2__14375_ vdd gnd FILL
XFILL_2__11587_ vdd gnd FILL
X_9700_ _9700_/A _9700_/B _9700_/Y vdd gnd NAND2X1
XFILL_0__12766_ vdd gnd FILL
XFILL_0__7264_ vdd gnd FILL
X_7892_ _7892_/A _7892_/B _7892_/Y vdd gnd NAND2X1
XFILL_0__9003_ vdd gnd FILL
XFILL_0__11717_ vdd gnd FILL
X_9631_ _9631_/A _9631_/Y vdd gnd INVX1
XFILL_0__12697_ vdd gnd FILL
XFILL_0__7195_ vdd gnd FILL
XFILL_0__14436_ vdd gnd FILL
XFILL_1__13987_ vdd gnd FILL
X_9562_ _9562_/A _9562_/B _9562_/Y vdd gnd OR2X2
XFILL_2__12208_ vdd gnd FILL
XFILL_1__12938_ vdd gnd FILL
XFILL_0__14367_ vdd gnd FILL
X_8513_ _8513_/A _8513_/B _8513_/Y vdd gnd NOR2X1
XFILL_0__11579_ vdd gnd FILL
X_9493_ _9493_/A _9493_/B _9493_/Y vdd gnd NAND2X1
XFILL_2__12139_ vdd gnd FILL
XFILL_0__13318_ vdd gnd FILL
XFILL_1__12869_ vdd gnd FILL
XFILL_0__9905_ vdd gnd FILL
XFILL_0__14298_ vdd gnd FILL
X_8444_ _8444_/A _8444_/B _8444_/C _8444_/Y vdd gnd OAI21X1
XFILL_1__14608_ vdd gnd FILL
XFILL_0__13249_ vdd gnd FILL
X_8375_ _8375_/A _8375_/B _8375_/Y vdd gnd NAND2X1
X_7326_ _7326_/A _7326_/B _7326_/C _7326_/Y vdd gnd OAI21X1
XFILL_1__8560_ vdd gnd FILL
XFILL_1__7511_ vdd gnd FILL
XFILL_0__8718_ vdd gnd FILL
X_7257_ _7257_/A _7257_/B _7257_/C _7257_/Y vdd gnd AOI21X1
XFILL_1__8491_ vdd gnd FILL
XFILL_0__9698_ vdd gnd FILL
XFILL_1__7442_ vdd gnd FILL
XFILL_0__8649_ vdd gnd FILL
X_7188_ _7188_/A _7188_/B _7188_/S _7188_/Y vdd gnd MUX2X1
XFILL_1__7373_ vdd gnd FILL
XFILL_1_BUFX2_insert1 vdd gnd FILL
XFILL_2_BUFX2_insert306 vdd gnd FILL
XFILL_1__9112_ vdd gnd FILL
XFILL_2_BUFX2_insert339 vdd gnd FILL
XFILL_1__9043_ vdd gnd FILL
X_11760_ _11760_/A _11760_/B _11760_/S _11760_/Y vdd gnd MUX2X1
X_9829_ _9829_/D _9829_/CLK _9829_/Q vdd gnd DFFPOSX1
X_10711_ _10711_/D _10711_/CLK _10711_/Q vdd gnd DFFPOSX1
X_11691_ _11691_/D _11691_/CLK _11691_/Q vdd gnd DFFPOSX1
XBUFX2_insert305 BUFX2_insert305/A BUFX2_insert305/Y vdd gnd BUFX2
XBUFX2_insert316 BUFX2_insert316/A BUFX2_insert316/Y vdd gnd BUFX2
X_10642_ _10642_/A _10642_/B _10642_/C _10642_/Y vdd gnd OAI21X1
X_13430_ _13430_/D _13430_/CLK _13430_/Q vdd gnd DFFPOSX1
XBUFX2_insert327 BUFX2_insert327/A BUFX2_insert327/Y vdd gnd BUFX2
XBUFX2_insert338 BUFX2_insert338/A BUFX2_insert338/Y vdd gnd BUFX2
XBUFX2_insert349 BUFX2_insert349/A BUFX2_insert349/Y vdd gnd BUFX2
XFILL_1__9945_ vdd gnd FILL
X_13361_ _13361_/A _13361_/B _13361_/Y vdd gnd NAND2X1
X_10573_ _10573_/A _10573_/B _10573_/C _10573_/Y vdd gnd OAI21X1
XFILL_1__9876_ vdd gnd FILL
X_12312_ _12312_/A _12312_/B _12312_/C _12312_/Y vdd gnd OAI21X1
X_13292_ _13292_/A _13292_/B _13292_/C _13292_/Y vdd gnd OAI21X1
XFILL_2__7620_ vdd gnd FILL
XFILL_1__8827_ vdd gnd FILL
X_12243_ _12243_/A _12243_/B _12243_/C _12243_/Y vdd gnd NAND3X1
XFILL_2__7551_ vdd gnd FILL
XFILL_1__8758_ vdd gnd FILL
X_12174_ _12174_/A _12174_/B _12174_/Y vdd gnd NOR2X1
XFILL_1__7709_ vdd gnd FILL
XFILL_2__7482_ vdd gnd FILL
XFILL_1__8689_ vdd gnd FILL
X_11125_ _11125_/A _11125_/B _11125_/C _11125_/Y vdd gnd NOR3X1
XFILL_1__10220_ vdd gnd FILL
XFILL_0__10950_ vdd gnd FILL
X_11056_ _11056_/A _11056_/Y vdd gnd INVX1
XFILL_2__9152_ vdd gnd FILL
XFILL_1__10151_ vdd gnd FILL
X_10007_ _10007_/A _10007_/Y vdd gnd INVX1
XFILL_0__10881_ vdd gnd FILL
XFILL_2__8103_ vdd gnd FILL
XFILL_2__9083_ vdd gnd FILL
XFILL_2__11441_ vdd gnd FILL
XFILL_0__12620_ vdd gnd FILL
XFILL_1__10082_ vdd gnd FILL
X_14815_ _14815_/A _14815_/B _14815_/C _14815_/Y vdd gnd OAI21X1
XFILL_1__13910_ vdd gnd FILL
XFILL_2__11372_ vdd gnd FILL
X_14746_ _14746_/A _14746_/B _14746_/Y vdd gnd AND2X2
X_11958_ _11958_/A _11958_/B _11958_/C _11958_/Y vdd gnd NAND3X1
XFILL_0__11502_ vdd gnd FILL
XFILL_1__13841_ vdd gnd FILL
XFILL_0__12482_ vdd gnd FILL
X_10909_ _10909_/A _10909_/B _10909_/C _10909_/D _10909_/Y vdd gnd OAI22X1
X_14677_ _14677_/A _14677_/B _14677_/C _14677_/Y vdd gnd AOI21X1
X_11889_ _11889_/A _11889_/B _11889_/Y vdd gnd NOR2X1
XFILL_0__14221_ vdd gnd FILL
XFILL_0__11433_ vdd gnd FILL
XFILL_1__13772_ vdd gnd FILL
XFILL_1__10984_ vdd gnd FILL
X_13628_ _13628_/A _13628_/B _13628_/C _13628_/Y vdd gnd AOI21X1
XFILL_2__8936_ vdd gnd FILL
XFILL_1__12723_ vdd gnd FILL
XFILL_0__14152_ vdd gnd FILL
XFILL_0__11364_ vdd gnd FILL
X_13559_ _13559_/A _13559_/B _13559_/Y vdd gnd NAND2X1
XFILL_0__13103_ vdd gnd FILL
XFILL_1__12654_ vdd gnd FILL
XFILL_0__10315_ vdd gnd FILL
XFILL_0__14083_ vdd gnd FILL
XFILL_0__11295_ vdd gnd FILL
XFILL_0__7882_ vdd gnd FILL
XFILL_2__7818_ vdd gnd FILL
XFILL256950x72150 vdd gnd FILL
XFILL_1__11605_ vdd gnd FILL
XFILL_0__13034_ vdd gnd FILL
XFILL_2__13944_ vdd gnd FILL
XFILL_0__10246_ vdd gnd FILL
XFILL_2__8798_ vdd gnd FILL
XFILL_0__9621_ vdd gnd FILL
X_8160_ _8160_/A _8160_/B _8160_/C _8160_/Y vdd gnd NAND3X1
XFILL_1__14324_ vdd gnd FILL
XFILL_2__7749_ vdd gnd FILL
XFILL_1__11536_ vdd gnd FILL
XFILL_2__13875_ vdd gnd FILL
X_7111_ _7111_/A _7111_/B _7111_/C _7111_/Y vdd gnd OAI21X1
XFILL_0__10177_ vdd gnd FILL
XFILL_0__9552_ vdd gnd FILL
X_8091_ _8091_/A _8091_/B _8091_/C _8091_/Y vdd gnd NAND3X1
XFILL_1__14255_ vdd gnd FILL
XFILL_2__12826_ vdd gnd FILL
XFILL_1__11467_ vdd gnd FILL
XFILL256950x244950 vdd gnd FILL
XFILL_0__8503_ vdd gnd FILL
XFILL_1__13206_ vdd gnd FILL
XFILL_2__9419_ vdd gnd FILL
XFILL_0__9483_ vdd gnd FILL
XFILL_1__10418_ vdd gnd FILL
XFILL_0__13936_ vdd gnd FILL
XFILL_2__12757_ vdd gnd FILL
XFILL_1__11398_ vdd gnd FILL
XFILL_0__8434_ vdd gnd FILL
XFILL_1__13137_ vdd gnd FILL
XFILL_1__10349_ vdd gnd FILL
XFILL_0__13867_ vdd gnd FILL
XFILL_2__12688_ vdd gnd FILL
XFILL_0__8365_ vdd gnd FILL
X_8993_ _8993_/A _8993_/B _8993_/Y vdd gnd NAND2X1
XFILL_0__12818_ vdd gnd FILL
XFILL_1__13068_ vdd gnd FILL
XFILL_0__7316_ vdd gnd FILL
XFILL_0__13798_ vdd gnd FILL
X_7944_ _7944_/D _7944_/CLK _7944_/Q vdd gnd DFFPOSX1
XFILL_0__8296_ vdd gnd FILL
XFILL_1__12019_ vdd gnd FILL
XFILL_0__12749_ vdd gnd FILL
XFILL_0__7247_ vdd gnd FILL
X_7875_ _7875_/A _7875_/B _7875_/C _7875_/Y vdd gnd OAI21X1
XFILL_0__7178_ vdd gnd FILL
X_9614_ _9614_/A _9614_/Y vdd gnd INVX1
XFILL_0__14419_ vdd gnd FILL
X_9545_ _9545_/A _9545_/B _9545_/Y vdd gnd NOR2X1
XFILL_1__9730_ vdd gnd FILL
X_9476_ _9476_/A _9476_/B _9476_/C _9476_/Y vdd gnd OAI21X1
X_8427_ _8427_/A _8427_/B _8427_/Y vdd gnd NOR2X1
XFILL_1__9661_ vdd gnd FILL
XFILL_1__8612_ vdd gnd FILL
X_8358_ _8358_/A _8358_/B _8358_/Y vdd gnd NAND2X1
XFILL_1__9592_ vdd gnd FILL
X_7309_ _7309_/A _7309_/B _7309_/C _7309_/Y vdd gnd NAND3X1
XFILL_1__8543_ vdd gnd FILL
X_8289_ _8289_/A _8289_/B _8289_/C _8289_/Y vdd gnd NAND3X1
XFILL_1__8474_ vdd gnd FILL
XFILL_1__7425_ vdd gnd FILL
X_12930_ _12930_/A _12930_/B _12930_/C _12930_/Y vdd gnd OAI21X1
XFILL_2_BUFX2_insert125 vdd gnd FILL
XFILL_1__7356_ vdd gnd FILL
XFILL_2_BUFX2_insert158 vdd gnd FILL
X_12861_ _12861_/A _12861_/B _12861_/C _12861_/Y vdd gnd NAND3X1
XFILL_1__7287_ vdd gnd FILL
X_14600_ _14600_/A _14600_/B _14600_/Y vdd gnd NAND2X1
X_11812_ _11812_/A _11812_/B _11812_/S _11812_/Y vdd gnd MUX2X1
XFILL_1__9026_ vdd gnd FILL
X_12792_ _12792_/A _12792_/B _12792_/C _12792_/Y vdd gnd OAI21X1
X_14531_ _14531_/D _14531_/CLK _14531_/Q vdd gnd DFFPOSX1
X_11743_ _11743_/A _11743_/Y vdd gnd INVX1
XBUFX2_insert113 BUFX2_insert113/A BUFX2_insert113/Y vdd gnd BUFX2
X_14462_ _14462_/A _14462_/B _14462_/C _14462_/Y vdd gnd OAI21X1
XBUFX2_insert124 BUFX2_insert124/A BUFX2_insert124/Y vdd gnd BUFX2
X_11674_ _11674_/D _11674_/CLK _11674_/Q vdd gnd DFFPOSX1
XBUFX2_insert135 BUFX2_insert135/A BUFX2_insert135/Y vdd gnd BUFX2
XBUFX2_insert146 BUFX2_insert146/A BUFX2_insert146/Y vdd gnd BUFX2
XBUFX2_insert157 BUFX2_insert157/A BUFX2_insert157/Y vdd gnd BUFX2
X_13413_ _13413_/A _13413_/B _13413_/C _13413_/Y vdd gnd OAI21X1
X_10625_ _10625_/A _10625_/B _10625_/C _10625_/Y vdd gnd OAI21X1
XBUFX2_insert168 BUFX2_insert168/A BUFX2_insert168/Y vdd gnd BUFX2
XFILL_1__9928_ vdd gnd FILL
X_14393_ _14393_/A _14393_/B _14393_/Y vdd gnd NAND2X1
XBUFX2_insert179 BUFX2_insert179/A BUFX2_insert179/Y vdd gnd BUFX2
X_10556_ _10556_/A _10556_/B _10556_/Y vdd gnd NAND2X1
X_13344_ _13344_/A _13344_/B _13344_/Y vdd gnd NAND2X1
XFILL_0__10100_ vdd gnd FILL
XFILL_1__9859_ vdd gnd FILL
XFILL_0__11080_ vdd gnd FILL
XFILL_2__7603_ vdd gnd FILL
X_10487_ _10487_/A _10487_/B _10487_/Y vdd gnd NAND2X1
X_13275_ _13275_/A _13275_/B _13275_/C _13275_/Y vdd gnd OAI21X1
XFILL_2__10941_ vdd gnd FILL
XFILL_0__10031_ vdd gnd FILL
XFILL_1__12370_ vdd gnd FILL
X_12226_ _12226_/A _12226_/Y vdd gnd INVX1
XFILL_1__11321_ vdd gnd FILL
XFILL_2__7534_ vdd gnd FILL
XFILL_2__10872_ vdd gnd FILL
X_12157_ _12157_/A _12157_/B _12157_/C _12157_/Y vdd gnd NAND3X1
XFILL_1__14040_ vdd gnd FILL
XFILL_1__11252_ vdd gnd FILL
XFILL_2__7465_ vdd gnd FILL
XFILL_2__13591_ vdd gnd FILL
XFILL_0__14770_ vdd gnd FILL
X_11108_ _11108_/A _11108_/B _11108_/Y vdd gnd AND2X2
XFILL_0__11982_ vdd gnd FILL
X_12088_ _12088_/A _12088_/B _12088_/Y vdd gnd NAND2X1
XFILL_1__10203_ vdd gnd FILL
XFILL_0__13721_ vdd gnd FILL
XFILL_2__7396_ vdd gnd FILL
XFILL_0__10933_ vdd gnd FILL
XFILL_1__11183_ vdd gnd FILL
X_11039_ _11039_/A _11039_/Y vdd gnd INVX1
XFILL_1__10134_ vdd gnd FILL
XFILL_0__13652_ vdd gnd FILL
XFILL_0__8150_ vdd gnd FILL
XFILL_0__10864_ vdd gnd FILL
XFILL_0__7101_ vdd gnd FILL
XFILL_1__10065_ vdd gnd FILL
XFILL_0__13583_ vdd gnd FILL
XFILL_0__8081_ vdd gnd FILL
XFILL_0__10795_ vdd gnd FILL
XFILL_2__8017_ vdd gnd FILL
XFILL_0__12534_ vdd gnd FILL
X_14729_ _14729_/A _14729_/Y vdd gnd INVX1
XFILL_2__10306_ vdd gnd FILL
X_7660_ _7660_/A _7660_/B _7660_/C _7660_/Y vdd gnd OAI21X1
XFILL_1__13824_ vdd gnd FILL
XFILL_0__12465_ vdd gnd FILL
X_7591_ _7591_/A _7591_/B _7591_/Y vdd gnd AND2X2
XFILL_2__10237_ vdd gnd FILL
XFILL_0__11416_ vdd gnd FILL
XFILL_1__10967_ vdd gnd FILL
XFILL_1__13755_ vdd gnd FILL
X_9330_ _9330_/A _9330_/B _9330_/Y vdd gnd OR2X2
XFILL_0__12396_ vdd gnd FILL
XFILL_0__8983_ vdd gnd FILL
XFILL_2__10168_ vdd gnd FILL
XFILL_1__12706_ vdd gnd FILL
XFILL_0__14135_ vdd gnd FILL
XFILL_0__11347_ vdd gnd FILL
XFILL_1__13686_ vdd gnd FILL
XFILL_1__10898_ vdd gnd FILL
X_9261_ _9261_/A _9261_/B _9261_/C _9261_/Y vdd gnd NAND3X1
XFILL_1__12637_ vdd gnd FILL
XFILL_0__14066_ vdd gnd FILL
X_8212_ _8212_/A _8212_/B _8212_/C _8212_/Y vdd gnd NOR3X1
XFILL_0__11278_ vdd gnd FILL
X_9192_ _9192_/A _9192_/B _9192_/Y vdd gnd NOR2X1
XFILL_0__7865_ vdd gnd FILL
XFILL_2__13927_ vdd gnd FILL
XFILL_0__13017_ vdd gnd FILL
XFILL_0__10229_ vdd gnd FILL
XFILL_0__9604_ vdd gnd FILL
X_8143_ _8143_/A _8143_/B _8143_/Y vdd gnd NAND2X1
XFILL_0__7796_ vdd gnd FILL
XFILL_1__14307_ vdd gnd FILL
XFILL_1__11519_ vdd gnd FILL
XFILL_2__13858_ vdd gnd FILL
XFILL_1__12499_ vdd gnd FILL
XFILL_0__9535_ vdd gnd FILL
X_8074_ _8074_/A _8074_/B _8074_/Y vdd gnd NAND2X1
XFILL_1__14238_ vdd gnd FILL
XFILL_2__13789_ vdd gnd FILL
XFILL_0__9466_ vdd gnd FILL
XFILL_0__13919_ vdd gnd FILL
XFILL_1__7210_ vdd gnd FILL
XFILL_0__8417_ vdd gnd FILL
XFILL_1__8190_ vdd gnd FILL
XFILL_0__9397_ vdd gnd FILL
XFILL_1__7141_ vdd gnd FILL
XFILL_0__8348_ vdd gnd FILL
X_8976_ _8976_/A _8976_/B _8976_/C _8976_/D _8976_/Y vdd gnd AOI22X1
XFILL_1__7072_ vdd gnd FILL
X_7927_ _7927_/D _7927_/CLK _7927_/Q vdd gnd DFFPOSX1
XFILL_0__8279_ vdd gnd FILL
X_7858_ _7858_/A _7858_/B _7858_/C _7858_/Y vdd gnd OAI21X1
X_7789_ _7789_/A _7789_/B _7789_/Y vdd gnd NAND2X1
X_9528_ _9528_/A _9528_/B _9528_/C _9528_/Y vdd gnd AOI21X1
X_10410_ _10410_/A _10410_/B _10410_/C _10410_/D _10410_/Y vdd gnd OAI22X1
XFILL_1__9713_ vdd gnd FILL
X_11390_ _11390_/A _11390_/Y vdd gnd INVX1
X_9459_ _9459_/A _9459_/B _9459_/Y vdd gnd NAND2X1
X_10341_ _10341_/A _10341_/B _10341_/Y vdd gnd AND2X2
XFILL_1__9644_ vdd gnd FILL
X_13060_ _13060_/A _13060_/B _13060_/C _13060_/Y vdd gnd NAND3X1
X_10272_ _10272_/A _10272_/B _10272_/C _10272_/Y vdd gnd NAND3X1
XFILL_1__9575_ vdd gnd FILL
X_12011_ _12011_/A _12011_/B _12011_/C _12011_/Y vdd gnd OAI21X1
XFILL_1__8526_ vdd gnd FILL
XFILL_2__7250_ vdd gnd FILL
XFILL_1__8457_ vdd gnd FILL
X_13962_ _13962_/A _13962_/B _13962_/Y vdd gnd NAND2X1
XFILL_1__7408_ vdd gnd FILL
XFILL_2__7181_ vdd gnd FILL
XFILL_1__8388_ vdd gnd FILL
X_12913_ _12913_/A _12913_/Y vdd gnd INVX1
X_13893_ _13893_/A _13893_/B _13893_/C _13893_/Y vdd gnd NAND3X1
XFILL_1__7339_ vdd gnd FILL
X_12844_ _12844_/A _12844_/B _12844_/C _12844_/Y vdd gnd OAI21X1
XFILL_0__10580_ vdd gnd FILL
XFILL_1__9009_ vdd gnd FILL
X_12775_ _12775_/A _12775_/B _12775_/Y vdd gnd NAND2X1
XFILL_1__11870_ vdd gnd FILL
X_14514_ _14514_/D _14514_/CLK _14514_/Q vdd gnd DFFPOSX1
X_11726_ _11726_/A _11726_/B _11726_/C _11726_/Y vdd gnd OAI21X1
XFILL_1__10821_ vdd gnd FILL
XFILL_0__12250_ vdd gnd FILL
X_14445_ _14445_/A _14445_/B _14445_/Y vdd gnd NOR2X1
XFILL_2__10022_ vdd gnd FILL
X_11657_ _11657_/D _11657_/CLK _11657_/Q vdd gnd DFFPOSX1
XFILL_2__9753_ vdd gnd FILL
XFILL_1__13540_ vdd gnd FILL
XFILL_0__11201_ vdd gnd FILL
XFILL_0__12181_ vdd gnd FILL
X_10608_ _10608_/A _10608_/B _10608_/C _10608_/Y vdd gnd OAI21X1
X_14376_ _14376_/A _14376_/B _14376_/C _14376_/Y vdd gnd OAI21X1
X_11588_ _11588_/A _11588_/B _11588_/Y vdd gnd NAND2X1
XFILL_2__9684_ vdd gnd FILL
XFILL_0__11132_ vdd gnd FILL
XFILL_1__10683_ vdd gnd FILL
X_13327_ _13327_/A _13327_/B _13327_/Y vdd gnd OR2X2
X_10539_ _10539_/A _10539_/B _10539_/C _10539_/Y vdd gnd OAI21X1
XFILL_1__12422_ vdd gnd FILL
XFILL_0__11063_ vdd gnd FILL
XFILL_0__7650_ vdd gnd FILL
X_13258_ _13258_/A _13258_/B _13258_/Y vdd gnd NOR2X1
XFILL_2__10924_ vdd gnd FILL
XFILL_0__10014_ vdd gnd FILL
XFILL_1__12353_ vdd gnd FILL
X_12209_ _12209_/A _12209_/B _12209_/Y vdd gnd NOR2X1
XFILL_0__7581_ vdd gnd FILL
X_13189_ _13189_/A _13189_/B _13189_/C _13189_/Y vdd gnd OAI21X1
XFILL_2__7517_ vdd gnd FILL
XFILL_1__11304_ vdd gnd FILL
XFILL_0__14822_ vdd gnd FILL
XFILL_1__12284_ vdd gnd FILL
XFILL_2__10855_ vdd gnd FILL
XFILL_0__9320_ vdd gnd FILL
XFILL_1__14023_ vdd gnd FILL
XFILL_2__7448_ vdd gnd FILL
XFILL_1__11235_ vdd gnd FILL
XFILL_0__14753_ vdd gnd FILL
XFILL_2__10786_ vdd gnd FILL
XFILL_0__11965_ vdd gnd FILL
XFILL_0__9251_ vdd gnd FILL
XFILL_2__12525_ vdd gnd FILL
XFILL_0__13704_ vdd gnd FILL
XFILL_1__11166_ vdd gnd FILL
XFILL_2__7379_ vdd gnd FILL
XFILL_0__10916_ vdd gnd FILL
XFILL_0__14684_ vdd gnd FILL
XFILL_0__8202_ vdd gnd FILL
XFILL_0__11896_ vdd gnd FILL
XFILL_0__9182_ vdd gnd FILL
X_8830_ _8830_/A _8830_/B _8830_/Y vdd gnd NAND2X1
XFILL_1__10117_ vdd gnd FILL
XFILL_0__13635_ vdd gnd FILL
XBUFX2_insert2 BUFX2_insert2/A BUFX2_insert2/Y vdd gnd BUFX2
XFILL_2__12456_ vdd gnd FILL
XFILL_0__10847_ vdd gnd FILL
XFILL_1__11097_ vdd gnd FILL
XFILL_0__8133_ vdd gnd FILL
X_8761_ _8761_/A _8761_/B _8761_/Y vdd gnd NAND2X1
XFILL_1__10048_ vdd gnd FILL
XFILL_2__12387_ vdd gnd FILL
XFILL_0__13566_ vdd gnd FILL
X_7712_ _7712_/A _7712_/B _7712_/S _7712_/Y vdd gnd MUX2X1
XFILL_0__8064_ vdd gnd FILL
XFILL_0__10778_ vdd gnd FILL
X_8692_ _8692_/A _8692_/B _8692_/C _8692_/Y vdd gnd OAI21X1
XFILL_0__12517_ vdd gnd FILL
XFILL_1__14856_ vdd gnd FILL
X_7643_ _7643_/A _7643_/Y vdd gnd INVX1
XFILL_1__13807_ vdd gnd FILL
XFILL_0__12448_ vdd gnd FILL
XFILL_1__14787_ vdd gnd FILL
XFILL_1__11999_ vdd gnd FILL
X_7574_ _7574_/A _7574_/B _7574_/C _7574_/Y vdd gnd AOI21X1
XFILL_1__13738_ vdd gnd FILL
X_9313_ _9313_/A _9313_/B _9313_/Y vdd gnd NAND2X1
XFILL_0__12379_ vdd gnd FILL
XFILL_0__8966_ vdd gnd FILL
XFILL_0__14118_ vdd gnd FILL
XFILL_1__13669_ vdd gnd FILL
X_9244_ _9244_/A _9244_/Y vdd gnd INVX1
XFILL_1__7690_ vdd gnd FILL
XFILL_0__14049_ vdd gnd FILL
XFILL_0__7848_ vdd gnd FILL
X_9175_ _9175_/A _9175_/B _9175_/C _9175_/Y vdd gnd AOI21X1
X_8126_ _8126_/A _8126_/B _8126_/C _8126_/Y vdd gnd AOI21X1
XFILL_1__9360_ vdd gnd FILL
XFILL_0__7779_ vdd gnd FILL
XFILL_0__9518_ vdd gnd FILL
XFILL_1__8311_ vdd gnd FILL
X_8057_ _8057_/A _8057_/Y vdd gnd INVX8
XFILL_1__9291_ vdd gnd FILL
XFILL_0__9449_ vdd gnd FILL
XFILL_1__8242_ vdd gnd FILL
XFILL_1__8173_ vdd gnd FILL
XFILL_1__7124_ vdd gnd FILL
X_10890_ _10890_/A _10890_/B _10890_/S _10890_/Y vdd gnd MUX2X1
X_8959_ _8959_/A _8959_/B _8959_/C _8959_/Y vdd gnd OAI21X1
XFILL_1_CLKBUF1_insert40 vdd gnd FILL
X_12560_ _12560_/D _12560_/CLK _12560_/Q vdd gnd DFFPOSX1
XFILL_1_CLKBUF1_insert51 vdd gnd FILL
XFILL_1_CLKBUF1_insert62 vdd gnd FILL
XFILL_1_CLKBUF1_insert73 vdd gnd FILL
XFILL_1_CLKBUF1_insert84 vdd gnd FILL
X_11511_ _11511_/A _11511_/B _11511_/C _11511_/Y vdd gnd OAI21X1
XFILL_1_CLKBUF1_insert95 vdd gnd FILL
X_12491_ _12491_/A _12491_/Y vdd gnd INVX1
X_14230_ _14230_/A _14230_/B _14230_/C _14230_/Y vdd gnd OAI21X1
X_11442_ _11442_/A _11442_/B _11442_/C _11442_/Y vdd gnd OAI21X1
X_14161_ _14161_/D _14161_/CLK _14161_/Q vdd gnd DFFPOSX1
X_11373_ _11373_/A _11373_/B _11373_/C _11373_/Y vdd gnd AOI21X1
XFILL_1__7888_ vdd gnd FILL
X_13112_ _13112_/A _13112_/B _13112_/Y vdd gnd NAND2X1
X_10324_ _10324_/A _10324_/B _10324_/C _10324_/Y vdd gnd OAI21X1
XFILL_1__9627_ vdd gnd FILL
XFILL_2__8420_ vdd gnd FILL
X_14092_ _14092_/A _14092_/B _14092_/Y vdd gnd NAND2X1
X_10255_ _10255_/A _10255_/B _10255_/C _10255_/Y vdd gnd AOI21X1
X_13043_ _13043_/A _13043_/B _13043_/C _13043_/Y vdd gnd OAI21X1
XFILL_1__9558_ vdd gnd FILL
XFILL257550x79350 vdd gnd FILL
X_10186_ _10186_/A _10186_/B _10186_/C _10186_/Y vdd gnd OAI21X1
XFILL_1__8509_ vdd gnd FILL
XFILL_1__9489_ vdd gnd FILL
XFILL_1__11020_ vdd gnd FILL
XFILL_0__11750_ vdd gnd FILL
X_13945_ _13945_/A _13945_/B _13945_/C _13945_/Y vdd gnd OAI21X1
XFILL_2__12310_ vdd gnd FILL
X_13876_ _13876_/A _13876_/B _13876_/C _13876_/Y vdd gnd OAI21X1
XFILL_2__12241_ vdd gnd FILL
XFILL_0__13420_ vdd gnd FILL
XFILL_0__10632_ vdd gnd FILL
XFILL_1__12971_ vdd gnd FILL
X_12827_ _12827_/A _12827_/B _12827_/C _12827_/Y vdd gnd OAI21X1
XFILL_1__14710_ vdd gnd FILL
XFILL_2__12172_ vdd gnd FILL
XFILL_1__11922_ vdd gnd FILL
XFILL_0__13351_ vdd gnd FILL
XFILL_0__10563_ vdd gnd FILL
X_12758_ _12758_/A _12758_/B _12758_/C _12758_/Y vdd gnd NAND3X1
XFILL_0__12302_ vdd gnd FILL
XFILL_1__14641_ vdd gnd FILL
XFILL_1__11853_ vdd gnd FILL
XFILL_0__13282_ vdd gnd FILL
XFILL_0__10494_ vdd gnd FILL
X_11709_ _11709_/A _11709_/B _11709_/C _11709_/Y vdd gnd AOI21X1
X_12689_ _12689_/A _12689_/B _12689_/Y vdd gnd NAND2X1
XFILL_1__10804_ vdd gnd FILL
XFILL_0__12233_ vdd gnd FILL
XFILL_1__14572_ vdd gnd FILL
XFILL_1__11784_ vdd gnd FILL
XFILL_0__8820_ vdd gnd FILL
X_14428_ _14428_/A _14428_/B _14428_/C _14428_/Y vdd gnd OAI21X1
XFILL_2__10005_ vdd gnd FILL
XFILL_2__9736_ vdd gnd FILL
XFILL_1__13523_ vdd gnd FILL
XFILL_0__12164_ vdd gnd FILL
XFILL_0__8751_ vdd gnd FILL
X_14359_ _14359_/A _14359_/B _14359_/Y vdd gnd NOR2X1
XFILL_2__14813_ vdd gnd FILL
X_7290_ _7290_/A _7290_/B _7290_/C _7290_/Y vdd gnd OAI21X1
XFILL_2__9667_ vdd gnd FILL
XFILL_0__11115_ vdd gnd FILL
XFILL_1__10666_ vdd gnd FILL
XFILL_0__7702_ vdd gnd FILL
XFILL_0__12095_ vdd gnd FILL
XFILL_0__8682_ vdd gnd FILL
XFILL_1__12405_ vdd gnd FILL
XFILL_2__9598_ vdd gnd FILL
XFILL_1__13385_ vdd gnd FILL
XFILL_0__11046_ vdd gnd FILL
XFILL_1__10597_ vdd gnd FILL
XFILL_0__7633_ vdd gnd FILL
XFILL_1__12336_ vdd gnd FILL
XFILL_0__7564_ vdd gnd FILL
XFILL_0__14805_ vdd gnd FILL
XFILL_1__12267_ vdd gnd FILL
XFILL_0__9303_ vdd gnd FILL
XFILL_0__12997_ vdd gnd FILL
X_9931_ _9931_/A _9931_/B _9931_/Y vdd gnd NOR2X1
XFILL_1__14006_ vdd gnd FILL
XFILL_0__7495_ vdd gnd FILL
XFILL_1__11218_ vdd gnd FILL
XFILL_0__14736_ vdd gnd FILL
XFILL_0__11948_ vdd gnd FILL
XFILL_1__12198_ vdd gnd FILL
XFILL_2__10769_ vdd gnd FILL
XFILL_0__9234_ vdd gnd FILL
X_9862_ _9862_/A _9862_/Y vdd gnd INVX1
XFILL_2__12508_ vdd gnd FILL
XFILL_1__11149_ vdd gnd FILL
XFILL_0__14667_ vdd gnd FILL
XFILL_0__11879_ vdd gnd FILL
XFILL_0__9165_ vdd gnd FILL
X_8813_ _8813_/A _8813_/B _8813_/C _8813_/Y vdd gnd OAI21X1
X_9793_ _9793_/D _9793_/CLK _9793_/Q vdd gnd DFFPOSX1
XFILL_2__12439_ vdd gnd FILL
XFILL_0__13618_ vdd gnd FILL
XFILL_0__14598_ vdd gnd FILL
XFILL_0__8116_ vdd gnd FILL
XFILL_0__9096_ vdd gnd FILL
X_8744_ _8744_/A _8744_/Y vdd gnd INVX1
XFILL_1__14908_ vdd gnd FILL
XFILL_0__13549_ vdd gnd FILL
XFILL_0__8047_ vdd gnd FILL
X_8675_ _8675_/A _8675_/B _8675_/C _8675_/Y vdd gnd OAI21X1
XFILL_2__14109_ vdd gnd FILL
XFILL_1__14839_ vdd gnd FILL
X_7626_ _7626_/A _7626_/Y vdd gnd INVX1
XFILL_1__7811_ vdd gnd FILL
X_7557_ _7557_/A _7557_/B _7557_/C _7557_/Y vdd gnd OAI21X1
XFILL_1_CLKBUF1_insert106 vdd gnd FILL
XFILL_0__9998_ vdd gnd FILL
XFILL_1__8791_ vdd gnd FILL
XFILL_0__8949_ vdd gnd FILL
XFILL_1__7742_ vdd gnd FILL
X_7488_ _7488_/A _7488_/B _7488_/Y vdd gnd NAND2X1
X_9227_ _9227_/A _9227_/B _9227_/C _9227_/Y vdd gnd NOR3X1
XFILL_1__7673_ vdd gnd FILL
XFILL_1__9412_ vdd gnd FILL
X_9158_ _9158_/A _9158_/B _9158_/C _9158_/Y vdd gnd NAND3X1
X_10040_ _10040_/A _10040_/B _10040_/Y vdd gnd OR2X2
X_8109_ _8109_/A _8109_/B _8109_/S _8109_/Y vdd gnd MUX2X1
XFILL_1__9343_ vdd gnd FILL
X_9089_ _9089_/A _9089_/B _9089_/C _9089_/Y vdd gnd OAI21X1
XFILL_1__9274_ vdd gnd FILL
XFILL_1__8225_ vdd gnd FILL
X_11991_ _11991_/A _11991_/B _11991_/Y vdd gnd NAND2X1
X_13730_ _13730_/A _13730_/B _13730_/C _13730_/Y vdd gnd OAI21X1
X_10942_ _10942_/A _10942_/B _10942_/C _10942_/Y vdd gnd NAND3X1
XFILL_1__8156_ vdd gnd FILL
X_13661_ _13661_/A _13661_/Y vdd gnd INVX1
XFILL_1__7107_ vdd gnd FILL
X_10873_ _10873_/A _10873_/B _10873_/C _10873_/Y vdd gnd OAI21X1
XFILL_1__8087_ vdd gnd FILL
X_12612_ _12612_/D _12612_/CLK _12612_/Q vdd gnd DFFPOSX1
X_13592_ _13592_/A _13592_/B _13592_/S _13592_/Y vdd gnd MUX2X1
XFILL257550x54150 vdd gnd FILL
X_12543_ _12543_/D _12543_/CLK _12543_/Q vdd gnd DFFPOSX1
XFILL_2__7851_ vdd gnd FILL
X_12474_ _12474_/A _12474_/B _12474_/Y vdd gnd NAND2X1
XFILL_1__8989_ vdd gnd FILL
XFILL_2__7782_ vdd gnd FILL
X_14213_ _14213_/D _14213_/CLK _14213_/Q vdd gnd DFFPOSX1
X_11425_ _11425_/A _11425_/B _11425_/Y vdd gnd NOR2X1
XFILL_1__10520_ vdd gnd FILL
X_14144_ _14144_/A _14144_/B _14144_/C _14144_/Y vdd gnd OAI21X1
X_11356_ _11356_/A _11356_/B _11356_/C _11356_/Y vdd gnd OAI21X1
XFILL_2__11810_ vdd gnd FILL
XFILL_1__10451_ vdd gnd FILL
X_10307_ _10307_/A _10307_/B _10307_/C _10307_/Y vdd gnd OAI21X1
XCLKBUF1_insert105 CLKBUF1_insert105/A CLKBUF1_insert105/Y vdd gnd CLKBUF1
XFILL_2__8403_ vdd gnd FILL
X_14075_ _14075_/A _14075_/Y vdd gnd INVX1
X_11287_ _11287_/A _11287_/B _11287_/Y vdd gnd AND2X2
XFILL_1__13170_ vdd gnd FILL
XFILL_2__11741_ vdd gnd FILL
XFILL_0__12920_ vdd gnd FILL
XFILL_1__10382_ vdd gnd FILL
X_13026_ _13026_/A _13026_/B _13026_/C _13026_/Y vdd gnd OAI21X1
X_10238_ _10238_/A _10238_/B _10238_/C _10238_/Y vdd gnd OAI21X1
XFILL_2__8334_ vdd gnd FILL
XFILL_1__12121_ vdd gnd FILL
XFILL_0__12851_ vdd gnd FILL
X_10169_ _10169_/A _10169_/B _10169_/C _10169_/Y vdd gnd AOI21X1
XFILL_2__10623_ vdd gnd FILL
XFILL_1__12052_ vdd gnd FILL
XFILL_0__11802_ vdd gnd FILL
XFILL_2__8265_ vdd gnd FILL
XFILL_0__12782_ vdd gnd FILL
XFILL_0__7280_ vdd gnd FILL
XFILL_1__11003_ vdd gnd FILL
XFILL_2__10554_ vdd gnd FILL
XFILL_0__11733_ vdd gnd FILL
XFILL_2__8196_ vdd gnd FILL
X_13928_ _13928_/A _13928_/B _13928_/Y vdd gnd NAND2X1
XFILL_0__14452_ vdd gnd FILL
X_13859_ _13859_/A _13859_/B _13859_/Y vdd gnd NAND2X1
XFILL_2__12224_ vdd gnd FILL
XFILL_0__13403_ vdd gnd FILL
XFILL_0__10615_ vdd gnd FILL
XFILL_1__12954_ vdd gnd FILL
XFILL_0__14383_ vdd gnd FILL
XFILL_1_BUFX2_insert260 vdd gnd FILL
XFILL_0__11595_ vdd gnd FILL
XFILL_1_BUFX2_insert271 vdd gnd FILL
XCLKBUF1_insert31 CLKBUF1_insert31/A CLKBUF1_insert31/Y vdd gnd CLKBUF1
XFILL_1__11905_ vdd gnd FILL
XFILL_2__12155_ vdd gnd FILL
XCLKBUF1_insert42 CLKBUF1_insert42/A CLKBUF1_insert42/Y vdd gnd CLKBUF1
XFILL_0__13334_ vdd gnd FILL
XFILL_1_BUFX2_insert282 vdd gnd FILL
XFILL_0__10546_ vdd gnd FILL
XFILL_1_BUFX2_insert293 vdd gnd FILL
XFILL_1__12885_ vdd gnd FILL
XFILL_0__9921_ vdd gnd FILL
XCLKBUF1_insert53 CLKBUF1_insert53/A CLKBUF1_insert53/Y vdd gnd CLKBUF1
XCLKBUF1_insert64 CLKBUF1_insert64/A CLKBUF1_insert64/Y vdd gnd CLKBUF1
X_8460_ _8460_/A _8460_/Y vdd gnd INVX1
XCLKBUF1_insert75 CLKBUF1_insert75/A CLKBUF1_insert75/Y vdd gnd CLKBUF1
XCLKBUF1_insert86 CLKBUF1_insert86/A CLKBUF1_insert86/Y vdd gnd CLKBUF1
XFILL_1__14624_ vdd gnd FILL
XFILL_2__12086_ vdd gnd FILL
XFILL_1__11836_ vdd gnd FILL
XFILL_0__13265_ vdd gnd FILL
XCLKBUF1_insert97 CLKBUF1_insert97/A CLKBUF1_insert97/Y vdd gnd CLKBUF1
X_7411_ _7411_/A _7411_/B _7411_/C _7411_/Y vdd gnd AOI21X1
XFILL_0__10477_ vdd gnd FILL
XFILL_0__9852_ vdd gnd FILL
X_8391_ _8391_/A _8391_/Y vdd gnd INVX1
XFILL_0__12216_ vdd gnd FILL
XFILL_0__13196_ vdd gnd FILL
XFILL_1__11767_ vdd gnd FILL
XFILL_0__8803_ vdd gnd FILL
X_7342_ _7342_/A _7342_/B _7342_/Y vdd gnd NAND2X1
XFILL_1__13506_ vdd gnd FILL
XFILL_0__12147_ vdd gnd FILL
XFILL_1__14486_ vdd gnd FILL
XFILL_1__11698_ vdd gnd FILL
XFILL_0__8734_ vdd gnd FILL
X_7273_ _7273_/A _7273_/B _7273_/Y vdd gnd AND2X2
XFILL_1__10649_ vdd gnd FILL
X_9012_ _9012_/A _9012_/B _9012_/Y vdd gnd NAND2X1
XFILL_0__12078_ vdd gnd FILL
XFILL_2__12988_ vdd gnd FILL
XFILL_0__8665_ vdd gnd FILL
XFILL_2__14727_ vdd gnd FILL
XFILL_0__11029_ vdd gnd FILL
XFILL_1__13368_ vdd gnd FILL
XFILL_0__7616_ vdd gnd FILL
XFILL_0__8596_ vdd gnd FILL
XFILL_2__14658_ vdd gnd FILL
XFILL_1__12319_ vdd gnd FILL
XFILL_1__13299_ vdd gnd FILL
XFILL_0__7547_ vdd gnd FILL
XFILL_2__14589_ vdd gnd FILL
X_9914_ _9914_/A _9914_/B _9914_/Y vdd gnd NAND2X1
XFILL_0__7478_ vdd gnd FILL
XFILL_0__14719_ vdd gnd FILL
XFILL_0__9217_ vdd gnd FILL
XFILL_1__8010_ vdd gnd FILL
X_9845_ _9845_/A _9845_/Y vdd gnd INVX2
XFILL_0__9148_ vdd gnd FILL
X_9776_ _9776_/D _9776_/CLK _9776_/Q vdd gnd DFFPOSX1
XFILL_0__9079_ vdd gnd FILL
XFILL_1__9961_ vdd gnd FILL
X_8727_ _8727_/A _8727_/B _8727_/C _8727_/Y vdd gnd AOI21X1
XFILL_1__9892_ vdd gnd FILL
X_8658_ _8658_/A _8658_/B _8658_/C _8658_/Y vdd gnd AOI21X1
X_7609_ _7609_/A _7609_/B _7609_/C _7609_/Y vdd gnd NAND3X1
X_8589_ _8589_/A _8589_/B _8589_/Y vdd gnd OR2X2
XFILL_1__8774_ vdd gnd FILL
X_11210_ _11210_/A _11210_/B _11210_/Y vdd gnd NAND2X1
X_12190_ _12190_/A _12190_/B _12190_/C _12190_/Y vdd gnd OAI21X1
XFILL_1__7725_ vdd gnd FILL
X_11141_ _11141_/A _11141_/B _11141_/Y vdd gnd NAND2X1
XFILL_1__7656_ vdd gnd FILL
X_11072_ _11072_/A _11072_/Y vdd gnd INVX1
XFILL_1__7587_ vdd gnd FILL
X_14900_ _14900_/D _14900_/CLK _14900_/Q vdd gnd DFFPOSX1
X_10023_ _10023_/A _10023_/B _10023_/C _10023_/Y vdd gnd AOI21X1
XFILL_1__9326_ vdd gnd FILL
X_14831_ _14831_/A _14831_/B _14831_/C _14831_/Y vdd gnd AOI21X1
XFILL_1__9257_ vdd gnd FILL
XFILL_2__8050_ vdd gnd FILL
X_14762_ _14762_/A _14762_/B _14762_/Y vdd gnd AND2X2
XFILL_1__8208_ vdd gnd FILL
X_11974_ _11974_/A _11974_/B _11974_/C _11974_/Y vdd gnd AOI21X1
XFILL_1__9188_ vdd gnd FILL
X_13713_ _13713_/A _13713_/Y vdd gnd INVX1
X_10925_ _10925_/A _10925_/B _10925_/C _10925_/Y vdd gnd OAI21X1
X_14693_ _14693_/A _14693_/B _14693_/Y vdd gnd OR2X2
XFILL_1__8139_ vdd gnd FILL
XFILL_2__10270_ vdd gnd FILL
X_13644_ _13644_/A _13644_/B _13644_/C _13644_/Y vdd gnd OAI21X1
X_10856_ _10856_/A _10856_/B _10856_/S _10856_/Y vdd gnd MUX2X1
XFILL_0__10400_ vdd gnd FILL
XFILL_2__8952_ vdd gnd FILL
XFILL_0_BUFX2_insert201 vdd gnd FILL
XFILL_0__11380_ vdd gnd FILL
XFILL_0_BUFX2_insert212 vdd gnd FILL
XFILL_2__7903_ vdd gnd FILL
XFILL_0_BUFX2_insert223 vdd gnd FILL
X_13575_ _13575_/A _13575_/B _13575_/S _13575_/Y vdd gnd MUX2X1
X_10787_ _10787_/A _10787_/B _10787_/Y vdd gnd NAND2X1
XFILL_0__10331_ vdd gnd FILL
XFILL_0_BUFX2_insert234 vdd gnd FILL
XFILL_0_BUFX2_insert245 vdd gnd FILL
XFILL_1__12670_ vdd gnd FILL
XFILL_0_BUFX2_insert256 vdd gnd FILL
X_12526_ _12526_/A _12526_/B _12526_/Y vdd gnd NAND2X1
XFILL_0_BUFX2_insert267 vdd gnd FILL
XFILL_2__7834_ vdd gnd FILL
XFILL_0_BUFX2_insert278 vdd gnd FILL
XFILL_0__13050_ vdd gnd FILL
XFILL_0__10262_ vdd gnd FILL
XFILL_0_BUFX2_insert289 vdd gnd FILL
X_12457_ _12457_/A _12457_/B _12457_/Y vdd gnd NAND2X1
XFILL_0__12001_ vdd gnd FILL
XFILL_2__7765_ vdd gnd FILL
XFILL_1__14340_ vdd gnd FILL
XFILL_1__11552_ vdd gnd FILL
XFILL_0__10193_ vdd gnd FILL
X_11408_ _11408_/A _11408_/B _11408_/S _11408_/Y vdd gnd MUX2X1
XFILL_1__10503_ vdd gnd FILL
X_12388_ _12388_/A _12388_/B _12388_/C _12388_/Y vdd gnd OAI21X1
XFILL_2__7696_ vdd gnd FILL
XFILL_1__14271_ vdd gnd FILL
XFILL_1__11483_ vdd gnd FILL
XFILL_2_BUFX2_insert27 vdd gnd FILL
X_14127_ _14127_/A _14127_/B _14127_/Y vdd gnd NAND2X1
X_11339_ _11339_/A _11339_/Y vdd gnd INVX1
XFILL_1__10434_ vdd gnd FILL
XFILL_1__13222_ vdd gnd FILL
XFILL_0__13952_ vdd gnd FILL
XFILL_0__8450_ vdd gnd FILL
X_14058_ _14058_/A _14058_/B _14058_/C _14058_/Y vdd gnd OAI21X1
XFILL_1__13153_ vdd gnd FILL
XFILL_2__11724_ vdd gnd FILL
XFILL_0__12903_ vdd gnd FILL
XFILL_1__10365_ vdd gnd FILL
XFILL_0__7401_ vdd gnd FILL
X_13009_ _13009_/A _13009_/B _13009_/C _13009_/Y vdd gnd OAI21X1
XFILL_0__13883_ vdd gnd FILL
XFILL_2__8317_ vdd gnd FILL
XFILL_0__8381_ vdd gnd FILL
XFILL_1__12104_ vdd gnd FILL
XFILL_1__13084_ vdd gnd FILL
XFILL_1__10296_ vdd gnd FILL
XFILL_0__12834_ vdd gnd FILL
XFILL_0__7332_ vdd gnd FILL
X_7960_ _7960_/D _7960_/CLK _7960_/Q vdd gnd DFFPOSX1
XFILL_2__10606_ vdd gnd FILL
XFILL_1__12035_ vdd gnd FILL
XFILL_2__8248_ vdd gnd FILL
XFILL_0__12765_ vdd gnd FILL
XFILL_0__7263_ vdd gnd FILL
X_7891_ _7891_/A _7891_/B _7891_/C _7891_/Y vdd gnd OAI21X1
XFILL_2__10537_ vdd gnd FILL
XFILL_0__11716_ vdd gnd FILL
XFILL_2__8179_ vdd gnd FILL
XFILL_0__9002_ vdd gnd FILL
XFILL_0__12696_ vdd gnd FILL
XFILL_0__7194_ vdd gnd FILL
X_9630_ _9630_/A _9630_/B _9630_/Y vdd gnd NAND2X1
XFILL_2__10468_ vdd gnd FILL
XFILL_0__14435_ vdd gnd FILL
XFILL_1__13986_ vdd gnd FILL
X_9561_ _9561_/A _9561_/B _9561_/Y vdd gnd NAND2X1
XFILL_1__12937_ vdd gnd FILL
XFILL_2__10399_ vdd gnd FILL
XFILL_0__14366_ vdd gnd FILL
XFILL_0__11578_ vdd gnd FILL
X_8512_ _8512_/A _8512_/B _8512_/Y vdd gnd NAND2X1
X_9492_ _9492_/A _9492_/B _9492_/C _9492_/Y vdd gnd OAI21X1
XFILL_0__13317_ vdd gnd FILL
XFILL_0__10529_ vdd gnd FILL
XFILL_0__9904_ vdd gnd FILL
XFILL_0__14297_ vdd gnd FILL
XFILL_1__12868_ vdd gnd FILL
X_8443_ _8443_/A _8443_/B _8443_/Y vdd gnd OR2X2
XFILL_1__14607_ vdd gnd FILL
XFILL_1__11819_ vdd gnd FILL
XFILL_0__13248_ vdd gnd FILL
XFILL_1__12799_ vdd gnd FILL
X_8374_ _8374_/A _8374_/B _8374_/Y vdd gnd NOR2X1
XFILL_0__13179_ vdd gnd FILL
X_7325_ _7325_/A _7325_/B _7325_/C _7325_/Y vdd gnd AOI21X1
XFILL_1__14469_ vdd gnd FILL
XFILL_1__7510_ vdd gnd FILL
XFILL_0__8717_ vdd gnd FILL
X_7256_ _7256_/A _7256_/B _7256_/C _7256_/D _7256_/Y vdd gnd AOI22X1
XFILL_0__9697_ vdd gnd FILL
XFILL_1__8490_ vdd gnd FILL
XFILL_1__7441_ vdd gnd FILL
XFILL_0__8648_ vdd gnd FILL
X_7187_ _7187_/A _7187_/B _7187_/C _7187_/Y vdd gnd NAND3X1
XFILL_1__7372_ vdd gnd FILL
XFILL_0__8579_ vdd gnd FILL
XFILL_1_BUFX2_insert2 vdd gnd FILL
XFILL_1__9111_ vdd gnd FILL
XFILL_2_BUFX2_insert318 vdd gnd FILL
XFILL_1__9042_ vdd gnd FILL
X_9828_ _9828_/D _9828_/CLK _9828_/Q vdd gnd DFFPOSX1
X_10710_ _10710_/D _10710_/CLK _10710_/Q vdd gnd DFFPOSX1
X_11690_ _11690_/D _11690_/CLK _11690_/Q vdd gnd DFFPOSX1
X_9759_ _9759_/A _9759_/B _9759_/C _9759_/Y vdd gnd OAI21X1
XBUFX2_insert306 BUFX2_insert306/A BUFX2_insert306/Y vdd gnd BUFX2
XBUFX2_insert317 BUFX2_insert317/A BUFX2_insert317/Y vdd gnd BUFX2
X_10641_ _10641_/A _10641_/B _10641_/C _10641_/Y vdd gnd OAI21X1
XFILL_1__9944_ vdd gnd FILL
XBUFX2_insert328 BUFX2_insert328/A BUFX2_insert328/Y vdd gnd BUFX2
XBUFX2_insert339 BUFX2_insert339/A BUFX2_insert339/Y vdd gnd BUFX2
X_13360_ _13360_/A _13360_/B _13360_/C _13360_/Y vdd gnd OAI21X1
X_10572_ _10572_/A _10572_/B _10572_/Y vdd gnd NOR2X1
XFILL_1__9875_ vdd gnd FILL
X_12311_ _12311_/A _12311_/B _12311_/Y vdd gnd NAND2X1
XFILL_1__8826_ vdd gnd FILL
X_13291_ _13291_/A _13291_/B _13291_/C _13291_/Y vdd gnd OAI21X1
X_12242_ _12242_/A _12242_/Y vdd gnd INVX1
XFILL_1__8757_ vdd gnd FILL
XFILL_1__7708_ vdd gnd FILL
X_12173_ _12173_/A _12173_/B _12173_/Y vdd gnd NAND2X1
XFILL_1__8688_ vdd gnd FILL
X_11124_ _11124_/A _11124_/Y vdd gnd INVX1
XFILL_1__7639_ vdd gnd FILL
X_11055_ _11055_/A _11055_/B _11055_/Y vdd gnd NOR2X1
XFILL_1__10150_ vdd gnd FILL
X_10006_ _10006_/A _10006_/Y vdd gnd INVX1
XFILL_0__10880_ vdd gnd FILL
XFILL_1__9309_ vdd gnd FILL
XFILL_1__10081_ vdd gnd FILL
X_14814_ _14814_/A _14814_/B _14814_/C _14814_/Y vdd gnd AOI21X1
XFILL_2__8033_ vdd gnd FILL
X_14745_ _14745_/A _14745_/B _14745_/Y vdd gnd NOR2X1
XFILL_2__13110_ vdd gnd FILL
X_11957_ _11957_/A _11957_/B _11957_/Y vdd gnd NAND2X1
XFILL_2__10322_ vdd gnd FILL
XFILL_0__11501_ vdd gnd FILL
XFILL_2__14090_ vdd gnd FILL
XFILL_1__13840_ vdd gnd FILL
XFILL_0__12481_ vdd gnd FILL
X_10908_ _10908_/A _10908_/B _10908_/Y vdd gnd NAND2X1
X_14676_ _14676_/A _14676_/B _14676_/Y vdd gnd OR2X2
XFILL_2__10253_ vdd gnd FILL
X_11888_ _11888_/A _11888_/B _11888_/Y vdd gnd OR2X2
XFILL_0__14220_ vdd gnd FILL
XFILL_2__13041_ vdd gnd FILL
XFILL_0__11432_ vdd gnd FILL
XFILL_1__13771_ vdd gnd FILL
XFILL_1__10983_ vdd gnd FILL
X_13627_ _13627_/A _13627_/B _13627_/C _13627_/D _13627_/Y vdd gnd OAI22X1
X_10839_ _10839_/A _10839_/B _10839_/C _10839_/Y vdd gnd OAI21X1
XFILL_2__10184_ vdd gnd FILL
XFILL_0__14151_ vdd gnd FILL
XFILL_1__12722_ vdd gnd FILL
XFILL_0__11363_ vdd gnd FILL
X_13558_ _13558_/A _13558_/Y vdd gnd INVX1
XFILL_0__13102_ vdd gnd FILL
XFILL_0__10314_ vdd gnd FILL
XFILL_1__12653_ vdd gnd FILL
XFILL_0__14082_ vdd gnd FILL
X_12509_ _12509_/A _12509_/B _12509_/C _12509_/Y vdd gnd OAI21X1
XFILL_0__11294_ vdd gnd FILL
XFILL_0__7881_ vdd gnd FILL
X_13489_ _13489_/D _13489_/CLK _13489_/Q vdd gnd DFFPOSX1
XFILL_1__11604_ vdd gnd FILL
XFILL_0__13033_ vdd gnd FILL
XFILL_0__10245_ vdd gnd FILL
XFILL_0__9620_ vdd gnd FILL
XFILL_1__14323_ vdd gnd FILL
XFILL_1__11535_ vdd gnd FILL
XFILL_0__10176_ vdd gnd FILL
X_7110_ _7110_/A _7110_/B _7110_/C _7110_/Y vdd gnd OAI21X1
XFILL_0__9551_ vdd gnd FILL
X_8090_ _8090_/A _8090_/B _8090_/C _8090_/Y vdd gnd NAND3X1
XFILL_2__7679_ vdd gnd FILL
XFILL_1__14254_ vdd gnd FILL
XFILL_1__11466_ vdd gnd FILL
XFILL_0__8502_ vdd gnd FILL
XFILL_0__9482_ vdd gnd FILL
XFILL_1__13205_ vdd gnd FILL
XFILL_1__10417_ vdd gnd FILL
XFILL_0__13935_ vdd gnd FILL
XFILL_1__11397_ vdd gnd FILL
XFILL_0__8433_ vdd gnd FILL
XFILL_2__11707_ vdd gnd FILL
XFILL_1__13136_ vdd gnd FILL
XFILL_1__10348_ vdd gnd FILL
XFILL_0__13866_ vdd gnd FILL
XFILL_0__8364_ vdd gnd FILL
X_8992_ _8992_/A _8992_/Y vdd gnd INVX1
XFILL_1__10279_ vdd gnd FILL
XFILL_0__12817_ vdd gnd FILL
XFILL_1__13067_ vdd gnd FILL
XFILL_0__7315_ vdd gnd FILL
XFILL_0__13797_ vdd gnd FILL
X_7943_ _7943_/D _7943_/CLK _7943_/Q vdd gnd DFFPOSX1
XFILL_0__8295_ vdd gnd FILL
XFILL_1__12018_ vdd gnd FILL
XFILL_0__12748_ vdd gnd FILL
XFILL_0__7246_ vdd gnd FILL
XFILL_2__13308_ vdd gnd FILL
X_7874_ _7874_/A _7874_/B _7874_/Y vdd gnd NAND2X1
X_9613_ _9613_/A _9613_/B _9613_/C _9613_/Y vdd gnd OAI21X1
XFILL_0__12679_ vdd gnd FILL
XFILL_0__7177_ vdd gnd FILL
XFILL_2__13239_ vdd gnd FILL
XFILL_0__14418_ vdd gnd FILL
XFILL_1__13969_ vdd gnd FILL
X_9544_ _9544_/A _9544_/B _9544_/C _9544_/Y vdd gnd AOI21X1
XFILL_0__14349_ vdd gnd FILL
X_9475_ _9475_/A _9475_/B _9475_/C _9475_/Y vdd gnd NAND3X1
XFILL_1__9660_ vdd gnd FILL
X_8426_ _8426_/A _8426_/B _8426_/C _8426_/Y vdd gnd AOI21X1
XFILL_1__8611_ vdd gnd FILL
XFILL257250x100950 vdd gnd FILL
XFILL_1__9591_ vdd gnd FILL
X_8357_ _8357_/A _8357_/B _8357_/Y vdd gnd NAND2X1
X_7308_ _7308_/A _7308_/B _7308_/Y vdd gnd NAND2X1
XFILL_0__9749_ vdd gnd FILL
XFILL_1__8542_ vdd gnd FILL
X_8288_ _8288_/A _8288_/B _8288_/C _8288_/Y vdd gnd OAI21X1
X_7239_ _7239_/A _7239_/B _7239_/C _7239_/Y vdd gnd OAI21X1
XFILL_1__8473_ vdd gnd FILL
XFILL_1__7424_ vdd gnd FILL
XFILL_1__7355_ vdd gnd FILL
XFILL_2_BUFX2_insert115 vdd gnd FILL
XFILL_2_BUFX2_insert137 vdd gnd FILL
XFILL_2_BUFX2_insert148 vdd gnd FILL
X_12860_ _12860_/A _12860_/B _12860_/Y vdd gnd AND2X2
XFILL_1__7286_ vdd gnd FILL
X_11811_ _11811_/A _11811_/B _11811_/S _11811_/Y vdd gnd MUX2X1
XFILL_1__9025_ vdd gnd FILL
X_12791_ _12791_/A _12791_/B _12791_/C _12791_/Y vdd gnd AOI21X1
X_14530_ _14530_/D _14530_/CLK _14530_/Q vdd gnd DFFPOSX1
X_11742_ _11742_/A _11742_/B _11742_/Y vdd gnd NAND2X1
X_14461_ _14461_/A _14461_/B _14461_/Y vdd gnd NAND2X1
X_11673_ _11673_/D _11673_/CLK _11673_/Q vdd gnd DFFPOSX1
XFILL257550x180150 vdd gnd FILL
XBUFX2_insert114 BUFX2_insert114/A BUFX2_insert114/Y vdd gnd BUFX2
XBUFX2_insert125 BUFX2_insert125/A BUFX2_insert125/Y vdd gnd BUFX2
XBUFX2_insert136 BUFX2_insert136/A BUFX2_insert136/Y vdd gnd BUFX2
X_13412_ _13412_/A _13412_/B _13412_/Y vdd gnd NAND2X1
XBUFX2_insert147 BUFX2_insert147/A BUFX2_insert147/Y vdd gnd BUFX2
X_10624_ _10624_/A _10624_/B _10624_/Y vdd gnd NAND2X1
XFILL_2__8720_ vdd gnd FILL
X_14392_ _14392_/A _14392_/Y vdd gnd INVX1
XBUFX2_insert158 BUFX2_insert158/A BUFX2_insert158/Y vdd gnd BUFX2
XFILL_1__9927_ vdd gnd FILL
XBUFX2_insert169 BUFX2_insert169/A BUFX2_insert169/Y vdd gnd BUFX2
X_13343_ _13343_/A _13343_/B _13343_/C _13343_/Y vdd gnd OAI21X1
X_10555_ _10555_/A _10555_/Y vdd gnd INVX1
XFILL_1__9858_ vdd gnd FILL
XFILL_2__8651_ vdd gnd FILL
X_13274_ _13274_/A _13274_/Y vdd gnd INVX1
X_10486_ _10486_/A _10486_/B _10486_/Y vdd gnd OR2X2
XFILL_1__8809_ vdd gnd FILL
XFILL_0__10030_ vdd gnd FILL
XFILL_2__8582_ vdd gnd FILL
X_12225_ _12225_/A _12225_/B _12225_/C _12225_/Y vdd gnd NAND3X1
XFILL_1__11320_ vdd gnd FILL
X_12156_ _12156_/A _12156_/Y vdd gnd INVX1
XFILL_1__11251_ vdd gnd FILL
XFILL_0__11981_ vdd gnd FILL
X_11107_ _11107_/A _11107_/B _11107_/C _11107_/Y vdd gnd AOI21X1
XFILL_2__9203_ vdd gnd FILL
XFILL_1__10202_ vdd gnd FILL
X_12087_ _12087_/A _12087_/Y vdd gnd INVX1
XFILL_2_CLKBUF1_insert384 vdd gnd FILL
XFILL_0__10932_ vdd gnd FILL
XFILL_0__13720_ vdd gnd FILL
XFILL_1__11182_ vdd gnd FILL
X_11038_ _11038_/A _11038_/B _11038_/Y vdd gnd NAND2X1
XFILL_1__10133_ vdd gnd FILL
XFILL_2__12472_ vdd gnd FILL
XFILL_0__13651_ vdd gnd FILL
XFILL_0__10863_ vdd gnd FILL
XFILL_1__10064_ vdd gnd FILL
XFILL_0__7100_ vdd gnd FILL
XFILL_0__13582_ vdd gnd FILL
XFILL_0__10794_ vdd gnd FILL
XFILL_0__8080_ vdd gnd FILL
XFILL_2__14142_ vdd gnd FILL
X_12989_ _12989_/A _12989_/B _12989_/Y vdd gnd NAND2X1
XFILL_0__12533_ vdd gnd FILL
X_14728_ _14728_/A _14728_/B _14728_/Y vdd gnd NOR2X1
XFILL_2__14073_ vdd gnd FILL
XFILL_1__13823_ vdd gnd FILL
XFILL_0__12464_ vdd gnd FILL
X_14659_ _14659_/A _14659_/B _14659_/C _14659_/Y vdd gnd OAI21X1
XFILL_2__13024_ vdd gnd FILL
X_7590_ _7590_/A _7590_/B _7590_/Y vdd gnd AND2X2
XFILL_0__11415_ vdd gnd FILL
XFILL_1__13754_ vdd gnd FILL
XFILL_1__10966_ vdd gnd FILL
XFILL_0__12395_ vdd gnd FILL
XFILL_0__8982_ vdd gnd FILL
XFILL_1__12705_ vdd gnd FILL
XFILL_0__11346_ vdd gnd FILL
XFILL_0__14134_ vdd gnd FILL
XFILL_1__13685_ vdd gnd FILL
XFILL_1__10897_ vdd gnd FILL
X_9260_ _9260_/A _9260_/B _9260_/Y vdd gnd AND2X2
XFILL_2__10098_ vdd gnd FILL
XFILL_0__14065_ vdd gnd FILL
XFILL_1__12636_ vdd gnd FILL
XFILL_0__11277_ vdd gnd FILL
X_8211_ _8211_/A _8211_/B _8211_/C _8211_/Y vdd gnd NAND3X1
X_9191_ _9191_/A _9191_/Y vdd gnd INVX1
XFILL_0__7864_ vdd gnd FILL
XFILL_0__13016_ vdd gnd FILL
XFILL_0__10228_ vdd gnd FILL
XFILL_0__9603_ vdd gnd FILL
X_8142_ _8142_/A _8142_/B _8142_/C _8142_/Y vdd gnd OAI21X1
XFILL_0__7795_ vdd gnd FILL
XFILL_1__14306_ vdd gnd FILL
XFILL_1__11518_ vdd gnd FILL
XFILL_0__10159_ vdd gnd FILL
XFILL_0__9534_ vdd gnd FILL
XFILL_1__12498_ vdd gnd FILL
X_8073_ _8073_/A _8073_/B _8073_/Y vdd gnd NOR2X1
XFILL_1__14237_ vdd gnd FILL
XFILL_1__11449_ vdd gnd FILL
XFILL_0__9465_ vdd gnd FILL
XFILL_0__13918_ vdd gnd FILL
XFILL_0__8416_ vdd gnd FILL
XFILL_0__9396_ vdd gnd FILL
XFILL_1__13119_ vdd gnd FILL
XFILL_0__13849_ vdd gnd FILL
XFILL_1__14099_ vdd gnd FILL
XFILL_1__7140_ vdd gnd FILL
XFILL_0__8347_ vdd gnd FILL
XFILL_2__14409_ vdd gnd FILL
X_8975_ _8975_/A _8975_/B _8975_/C _8975_/Y vdd gnd OAI21X1
X_7926_ _7926_/D _7926_/CLK _7926_/Q vdd gnd DFFPOSX1
XFILL_0__8278_ vdd gnd FILL
XFILL_0__7229_ vdd gnd FILL
X_7857_ _7857_/A _7857_/B _7857_/C _7857_/Y vdd gnd OAI21X1
X_7788_ _7788_/A _7788_/Y vdd gnd INVX1
X_9527_ _9527_/A _9527_/B _9527_/Y vdd gnd NOR2X1
XFILL_1__9712_ vdd gnd FILL
X_9458_ _9458_/A _9458_/B _9458_/C _9458_/Y vdd gnd NAND3X1
X_10340_ _10340_/A _10340_/B _10340_/Y vdd gnd NOR2X1
XFILL_1__9643_ vdd gnd FILL
X_8409_ _8409_/A _8409_/B _8409_/Y vdd gnd NAND2X1
X_9389_ _9389_/A _9389_/B _9389_/C _9389_/Y vdd gnd OAI21X1
X_10271_ _10271_/A _10271_/B _10271_/C _10271_/Y vdd gnd OAI21X1
XFILL_1__9574_ vdd gnd FILL
X_12010_ _12010_/A _12010_/B _12010_/Y vdd gnd AND2X2
XFILL_1__8525_ vdd gnd FILL
XFILL_1__8456_ vdd gnd FILL
X_13961_ _13961_/A _13961_/B _13961_/Y vdd gnd OR2X2
XFILL_1__7407_ vdd gnd FILL
XFILL_1__8387_ vdd gnd FILL
X_12912_ _12912_/A _12912_/B _12912_/C _12912_/Y vdd gnd OAI21X1
X_13892_ _13892_/A _13892_/Y vdd gnd INVX1
XFILL_1__7338_ vdd gnd FILL
X_12843_ _12843_/A _12843_/Y vdd gnd INVX1
XFILL_1__7269_ vdd gnd FILL
XFILL_1__9008_ vdd gnd FILL
X_12774_ _12774_/A _12774_/Y vdd gnd INVX1
X_14513_ _14513_/D _14513_/CLK _14513_/Q vdd gnd DFFPOSX1
X_11725_ _11725_/A _11725_/Y vdd gnd INVX1
XFILL_2__11070_ vdd gnd FILL
XFILL_1__10820_ vdd gnd FILL
X_14444_ _14444_/A _14444_/Y vdd gnd INVX1
X_11656_ _11656_/D _11656_/CLK _11656_/Q vdd gnd DFFPOSX1
XFILL_0__11200_ vdd gnd FILL
XFILL_0__12180_ vdd gnd FILL
X_10607_ _10607_/A _10607_/B _10607_/Y vdd gnd NAND2X1
X_14375_ _14375_/A _14375_/B _14375_/C _14375_/Y vdd gnd NAND3X1
XFILL_2__8703_ vdd gnd FILL
X_11587_ _11587_/A _11587_/B _11587_/C _11587_/Y vdd gnd OAI21X1
XFILL_0__11131_ vdd gnd FILL
XFILL_1__10682_ vdd gnd FILL
X_13326_ _13326_/A _13326_/B _13326_/C _13326_/Y vdd gnd AOI21X1
X_10538_ _10538_/A _10538_/Y vdd gnd INVX1
XFILL_2__8634_ vdd gnd FILL
XFILL_2__14760_ vdd gnd FILL
XFILL_1__12421_ vdd gnd FILL
XFILL_0__11062_ vdd gnd FILL
XFILL_2__11972_ vdd gnd FILL
X_13257_ _13257_/A _13257_/B _13257_/C _13257_/Y vdd gnd OAI21X1
X_10469_ _10469_/A _10469_/B _10469_/Y vdd gnd NOR2X1
XFILL_2__13711_ vdd gnd FILL
XFILL_0__10013_ vdd gnd FILL
XFILL_2__8565_ vdd gnd FILL
XFILL_2__14691_ vdd gnd FILL
XFILL_1__12352_ vdd gnd FILL
X_12208_ _12208_/A _12208_/B _12208_/Y vdd gnd NAND2X1
X_13188_ _13188_/A _13188_/B _13188_/Y vdd gnd AND2X2
XFILL_0__7580_ vdd gnd FILL
XFILL_2__13642_ vdd gnd FILL
XFILL_1__11303_ vdd gnd FILL
XFILL_0__14821_ vdd gnd FILL
XFILL_2__8496_ vdd gnd FILL
XFILL_1__12283_ vdd gnd FILL
X_12139_ _12139_/A _12139_/B _12139_/Y vdd gnd OR2X2
XFILL_1__14022_ vdd gnd FILL
XFILL_1__11234_ vdd gnd FILL
XFILL_0__14752_ vdd gnd FILL
XFILL_0__9250_ vdd gnd FILL
XFILL_0__11964_ vdd gnd FILL
XFILL_1__11165_ vdd gnd FILL
XFILL_0__13703_ vdd gnd FILL
XFILL_0__8201_ vdd gnd FILL
XFILL_0__10915_ vdd gnd FILL
XFILL_0__14683_ vdd gnd FILL
XFILL_2__9117_ vdd gnd FILL
XFILL_0__9181_ vdd gnd FILL
XFILL_0__11895_ vdd gnd FILL
XFILL_1__10116_ vdd gnd FILL
XFILL_0__13634_ vdd gnd FILL
XFILL_1__11096_ vdd gnd FILL
XBUFX2_insert3 BUFX2_insert3/A BUFX2_insert3/Y vdd gnd BUFX2
XFILL_0__8132_ vdd gnd FILL
XFILL_0__10846_ vdd gnd FILL
XFILL_2__9048_ vdd gnd FILL
X_8760_ _8760_/A _8760_/B _8760_/C _8760_/Y vdd gnd OAI21X1
XFILL_2__11406_ vdd gnd FILL
XFILL_1__10047_ vdd gnd FILL
XFILL_0__10777_ vdd gnd FILL
XFILL_0__13565_ vdd gnd FILL
X_7711_ _7711_/A _7711_/B _7711_/C _7711_/Y vdd gnd OAI21X1
XFILL_0__8063_ vdd gnd FILL
XFILL_2__14125_ vdd gnd FILL
X_8691_ _8691_/A _8691_/B _8691_/C _8691_/Y vdd gnd OAI21X1
XFILL_2__11337_ vdd gnd FILL
XFILL_1__14855_ vdd gnd FILL
XFILL_0__12516_ vdd gnd FILL
X_7642_ _7642_/A _7642_/B _7642_/C _7642_/Y vdd gnd OAI21X1
XFILL_1__13806_ vdd gnd FILL
XFILL_2__14056_ vdd gnd FILL
XFILL_1__14786_ vdd gnd FILL
XFILL_0__12447_ vdd gnd FILL
XFILL_1__11998_ vdd gnd FILL
XFILL_2__13007_ vdd gnd FILL
X_7573_ _7573_/A _7573_/B _7573_/C _7573_/Y vdd gnd NAND3X1
XFILL_1__13737_ vdd gnd FILL
XFILL_0__12378_ vdd gnd FILL
XFILL_1__10949_ vdd gnd FILL
X_9312_ _9312_/A _9312_/B _9312_/Y vdd gnd NAND2X1
XFILL_0__8965_ vdd gnd FILL
XFILL_0__14117_ vdd gnd FILL
XFILL_0__11329_ vdd gnd FILL
XFILL_1__13668_ vdd gnd FILL
X_9243_ _9243_/A _9243_/B _9243_/C _9243_/Y vdd gnd OAI21X1
XFILL_1__12619_ vdd gnd FILL
XFILL_0__14048_ vdd gnd FILL
XFILL_1__13599_ vdd gnd FILL
XFILL_0__7847_ vdd gnd FILL
X_9174_ _9174_/A _9174_/B _9174_/C _9174_/Y vdd gnd OAI21X1
X_8125_ _8125_/A _8125_/B _8125_/Y vdd gnd OR2X2
XFILL_0__7778_ vdd gnd FILL
XFILL_0__9517_ vdd gnd FILL
XFILL_1__8310_ vdd gnd FILL
XFILL_1__9290_ vdd gnd FILL
X_8056_ _8056_/A _8056_/Y vdd gnd INVX8
XFILL_0__9448_ vdd gnd FILL
XFILL_1__8241_ vdd gnd FILL
XFILL_0__9379_ vdd gnd FILL
XFILL_1__8172_ vdd gnd FILL
XFILL_1__7123_ vdd gnd FILL
X_8958_ _8958_/A _8958_/B _8958_/C _8958_/Y vdd gnd OAI21X1
X_7909_ _7909_/A _7909_/B _7909_/C _7909_/Y vdd gnd OAI21X1
X_8889_ _8889_/D _8889_/CLK _8889_/Q vdd gnd DFFPOSX1
XFILL_1_CLKBUF1_insert30 vdd gnd FILL
XFILL_1_CLKBUF1_insert41 vdd gnd FILL
XFILL_1_CLKBUF1_insert52 vdd gnd FILL
XFILL_1_CLKBUF1_insert63 vdd gnd FILL
XFILL_1_CLKBUF1_insert74 vdd gnd FILL
X_11510_ _11510_/A _11510_/B _11510_/Y vdd gnd AND2X2
XFILL_1_CLKBUF1_insert85 vdd gnd FILL
XFILL_1_CLKBUF1_insert96 vdd gnd FILL
X_12490_ _12490_/A _12490_/B _12490_/C _12490_/Y vdd gnd OAI21X1
X_11441_ _11441_/A _11441_/B _11441_/Y vdd gnd AND2X2
X_14160_ _14160_/D _14160_/CLK _14160_/Q vdd gnd DFFPOSX1
X_11372_ _11372_/A _11372_/Y vdd gnd INVX1
XFILL_1__7887_ vdd gnd FILL
X_13111_ _13111_/A _13111_/B _13111_/C _13111_/Y vdd gnd AOI21X1
X_10323_ _10323_/A _10323_/Y vdd gnd INVX1
X_14091_ _14091_/A _14091_/B _14091_/C _14091_/Y vdd gnd AOI21X1
XFILL_1__9626_ vdd gnd FILL
X_13042_ _13042_/A _13042_/B _13042_/Y vdd gnd NOR2X1
X_10254_ _10254_/A _10254_/B _10254_/Y vdd gnd OR2X2
XFILL_1__9557_ vdd gnd FILL
XFILL_2__8350_ vdd gnd FILL
XFILL_1__8508_ vdd gnd FILL
X_10185_ _10185_/A _10185_/B _10185_/C _10185_/Y vdd gnd NAND3X1
XFILL_1__9488_ vdd gnd FILL
XFILL_2__8281_ vdd gnd FILL
XFILL_1__8439_ vdd gnd FILL
XFILL_2__10570_ vdd gnd FILL
X_13944_ _13944_/A _13944_/B _13944_/Y vdd gnd NAND2X1
X_13875_ _13875_/A _13875_/B _13875_/Y vdd gnd NAND2X1
XFILL_0__10631_ vdd gnd FILL
XFILL_1__12970_ vdd gnd FILL
X_12826_ _12826_/A _12826_/Y vdd gnd INVX1
XFILL_1__11921_ vdd gnd FILL
XFILL_0__10562_ vdd gnd FILL
XFILL_0__13350_ vdd gnd FILL
X_12757_ _12757_/A _12757_/B _12757_/C _12757_/Y vdd gnd AOI21X1
XFILL_2__11122_ vdd gnd FILL
XFILL_1__14640_ vdd gnd FILL
XFILL_0__12301_ vdd gnd FILL
XFILL_1__11852_ vdd gnd FILL
XFILL_0__13281_ vdd gnd FILL
XFILL_0__10493_ vdd gnd FILL
X_11708_ _11708_/A _11708_/B _11708_/C _11708_/Y vdd gnd OAI21X1
X_12688_ _12688_/A _12688_/Y vdd gnd INVX1
XFILL_2__11053_ vdd gnd FILL
XFILL_0__12232_ vdd gnd FILL
XFILL_1__10803_ vdd gnd FILL
XFILL_1__14571_ vdd gnd FILL
X_14427_ _14427_/A _14427_/B _14427_/C _14427_/Y vdd gnd NAND3X1
XFILL_1__11783_ vdd gnd FILL
X_11639_ _11639_/D _11639_/CLK _11639_/Q vdd gnd DFFPOSX1
XFILL_1__13522_ vdd gnd FILL
XFILL_0__12163_ vdd gnd FILL
XFILL_0__8750_ vdd gnd FILL
X_14358_ _14358_/A _14358_/B _14358_/Y vdd gnd OR2X2
XFILL_0__11114_ vdd gnd FILL
XFILL_1__10665_ vdd gnd FILL
XFILL_0__7701_ vdd gnd FILL
XFILL_0__12094_ vdd gnd FILL
X_13309_ _13309_/A _13309_/Y vdd gnd INVX1
X_14289_ _14289_/A _14289_/B _14289_/Y vdd gnd NOR2X1
XFILL_0__8681_ vdd gnd FILL
XFILL_2__14743_ vdd gnd FILL
XFILL_2__8617_ vdd gnd FILL
XFILL_1__12404_ vdd gnd FILL
XFILL_0__11045_ vdd gnd FILL
XFILL_2__11955_ vdd gnd FILL
XFILL_1__13384_ vdd gnd FILL
XFILL_0__7632_ vdd gnd FILL
XFILL_1__10596_ vdd gnd FILL
XFILL_2__8548_ vdd gnd FILL
XFILL_2__14674_ vdd gnd FILL
XFILL_1__12335_ vdd gnd FILL
XFILL_2__11886_ vdd gnd FILL
XFILL_0__7563_ vdd gnd FILL
XFILL_2__13625_ vdd gnd FILL
XFILL_0__14804_ vdd gnd FILL
XFILL_2__8479_ vdd gnd FILL
XFILL_0__9302_ vdd gnd FILL
XFILL_1__12266_ vdd gnd FILL
X_9930_ _9930_/A _9930_/B _9930_/Y vdd gnd NAND2X1
XFILL_0__12996_ vdd gnd FILL
XFILL_1__14005_ vdd gnd FILL
XFILL_0__7494_ vdd gnd FILL
XFILL_1__11217_ vdd gnd FILL
XFILL_2__13556_ vdd gnd FILL
XFILL_0__14735_ vdd gnd FILL
XFILL_0__9233_ vdd gnd FILL
XFILL_0__11947_ vdd gnd FILL
XFILL_1__12197_ vdd gnd FILL
X_9861_ _9861_/A _9861_/B _9861_/C _9861_/Y vdd gnd AOI21X1
XFILL_1__11148_ vdd gnd FILL
XFILL_0__14666_ vdd gnd FILL
XFILL_0__9164_ vdd gnd FILL
XFILL_0__11878_ vdd gnd FILL
X_8812_ _8812_/A _8812_/B _8812_/Y vdd gnd NAND2X1
X_9792_ _9792_/D _9792_/CLK _9792_/Q vdd gnd DFFPOSX1
XFILL_1__11079_ vdd gnd FILL
XFILL_0__13617_ vdd gnd FILL
XFILL_0__10829_ vdd gnd FILL
XFILL_0__8115_ vdd gnd FILL
XFILL_0__14597_ vdd gnd FILL
XFILL_0__9095_ vdd gnd FILL
X_8743_ _8743_/A _8743_/B _8743_/C _8743_/Y vdd gnd NAND3X1
XFILL_0__13548_ vdd gnd FILL
XFILL_0__8046_ vdd gnd FILL
X_8674_ _8674_/A _8674_/B _8674_/C _8674_/Y vdd gnd OAI21X1
XFILL_1__14838_ vdd gnd FILL
X_7625_ _7625_/A _7625_/B _7625_/C _7625_/Y vdd gnd OAI21X1
XFILL_2__14039_ vdd gnd FILL
XFILL_1__14769_ vdd gnd FILL
XFILL_1__7810_ vdd gnd FILL
X_7556_ _7556_/A _7556_/B _7556_/Y vdd gnd NAND2X1
XFILL_1__8790_ vdd gnd FILL
XFILL_0__9997_ vdd gnd FILL
XFILL_1_CLKBUF1_insert107 vdd gnd FILL
XFILL256350x108150 vdd gnd FILL
XFILL_1__7741_ vdd gnd FILL
XFILL_0__8948_ vdd gnd FILL
X_7487_ _7487_/A _7487_/B _7487_/Y vdd gnd NAND2X1
X_9226_ _9226_/A _9226_/Y vdd gnd INVX1
XFILL_1__7672_ vdd gnd FILL
XFILL_1__9411_ vdd gnd FILL
X_9157_ _9157_/A _9157_/B _9157_/C _9157_/Y vdd gnd NAND3X1
XFILL_1__9342_ vdd gnd FILL
X_8108_ _8108_/A _8108_/B _8108_/C _8108_/Y vdd gnd OAI21X1
X_9088_ _9088_/A _9088_/B _9088_/Y vdd gnd NAND2X1
XFILL_1__9273_ vdd gnd FILL
X_8039_ _8039_/A _8039_/B _8039_/C _8039_/Y vdd gnd OAI21X1
XFILL_1__8224_ vdd gnd FILL
X_11990_ _11990_/A _11990_/B _11990_/C _11990_/D _11990_/Y vdd gnd AOI22X1
X_10941_ _10941_/A _10941_/B _10941_/C _10941_/Y vdd gnd OAI21X1
XFILL_1__8155_ vdd gnd FILL
X_13660_ _13660_/A _13660_/B _13660_/C _13660_/Y vdd gnd NAND3X1
XFILL_1__7106_ vdd gnd FILL
X_10872_ _10872_/A _10872_/B _10872_/Y vdd gnd NAND2X1
XFILL_1__8086_ vdd gnd FILL
X_12611_ _12611_/D _12611_/CLK _12611_/Q vdd gnd DFFPOSX1
X_13591_ _13591_/A _13591_/B _13591_/C _13591_/Y vdd gnd OAI21X1
X_12542_ _12542_/D _12542_/CLK _12542_/Q vdd gnd DFFPOSX1
X_12473_ _12473_/A _12473_/B _12473_/C _12473_/Y vdd gnd OAI21X1
XFILL_1__8988_ vdd gnd FILL
X_14212_ _14212_/D _14212_/CLK _14212_/Q vdd gnd DFFPOSX1
X_11424_ _11424_/A _11424_/B _11424_/C _11424_/Y vdd gnd OAI21X1
X_14143_ _14143_/A _14143_/B _14143_/Y vdd gnd NAND2X1
X_11355_ _11355_/A _11355_/B _11355_/C _11355_/Y vdd gnd OAI21X1
XFILL_1__10450_ vdd gnd FILL
X_10306_ _10306_/A _10306_/B _10306_/Y vdd gnd NAND2X1
X_14074_ _14074_/A _14074_/B _14074_/C _14074_/Y vdd gnd OAI21X1
XCLKBUF1_insert106 CLKBUF1_insert106/A CLKBUF1_insert106/Y vdd gnd CLKBUF1
XFILL_1__9609_ vdd gnd FILL
X_11286_ _11286_/A _11286_/B _11286_/Y vdd gnd AND2X2
XFILL_1__10381_ vdd gnd FILL
X_13025_ _13025_/A _13025_/B _13025_/Y vdd gnd NAND2X1
X_10237_ _10237_/A _10237_/B _10237_/Y vdd gnd NAND2X1
XFILL_1__12120_ vdd gnd FILL
XFILL_0__12850_ vdd gnd FILL
X_10168_ _10168_/A _10168_/Y vdd gnd INVX1
XFILL_2__13410_ vdd gnd FILL
XFILL_1__12051_ vdd gnd FILL
XFILL_2__14390_ vdd gnd FILL
XFILL_0__11801_ vdd gnd FILL
XFILL_0__12781_ vdd gnd FILL
XFILL_2__7215_ vdd gnd FILL
XFILL_1__11002_ vdd gnd FILL
X_10099_ _10099_/A _10099_/B _10099_/C _10099_/Y vdd gnd AOI21X1
XFILL_2__13341_ vdd gnd FILL
XFILL_0__11732_ vdd gnd FILL
X_13927_ _13927_/A _13927_/B _13927_/Y vdd gnd NOR2X1
XFILL_2__7146_ vdd gnd FILL
XFILL_2__13272_ vdd gnd FILL
XFILL_2__10484_ vdd gnd FILL
XFILL_0__14451_ vdd gnd FILL
X_13858_ _13858_/A _13858_/B _13858_/C _13858_/Y vdd gnd OAI21X1
XFILL_0__13402_ vdd gnd FILL
XFILL_1__12953_ vdd gnd FILL
XFILL256950x57750 vdd gnd FILL
XFILL_0__10614_ vdd gnd FILL
XFILL_0__14382_ vdd gnd FILL
XFILL_0__11594_ vdd gnd FILL
XFILL_1_BUFX2_insert250 vdd gnd FILL
X_12809_ _12809_/A _12809_/B _12809_/Y vdd gnd NOR2X1
XFILL_1_BUFX2_insert261 vdd gnd FILL
XFILL_1_BUFX2_insert272 vdd gnd FILL
XFILL_1__11904_ vdd gnd FILL
X_13789_ _13789_/A _13789_/B _13789_/C _13789_/Y vdd gnd OAI21X1
XFILL_0__10545_ vdd gnd FILL
XCLKBUF1_insert32 CLKBUF1_insert32/A CLKBUF1_insert32/Y vdd gnd CLKBUF1
XFILL_0__13333_ vdd gnd FILL
XFILL_1_BUFX2_insert283 vdd gnd FILL
XFILL_1__12884_ vdd gnd FILL
XFILL_1_BUFX2_insert294 vdd gnd FILL
XCLKBUF1_insert43 CLKBUF1_insert43/A CLKBUF1_insert43/Y vdd gnd CLKBUF1
XFILL_0__9920_ vdd gnd FILL
XCLKBUF1_insert54 CLKBUF1_insert54/A CLKBUF1_insert54/Y vdd gnd CLKBUF1
XFILL_2__11105_ vdd gnd FILL
XCLKBUF1_insert65 CLKBUF1_insert65/A CLKBUF1_insert65/Y vdd gnd CLKBUF1
XFILL_1__14623_ vdd gnd FILL
XCLKBUF1_insert76 CLKBUF1_insert76/A CLKBUF1_insert76/Y vdd gnd CLKBUF1
XFILL_1__11835_ vdd gnd FILL
XFILL_0__10476_ vdd gnd FILL
XCLKBUF1_insert87 CLKBUF1_insert87/A CLKBUF1_insert87/Y vdd gnd CLKBUF1
XFILL_0__13264_ vdd gnd FILL
X_7410_ _7410_/A _7410_/B _7410_/C _7410_/Y vdd gnd NAND3X1
XCLKBUF1_insert98 CLKBUF1_insert98/A CLKBUF1_insert98/Y vdd gnd CLKBUF1
XFILL_0__9851_ vdd gnd FILL
XFILL_2__11036_ vdd gnd FILL
X_8390_ _8390_/A _8390_/B _8390_/C _8390_/Y vdd gnd OAI21X1
XFILL_0__12215_ vdd gnd FILL
XFILL_0__13195_ vdd gnd FILL
XFILL_1__11766_ vdd gnd FILL
XFILL_0__8802_ vdd gnd FILL
X_7341_ _7341_/A _7341_/B _7341_/C _7341_/Y vdd gnd NAND3X1
XFILL_1__13505_ vdd gnd FILL
XFILL_1__14485_ vdd gnd FILL
XFILL_0__12146_ vdd gnd FILL
XFILL_0__8733_ vdd gnd FILL
XFILL_1__11697_ vdd gnd FILL
X_7272_ _7272_/A _7272_/B _7272_/Y vdd gnd NOR2X1
XFILL_1__10648_ vdd gnd FILL
XFILL_0__12077_ vdd gnd FILL
X_9011_ _9011_/A _9011_/Y vdd gnd INVX2
XFILL_0__8664_ vdd gnd FILL
XFILL_0__11028_ vdd gnd FILL
XFILL_2__11938_ vdd gnd FILL
XFILL_1__13367_ vdd gnd FILL
XFILL_0__7615_ vdd gnd FILL
XFILL_1__10579_ vdd gnd FILL
XFILL_0__8595_ vdd gnd FILL
XFILL_1__12318_ vdd gnd FILL
XFILL_2__11869_ vdd gnd FILL
XFILL_1__13298_ vdd gnd FILL
XFILL_0__7546_ vdd gnd FILL
XFILL_2__13608_ vdd gnd FILL
XFILL_1__12249_ vdd gnd FILL
X_9913_ _9913_/A _9913_/Y vdd gnd INVX1
XFILL_0__12979_ vdd gnd FILL
XFILL_0__7477_ vdd gnd FILL
XFILL_2__13539_ vdd gnd FILL
XFILL_0__14718_ vdd gnd FILL
XFILL_0__9216_ vdd gnd FILL
X_9844_ _9844_/A _9844_/Y vdd gnd INVX1
XFILL_0__14649_ vdd gnd FILL
XFILL_0__9147_ vdd gnd FILL
X_9775_ _9775_/D _9775_/CLK _9775_/Q vdd gnd DFFPOSX1
XFILL_0__9078_ vdd gnd FILL
X_8726_ _8726_/A _8726_/B _8726_/Y vdd gnd NOR2X1
XFILL_1__9960_ vdd gnd FILL
XFILL_0__8029_ vdd gnd FILL
X_8657_ _8657_/A _8657_/B _8657_/C _8657_/Y vdd gnd OAI21X1
XFILL_1__9891_ vdd gnd FILL
X_7608_ _7608_/A _7608_/B _7608_/Y vdd gnd NAND2X1
X_8588_ _8588_/A _8588_/B _8588_/Y vdd gnd NAND2X1
X_7539_ _7539_/A _7539_/B _7539_/Y vdd gnd OR2X2
XFILL_1__8773_ vdd gnd FILL
XFILL_1__7724_ vdd gnd FILL
X_11140_ _11140_/A _11140_/B _11140_/C _11140_/Y vdd gnd OAI21X1
X_9209_ _9209_/A _9209_/B _9209_/C _9209_/Y vdd gnd OAI21X1
XFILL_1__7655_ vdd gnd FILL
X_11071_ _11071_/A _11071_/B _11071_/C _11071_/Y vdd gnd OAI21X1
XFILL_1__7586_ vdd gnd FILL
X_10022_ _10022_/A _10022_/B _10022_/C _10022_/Y vdd gnd NAND3X1
XFILL_1__9325_ vdd gnd FILL
X_14830_ _14830_/A _14830_/B _14830_/C _14830_/Y vdd gnd OAI21X1
XFILL_1__9256_ vdd gnd FILL
XFILL_1__8207_ vdd gnd FILL
X_14761_ _14761_/A _14761_/B _14761_/C _14761_/Y vdd gnd AOI21X1
X_11973_ _11973_/A _11973_/B _11973_/Y vdd gnd NOR2X1
XFILL_1__9187_ vdd gnd FILL
X_10924_ _10924_/A _10924_/Y vdd gnd INVX2
X_13712_ _13712_/A _13712_/B _13712_/C _13712_/Y vdd gnd OAI21X1
X_14692_ _14692_/A _14692_/B _14692_/Y vdd gnd NAND2X1
XFILL_1__8138_ vdd gnd FILL
X_13643_ _13643_/A _13643_/B _13643_/C _13643_/Y vdd gnd OAI21X1
X_10855_ _10855_/A _10855_/B _10855_/Y vdd gnd NOR2X1
XFILL_1__8069_ vdd gnd FILL
XFILL_0_BUFX2_insert202 vdd gnd FILL
X_13574_ _13574_/A _13574_/B _13574_/S _13574_/Y vdd gnd MUX2X1
XFILL_0_BUFX2_insert213 vdd gnd FILL
X_10786_ _10786_/A _10786_/Y vdd gnd INVX1
XFILL_0__10330_ vdd gnd FILL
XFILL_0_BUFX2_insert224 vdd gnd FILL
XFILL_0_BUFX2_insert235 vdd gnd FILL
XFILL_0_BUFX2_insert246 vdd gnd FILL
X_12525_ _12525_/A _12525_/B _12525_/C _12525_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert257 vdd gnd FILL
XFILL_0_BUFX2_insert268 vdd gnd FILL
XFILL_0_BUFX2_insert279 vdd gnd FILL
XFILL_0__10261_ vdd gnd FILL
X_12456_ _12456_/A _12456_/B _12456_/C _12456_/Y vdd gnd OAI21X1
XFILL_2__12910_ vdd gnd FILL
XFILL_0__12000_ vdd gnd FILL
XFILL_1__11551_ vdd gnd FILL
XFILL_0__10192_ vdd gnd FILL
X_11407_ _11407_/A _11407_/B _11407_/C _11407_/Y vdd gnd OAI21X1
XFILL_2__9503_ vdd gnd FILL
X_12387_ _12387_/A _12387_/B _12387_/C _12387_/Y vdd gnd OAI21X1
XFILL_1__10502_ vdd gnd FILL
XFILL_2__12841_ vdd gnd FILL
XFILL_1__14270_ vdd gnd FILL
XFILL_1__11482_ vdd gnd FILL
X_14126_ _14126_/A _14126_/B _14126_/C _14126_/Y vdd gnd OAI21X1
X_11338_ _11338_/A _11338_/B _11338_/C _11338_/Y vdd gnd OAI21X1
XFILL_2_BUFX2_insert17 vdd gnd FILL
XFILL_1__13221_ vdd gnd FILL
XFILL_2__9434_ vdd gnd FILL
XFILL_1__10433_ vdd gnd FILL
XFILL_2__12772_ vdd gnd FILL
XFILL_0__13951_ vdd gnd FILL
X_14057_ _14057_/A _14057_/Y vdd gnd INVX1
X_11269_ _11269_/A _11269_/B _11269_/C _11269_/Y vdd gnd NAND3X1
XFILL_2__9365_ vdd gnd FILL
XFILL_1__13152_ vdd gnd FILL
XFILL_0__12902_ vdd gnd FILL
XFILL_1__10364_ vdd gnd FILL
XFILL_0__7400_ vdd gnd FILL
X_13008_ _13008_/A _13008_/B _13008_/C _13008_/Y vdd gnd OAI21X1
XFILL_0__13882_ vdd gnd FILL
XFILL_0__8380_ vdd gnd FILL
XFILL_1__12103_ vdd gnd FILL
XFILL_2__14442_ vdd gnd FILL
XFILL_1__13083_ vdd gnd FILL
XFILL_0__12833_ vdd gnd FILL
XFILL_1__10295_ vdd gnd FILL
XFILL_0__7331_ vdd gnd FILL
XFILL_1__12034_ vdd gnd FILL
XFILL_2__14373_ vdd gnd FILL
XFILL_0__12764_ vdd gnd FILL
XFILL_0__7262_ vdd gnd FILL
XFILL_2__13324_ vdd gnd FILL
X_7890_ _7890_/A _7890_/B _7890_/Y vdd gnd NAND2X1
XFILL_0__9001_ vdd gnd FILL
XFILL_0__11715_ vdd gnd FILL
XFILL_0__12695_ vdd gnd FILL
XFILL_0__7193_ vdd gnd FILL
XFILL_2__7129_ vdd gnd FILL
XFILL_2__13255_ vdd gnd FILL
XFILL_0__14434_ vdd gnd FILL
XFILL_1__13985_ vdd gnd FILL
X_9560_ _9560_/A _9560_/B _9560_/S _9560_/Y vdd gnd MUX2X1
XFILL_2__13186_ vdd gnd FILL
XFILL_1__12936_ vdd gnd FILL
XFILL_0__14365_ vdd gnd FILL
X_8511_ _8511_/A _8511_/B _8511_/C _8511_/Y vdd gnd OAI21X1
XFILL_0__11577_ vdd gnd FILL
X_9491_ _9491_/A _9491_/Y vdd gnd INVX1
XFILL_0__13316_ vdd gnd FILL
XFILL_0__10528_ vdd gnd FILL
XFILL_1__12867_ vdd gnd FILL
XFILL_0__9903_ vdd gnd FILL
XFILL_0__14296_ vdd gnd FILL
X_8442_ _8442_/A _8442_/B _8442_/C _8442_/Y vdd gnd OAI21X1
XFILL_1__14606_ vdd gnd FILL
XFILL_1__11818_ vdd gnd FILL
XFILL_0__13247_ vdd gnd FILL
XFILL_0__10459_ vdd gnd FILL
XFILL_1__12798_ vdd gnd FILL
X_8373_ _8373_/A _8373_/B _8373_/Y vdd gnd AND2X2
XFILL_1__11749_ vdd gnd FILL
XFILL_0__13178_ vdd gnd FILL
X_7324_ _7324_/A _7324_/B _7324_/C _7324_/Y vdd gnd NAND3X1
XFILL_1__14468_ vdd gnd FILL
XFILL_0__12129_ vdd gnd FILL
XFILL_0__8716_ vdd gnd FILL
X_7255_ _7255_/A _7255_/B _7255_/C _7255_/Y vdd gnd OAI21X1
XFILL_0__9696_ vdd gnd FILL
XFILL_1__13419_ vdd gnd FILL
XFILL_1__14399_ vdd gnd FILL
XFILL_1__7440_ vdd gnd FILL
XFILL_0__8647_ vdd gnd FILL
X_7186_ _7186_/A _7186_/B _7186_/S _7186_/Y vdd gnd MUX2X1
XFILL_1__7371_ vdd gnd FILL
XFILL_0__8578_ vdd gnd FILL
XFILL_1__9110_ vdd gnd FILL
XFILL_0__7529_ vdd gnd FILL
XFILL_2_BUFX2_insert308 vdd gnd FILL
XFILL_1_BUFX2_insert3 vdd gnd FILL
XFILL_1__9041_ vdd gnd FILL
X_9827_ _9827_/D _9827_/CLK _9827_/Q vdd gnd DFFPOSX1
X_9758_ _9758_/A _9758_/B _9758_/C _9758_/Y vdd gnd OAI21X1
X_10640_ _10640_/A _10640_/Y vdd gnd INVX1
XBUFX2_insert307 BUFX2_insert307/A BUFX2_insert307/Y vdd gnd BUFX2
XBUFX2_insert318 BUFX2_insert318/A BUFX2_insert318/Y vdd gnd BUFX2
X_8709_ _8709_/A _8709_/B _8709_/Y vdd gnd OR2X2
XBUFX2_insert329 BUFX2_insert329/A BUFX2_insert329/Y vdd gnd BUFX2
XFILL_1__9943_ vdd gnd FILL
X_9689_ _9689_/A _9689_/B _9689_/C _9689_/Y vdd gnd OAI21X1
X_10571_ _10571_/A _10571_/B _10571_/C _10571_/Y vdd gnd AOI21X1
XFILL_1__9874_ vdd gnd FILL
X_12310_ _12310_/A _12310_/B _12310_/Y vdd gnd NAND2X1
X_13290_ _13290_/A _13290_/Y vdd gnd INVX1
XFILL_1__8825_ vdd gnd FILL
X_12241_ _12241_/A _12241_/B _12241_/C _12241_/Y vdd gnd AOI21X1
XFILL_1__8756_ vdd gnd FILL
X_12172_ _12172_/A _12172_/B _12172_/C _12172_/Y vdd gnd OAI21X1
XFILL_1__7707_ vdd gnd FILL
XFILL_1__8687_ vdd gnd FILL
X_11123_ _11123_/A _11123_/B _11123_/Y vdd gnd NAND2X1
XFILL_1__7638_ vdd gnd FILL
X_11054_ _11054_/A _11054_/B _11054_/C _11054_/Y vdd gnd NAND3X1
XFILL_2__9150_ vdd gnd FILL
XFILL_1__7569_ vdd gnd FILL
X_10005_ _10005_/A _10005_/B _10005_/C _10005_/Y vdd gnd OAI21X1
XFILL_1__9308_ vdd gnd FILL
XFILL_2__9081_ vdd gnd FILL
XFILL_1__10080_ vdd gnd FILL
X_14813_ _14813_/A _14813_/B _14813_/Y vdd gnd OR2X2
XFILL_1__9239_ vdd gnd FILL
XFILL_2__11370_ vdd gnd FILL
X_14744_ _14744_/A _14744_/B _14744_/Y vdd gnd NAND2X1
X_11956_ _11956_/A _11956_/B _11956_/C _11956_/Y vdd gnd OAI21X1
XFILL_0__11500_ vdd gnd FILL
XFILL_0__12480_ vdd gnd FILL
X_10907_ _10907_/A _10907_/B _10907_/S _10907_/Y vdd gnd MUX2X1
X_14675_ _14675_/A _14675_/B _14675_/Y vdd gnd NAND2X1
X_11887_ _11887_/A _11887_/B _11887_/C _11887_/Y vdd gnd OAI21X1
XFILL_2__9983_ vdd gnd FILL
XFILL_0__11431_ vdd gnd FILL
XFILL_1__13770_ vdd gnd FILL
XFILL_1__10982_ vdd gnd FILL
X_10838_ _10838_/A _10838_/B _10838_/Y vdd gnd NAND2X1
X_13626_ _13626_/A _13626_/B _13626_/Y vdd gnd NAND2X1
XFILL_1__12721_ vdd gnd FILL
XFILL_0__14150_ vdd gnd FILL
XFILL_0__11362_ vdd gnd FILL
X_10769_ _10769_/A _10769_/Y vdd gnd INVX2
X_13557_ _13557_/A _13557_/B _13557_/C _13557_/Y vdd gnd OAI21X1
XFILL_0__13101_ vdd gnd FILL
XFILL_1__12652_ vdd gnd FILL
XFILL_0__10313_ vdd gnd FILL
XFILL_0__11293_ vdd gnd FILL
XFILL_0__14081_ vdd gnd FILL
X_12508_ _12508_/A _12508_/B _12508_/Y vdd gnd NAND2X1
XFILL_0__7880_ vdd gnd FILL
X_13488_ _13488_/D _13488_/CLK _13488_/Q vdd gnd DFFPOSX1
XFILL_1__11603_ vdd gnd FILL
XFILL_0__10244_ vdd gnd FILL
XFILL_2__13942_ vdd gnd FILL
XFILL_0__13032_ vdd gnd FILL
XFILL_2__8796_ vdd gnd FILL
X_12439_ _12439_/A _12439_/B _12439_/C _12439_/Y vdd gnd NAND3X1
XFILL_1__14322_ vdd gnd FILL
XFILL_1__11534_ vdd gnd FILL
XFILL_2__13873_ vdd gnd FILL
XFILL_0__10175_ vdd gnd FILL
XFILL_0__9550_ vdd gnd FILL
XFILL_1__14253_ vdd gnd FILL
XFILL_2__12824_ vdd gnd FILL
XFILL_1__11465_ vdd gnd FILL
XFILL_0__8501_ vdd gnd FILL
X_14109_ _14109_/A _14109_/B _14109_/C _14109_/Y vdd gnd OAI21X1
XFILL_0__9481_ vdd gnd FILL
XFILL_1__13204_ vdd gnd FILL
XFILL_2__9417_ vdd gnd FILL
XFILL_1__10416_ vdd gnd FILL
XFILL_2__12755_ vdd gnd FILL
XFILL_0__13934_ vdd gnd FILL
XFILL_0__8432_ vdd gnd FILL
XFILL_1__11396_ vdd gnd FILL
XFILL_1__13135_ vdd gnd FILL
XFILL_2__9348_ vdd gnd FILL
XFILL_1__10347_ vdd gnd FILL
XFILL_2__12686_ vdd gnd FILL
XFILL_0__13865_ vdd gnd FILL
XFILL_0__8363_ vdd gnd FILL
X_8991_ _8991_/A _8991_/B _8991_/C _8991_/Y vdd gnd OAI21X1
XFILL_2__14425_ vdd gnd FILL
XFILL_2__9279_ vdd gnd FILL
XFILL_0__12816_ vdd gnd FILL
XFILL_1__13066_ vdd gnd FILL
XFILL_0__7314_ vdd gnd FILL
XFILL_1__10278_ vdd gnd FILL
XFILL_0__13796_ vdd gnd FILL
X_7942_ _7942_/D _7942_/CLK _7942_/Q vdd gnd DFFPOSX1
XFILL_0__8294_ vdd gnd FILL
XFILL_1__12017_ vdd gnd FILL
XFILL_2__14356_ vdd gnd FILL
XFILL_2__11568_ vdd gnd FILL
XFILL_0__12747_ vdd gnd FILL
XFILL_0__7245_ vdd gnd FILL
X_7873_ _7873_/A _7873_/B _7873_/C _7873_/Y vdd gnd OAI21X1
XFILL_2__14287_ vdd gnd FILL
XFILL_2__11499_ vdd gnd FILL
X_9612_ _9612_/A _9612_/B _9612_/Y vdd gnd NAND2X1
XFILL_0__12678_ vdd gnd FILL
XFILL_0__7176_ vdd gnd FILL
XFILL_0__14417_ vdd gnd FILL
XFILL_1__13968_ vdd gnd FILL
X_9543_ _9543_/A _9543_/B _9543_/Y vdd gnd NOR2X1
XFILL_1__12919_ vdd gnd FILL
XFILL_0__14348_ vdd gnd FILL
XFILL_1__13899_ vdd gnd FILL
X_9474_ _9474_/A _9474_/Y vdd gnd INVX1
XFILL_0__14279_ vdd gnd FILL
X_8425_ _8425_/A _8425_/Y vdd gnd INVX1
XFILL_1__8610_ vdd gnd FILL
XFILL_1__9590_ vdd gnd FILL
X_8356_ _8356_/A _8356_/B _8356_/C _8356_/Y vdd gnd OAI21X1
X_7307_ _7307_/A _7307_/B _7307_/C _7307_/Y vdd gnd OAI21X1
XFILL_0__9748_ vdd gnd FILL
XFILL_1__8541_ vdd gnd FILL
X_8287_ _8287_/A _8287_/B _8287_/C _8287_/Y vdd gnd NAND3X1
X_7238_ _7238_/A _7238_/B _7238_/Y vdd gnd NAND2X1
XFILL_1__8472_ vdd gnd FILL
XFILL_0__9679_ vdd gnd FILL
XFILL_1__7423_ vdd gnd FILL
X_7169_ _7169_/A _7169_/B _7169_/C _7169_/D _7169_/Y vdd gnd OAI22X1
XFILL_1__7354_ vdd gnd FILL
XFILL_2_BUFX2_insert127 vdd gnd FILL
XFILL_1__7285_ vdd gnd FILL
XFILL_1__9024_ vdd gnd FILL
X_11810_ _11810_/A _11810_/B _11810_/S _11810_/Y vdd gnd MUX2X1
X_12790_ _12790_/A _12790_/B _12790_/Y vdd gnd NAND2X1
X_11741_ _11741_/A _11741_/B _11741_/C _11741_/D _11741_/Y vdd gnd AOI22X1
X_14460_ _14460_/A _14460_/B _14460_/C _14460_/Y vdd gnd OAI21X1
X_11672_ _11672_/D _11672_/CLK _11672_/Q vdd gnd DFFPOSX1
XBUFX2_insert115 BUFX2_insert115/A BUFX2_insert115/Y vdd gnd BUFX2
XBUFX2_insert126 BUFX2_insert126/A BUFX2_insert126/Y vdd gnd BUFX2
XBUFX2_insert137 BUFX2_insert137/A BUFX2_insert137/Y vdd gnd BUFX2
X_10623_ _10623_/A _10623_/B _10623_/Y vdd gnd AND2X2
X_13411_ _13411_/A _13411_/B _13411_/C _13411_/Y vdd gnd OAI21X1
XBUFX2_insert148 BUFX2_insert148/A BUFX2_insert148/Y vdd gnd BUFX2
X_14391_ _14391_/A _14391_/B _14391_/C _14391_/Y vdd gnd NAND3X1
XFILL_1__9926_ vdd gnd FILL
XBUFX2_insert159 BUFX2_insert159/A BUFX2_insert159/Y vdd gnd BUFX2
X_13342_ _13342_/A _13342_/B _13342_/C _13342_/Y vdd gnd OAI21X1
X_10554_ _10554_/A _10554_/B _10554_/Y vdd gnd NAND2X1
XFILL_1__9857_ vdd gnd FILL
X_13273_ _13273_/A _13273_/B _13273_/C _13273_/Y vdd gnd OAI21X1
XFILL_2__7601_ vdd gnd FILL
X_10485_ _10485_/A _10485_/B _10485_/Y vdd gnd NAND2X1
XFILL_1__8808_ vdd gnd FILL
X_12224_ _12224_/A _12224_/B _12224_/C _12224_/Y vdd gnd OAI21X1
XFILL_2__7532_ vdd gnd FILL
XFILL_1__8739_ vdd gnd FILL
XFILL_2__10870_ vdd gnd FILL
X_12155_ _12155_/A _12155_/B _12155_/C _12155_/Y vdd gnd OAI21X1
XFILL_2__7463_ vdd gnd FILL
XFILL_1__11250_ vdd gnd FILL
X_11106_ _11106_/A _11106_/B _11106_/C _11106_/Y vdd gnd NAND3X1
XFILL_0__11980_ vdd gnd FILL
X_12086_ _12086_/A _12086_/B _12086_/C _12086_/Y vdd gnd OAI21X1
XFILL_1__10201_ vdd gnd FILL
XFILL_1__11181_ vdd gnd FILL
XFILL_0__10931_ vdd gnd FILL
X_11037_ _11037_/A _11037_/B _11037_/C _11037_/Y vdd gnd NAND3X1
XFILL_2__9133_ vdd gnd FILL
XFILL_1__10132_ vdd gnd FILL
XFILL_0__13650_ vdd gnd FILL
XFILL_0__10862_ vdd gnd FILL
XFILL_2__9064_ vdd gnd FILL
XFILL_2__11422_ vdd gnd FILL
XFILL_1__10063_ vdd gnd FILL
XFILL_0__13581_ vdd gnd FILL
XFILL_0__10793_ vdd gnd FILL
XFILL_2__11353_ vdd gnd FILL
X_12988_ _12988_/A _12988_/B _12988_/Y vdd gnd NAND2X1
XFILL_0__12532_ vdd gnd FILL
X_14727_ _14727_/A _14727_/B _14727_/Y vdd gnd NOR2X1
X_11939_ _11939_/A _11939_/B _11939_/C _11939_/Y vdd gnd OAI21X1
XFILL_1__13822_ vdd gnd FILL
XFILL_2__11284_ vdd gnd FILL
XFILL_0__12463_ vdd gnd FILL
X_14658_ _14658_/A _14658_/Y vdd gnd INVX1
XFILL_2__9966_ vdd gnd FILL
XFILL_0__11414_ vdd gnd FILL
XFILL_1__13753_ vdd gnd FILL
XFILL_1__10965_ vdd gnd FILL
X_13609_ _13609_/A _13609_/B _13609_/C _13609_/Y vdd gnd OAI21X1
XFILL_0__12394_ vdd gnd FILL
XFILL_0__8981_ vdd gnd FILL
X_14589_ _14589_/A _14589_/B _14589_/Y vdd gnd NAND2X1
XFILL_1__12704_ vdd gnd FILL
XFILL_0__14133_ vdd gnd FILL
XFILL_2__9897_ vdd gnd FILL
XFILL_0__11345_ vdd gnd FILL
XFILL_1__13684_ vdd gnd FILL
XFILL_1__10896_ vdd gnd FILL
XFILL_1__12635_ vdd gnd FILL
XFILL_0__14064_ vdd gnd FILL
X_8210_ _8210_/A _8210_/B _8210_/C _8210_/Y vdd gnd OAI21X1
XFILL_0__11276_ vdd gnd FILL
XFILL_0__7863_ vdd gnd FILL
X_9190_ _9190_/A _9190_/B _9190_/Y vdd gnd NAND2X1
XFILL_2__13925_ vdd gnd FILL
XFILL_0__13015_ vdd gnd FILL
XFILL_0__10227_ vdd gnd FILL
XFILL_2__8779_ vdd gnd FILL
XFILL_0__9602_ vdd gnd FILL
X_8141_ _8141_/A _8141_/Y vdd gnd INVX1
XFILL256050x252150 vdd gnd FILL
XFILL_0__7794_ vdd gnd FILL
XFILL_1__14305_ vdd gnd FILL
XFILL_1__11517_ vdd gnd FILL
XFILL_0__10158_ vdd gnd FILL
XFILL_2__13856_ vdd gnd FILL
XFILL_1__12497_ vdd gnd FILL
XFILL_0__9533_ vdd gnd FILL
X_8072_ _8072_/A _8072_/B _8072_/S _8072_/Y vdd gnd MUX2X1
XFILL_1__14236_ vdd gnd FILL
XFILL_2__12807_ vdd gnd FILL
XFILL_1__11448_ vdd gnd FILL
XFILL_0__10089_ vdd gnd FILL
XFILL_2__13787_ vdd gnd FILL
XFILL_0__9464_ vdd gnd FILL
XFILL_0__13917_ vdd gnd FILL
XFILL_2__12738_ vdd gnd FILL
XFILL_1__11379_ vdd gnd FILL
XFILL_0__8415_ vdd gnd FILL
XFILL_0__9395_ vdd gnd FILL
XFILL_1__13118_ vdd gnd FILL
XFILL_1__14098_ vdd gnd FILL
XFILL_0__13848_ vdd gnd FILL
XFILL_2__12669_ vdd gnd FILL
XFILL_0__8346_ vdd gnd FILL
X_8974_ _8974_/A _8974_/B _8974_/C _8974_/D _8974_/Y vdd gnd AOI22X1
XFILL_1__13049_ vdd gnd FILL
XFILL_0__13779_ vdd gnd FILL
X_7925_ _7925_/D _7925_/CLK _7925_/Q vdd gnd DFFPOSX1
XFILL_0__8277_ vdd gnd FILL
XFILL_0__7228_ vdd gnd FILL
X_7856_ _7856_/A _7856_/B _7856_/C _7856_/Y vdd gnd OAI21X1
XFILL_0__7159_ vdd gnd FILL
X_7787_ _7787_/A _7787_/B _7787_/Y vdd gnd NOR2X1
X_9526_ _9526_/A _9526_/B _9526_/Y vdd gnd NAND2X1
XFILL_1__9711_ vdd gnd FILL
X_9457_ _9457_/A _9457_/B _9457_/C _9457_/Y vdd gnd NAND3X1
X_8408_ _8408_/A _8408_/B _8408_/C _8408_/Y vdd gnd OAI21X1
XFILL_1__9642_ vdd gnd FILL
X_9388_ _9388_/A _9388_/B _9388_/Y vdd gnd NOR2X1
X_10270_ _10270_/A _10270_/B _10270_/C _10270_/Y vdd gnd AOI21X1
X_8339_ _8339_/A _8339_/B _8339_/C _8339_/Y vdd gnd OAI21X1
XFILL_1__9573_ vdd gnd FILL
XFILL_1__8524_ vdd gnd FILL
XFILL_1__8455_ vdd gnd FILL
X_13960_ _13960_/A _13960_/B _13960_/Y vdd gnd NAND2X1
XFILL_1__7406_ vdd gnd FILL
XFILL_1__8386_ vdd gnd FILL
X_12911_ _12911_/A _12911_/B _12911_/C _12911_/Y vdd gnd NAND3X1
XFILL257550x39750 vdd gnd FILL
XFILL_1__7337_ vdd gnd FILL
X_13891_ _13891_/A _13891_/B _13891_/C _13891_/Y vdd gnd AOI21X1
X_12842_ _12842_/A _12842_/B _12842_/C _12842_/Y vdd gnd NAND3X1
XFILL_1__7268_ vdd gnd FILL
XFILL_1__9007_ vdd gnd FILL
X_12773_ _12773_/A _12773_/B _12773_/C _12773_/Y vdd gnd NAND3X1
XFILL_1__7199_ vdd gnd FILL
X_14512_ _14512_/D _14512_/CLK _14512_/Q vdd gnd DFFPOSX1
X_11724_ _11724_/A _11724_/B _11724_/Y vdd gnd NAND2X1
XFILL257550x82950 vdd gnd FILL
X_14443_ _14443_/A _14443_/B _14443_/C _14443_/Y vdd gnd OAI21X1
X_11655_ _11655_/D _11655_/CLK _11655_/Q vdd gnd DFFPOSX1
XFILL_2__10020_ vdd gnd FILL
XFILL_2__9751_ vdd gnd FILL
X_10606_ _10606_/A _10606_/B _10606_/Y vdd gnd NOR2X1
XFILL_1__9909_ vdd gnd FILL
X_14374_ _14374_/A _14374_/B _14374_/C _14374_/Y vdd gnd OAI21X1
X_11586_ _11586_/A _11586_/B _11586_/Y vdd gnd NAND2X1
XFILL_2__9682_ vdd gnd FILL
XFILL_0__11130_ vdd gnd FILL
XFILL_1__10681_ vdd gnd FILL
X_10537_ _10537_/A _10537_/B _10537_/C _10537_/Y vdd gnd OAI21X1
X_13325_ _13325_/A _13325_/B _13325_/C _13325_/Y vdd gnd OAI21X1
XFILL_1__12420_ vdd gnd FILL
XFILL_0__11061_ vdd gnd FILL
X_10468_ _10468_/A _10468_/B _10468_/C _10468_/Y vdd gnd AOI21X1
X_13256_ _13256_/A _13256_/B _13256_/C _13256_/Y vdd gnd OAI21X1
XFILL_0__10012_ vdd gnd FILL
XFILL_2__10922_ vdd gnd FILL
XFILL_1__12351_ vdd gnd FILL
X_12207_ _12207_/A _12207_/B _12207_/C _12207_/Y vdd gnd OAI21X1
X_13187_ _13187_/A _13187_/B _13187_/Y vdd gnd NAND2X1
X_10399_ _10399_/A _10399_/B _10399_/C _10399_/Y vdd gnd NAND3X1
XFILL_2__7515_ vdd gnd FILL
XFILL_1__11302_ vdd gnd FILL
XFILL_0__14820_ vdd gnd FILL
XFILL_2__10853_ vdd gnd FILL
XFILL_1__12282_ vdd gnd FILL
X_12138_ _12138_/A _12138_/B _12138_/C _12138_/Y vdd gnd OAI21X1
XFILL_1__14021_ vdd gnd FILL
XFILL_2__7446_ vdd gnd FILL
XFILL_2__13572_ vdd gnd FILL
XFILL_1__11233_ vdd gnd FILL
XFILL_0__14751_ vdd gnd FILL
XFILL_2__10784_ vdd gnd FILL
XFILL_0__11963_ vdd gnd FILL
X_12069_ _12069_/A _12069_/B _12069_/Y vdd gnd AND2X2
XFILL_2__7377_ vdd gnd FILL
XFILL_0__13702_ vdd gnd FILL
XFILL_1__11164_ vdd gnd FILL
XFILL_0__8200_ vdd gnd FILL
XFILL_0__10914_ vdd gnd FILL
XFILL_0__14682_ vdd gnd FILL
XFILL_0__9180_ vdd gnd FILL
XFILL_0__11894_ vdd gnd FILL
XFILL_1__10115_ vdd gnd FILL
XFILL_0__13633_ vdd gnd FILL
XFILL_0__8131_ vdd gnd FILL
XFILL_0__10845_ vdd gnd FILL
XFILL_1__11095_ vdd gnd FILL
XBUFX2_insert4 BUFX2_insert4/A BUFX2_insert4/Y vdd gnd BUFX2
XFILL_1__10046_ vdd gnd FILL
XFILL_0__13564_ vdd gnd FILL
X_7710_ _7710_/A _7710_/B _7710_/C _7710_/Y vdd gnd OAI21X1
XFILL_0__8062_ vdd gnd FILL
XFILL_0__10776_ vdd gnd FILL
X_8690_ _8690_/A _8690_/Y vdd gnd INVX1
XFILL_0__12515_ vdd gnd FILL
XFILL_1__14854_ vdd gnd FILL
X_7641_ _7641_/A _7641_/B _7641_/Y vdd gnd NOR2X1
XFILL_2__11267_ vdd gnd FILL
XFILL_1__13805_ vdd gnd FILL
XFILL_1__14785_ vdd gnd FILL
XFILL_0__12446_ vdd gnd FILL
XFILL_1__11997_ vdd gnd FILL
X_7572_ _7572_/A _7572_/Y vdd gnd INVX1
XFILL_2__10218_ vdd gnd FILL
XFILL_1__13736_ vdd gnd FILL
XFILL_2__11198_ vdd gnd FILL
XFILL_1__10948_ vdd gnd FILL
X_9311_ _9311_/A _9311_/B _9311_/S _9311_/Y vdd gnd MUX2X1
XFILL_0__12377_ vdd gnd FILL
XFILL_0__8964_ vdd gnd FILL
XFILL_0__14116_ vdd gnd FILL
XFILL_1__13667_ vdd gnd FILL
XFILL_0__11328_ vdd gnd FILL
XFILL_1__10879_ vdd gnd FILL
X_9242_ _9242_/A _9242_/Y vdd gnd INVX1
XFILL_0__7915_ vdd gnd FILL
XFILL_1__12618_ vdd gnd FILL
XFILL_0__14047_ vdd gnd FILL
XFILL_1__13598_ vdd gnd FILL
XFILL_0__11259_ vdd gnd FILL
X_9173_ _9173_/A _9173_/B _9173_/C _9173_/Y vdd gnd AOI21X1
XFILL_0__7846_ vdd gnd FILL
XFILL_2__13908_ vdd gnd FILL
X_8124_ _8124_/A _8124_/B _8124_/C _8124_/Y vdd gnd OAI21X1
XFILL_0__7777_ vdd gnd FILL
XFILL_2__13839_ vdd gnd FILL
XFILL_0__9516_ vdd gnd FILL
X_8055_ _8055_/A _8055_/Y vdd gnd INVX1
XFILL_1__14219_ vdd gnd FILL
XFILL_1__8240_ vdd gnd FILL
XFILL_0__9447_ vdd gnd FILL
XFILL_1__8171_ vdd gnd FILL
XFILL_0__9378_ vdd gnd FILL
XFILL_1__7122_ vdd gnd FILL
XFILL_0__8329_ vdd gnd FILL
X_8957_ _8957_/A _8957_/B _8957_/Y vdd gnd NAND2X1
X_7908_ _7908_/A _7908_/B _7908_/C _7908_/Y vdd gnd OAI21X1
X_8888_ _8888_/D _8888_/CLK _8888_/Q vdd gnd DFFPOSX1
XFILL_1_CLKBUF1_insert31 vdd gnd FILL
X_7839_ _7839_/A _7839_/Y vdd gnd INVX1
XFILL_1_CLKBUF1_insert42 vdd gnd FILL
XFILL_1_CLKBUF1_insert53 vdd gnd FILL
XFILL_1_CLKBUF1_insert64 vdd gnd FILL
XFILL_1_CLKBUF1_insert75 vdd gnd FILL
XFILL_1_CLKBUF1_insert86 vdd gnd FILL
XFILL_1_CLKBUF1_insert97 vdd gnd FILL
X_11440_ _11440_/A _11440_/B _11440_/C _11440_/Y vdd gnd AOI21X1
X_9509_ _9509_/A _9509_/Y vdd gnd INVX1
XFILL257550x14550 vdd gnd FILL
X_11371_ _11371_/A _11371_/B _11371_/Y vdd gnd NAND2X1
XFILL_1__7886_ vdd gnd FILL
X_13110_ _13110_/A _13110_/B _13110_/C _13110_/Y vdd gnd NAND3X1
X_10322_ _10322_/A _10322_/B _10322_/C _10322_/D _10322_/Y vdd gnd AOI22X1
X_14090_ _14090_/A _14090_/Y vdd gnd INVX1
XFILL_1__9625_ vdd gnd FILL
X_13041_ _13041_/A _13041_/B _13041_/Y vdd gnd AND2X2
X_10253_ _10253_/A _10253_/B _10253_/Y vdd gnd NAND2X1
XFILL_1__9556_ vdd gnd FILL
XFILL_2__7300_ vdd gnd FILL
X_10184_ _10184_/A _10184_/B _10184_/Y vdd gnd AND2X2
XFILL_1__8507_ vdd gnd FILL
XFILL_1__9487_ vdd gnd FILL
XFILL_2__7231_ vdd gnd FILL
XFILL_1__8438_ vdd gnd FILL
X_13943_ _13943_/A _13943_/B _13943_/C _13943_/Y vdd gnd AOI21X1
XFILL_2__7162_ vdd gnd FILL
XFILL_1__8369_ vdd gnd FILL
X_13874_ _13874_/A _13874_/B _13874_/C _13874_/Y vdd gnd OAI21X1
XFILL_2__7093_ vdd gnd FILL
XFILL_0__10630_ vdd gnd FILL
X_12825_ _12825_/A _12825_/B _12825_/C _12825_/Y vdd gnd NOR3X1
XFILL_1__11920_ vdd gnd FILL
XFILL_2__12170_ vdd gnd FILL
XFILL_0__10561_ vdd gnd FILL
X_12756_ _12756_/A _12756_/B _12756_/Y vdd gnd NAND2X1
XFILL_0__12300_ vdd gnd FILL
XFILL_1__11851_ vdd gnd FILL
XFILL_0__13280_ vdd gnd FILL
XFILL_0__10492_ vdd gnd FILL
X_11707_ _11707_/A _11707_/Y vdd gnd INVX1
X_12687_ _12687_/A _12687_/B _12687_/Y vdd gnd NAND2X1
XFILL_1__10802_ vdd gnd FILL
XFILL_1__14570_ vdd gnd FILL
XFILL_0__12231_ vdd gnd FILL
XFILL_1__11782_ vdd gnd FILL
X_14426_ _14426_/A _14426_/B _14426_/Y vdd gnd NAND2X1
XFILL_2__10003_ vdd gnd FILL
X_11638_ _11638_/D _11638_/CLK _11638_/Q vdd gnd DFFPOSX1
XFILL_2__9734_ vdd gnd FILL
XFILL_1__13521_ vdd gnd FILL
XFILL_0__12162_ vdd gnd FILL
X_14357_ _14357_/A _14357_/B _14357_/C _14357_/Y vdd gnd OAI21X1
X_11569_ _11569_/A _11569_/B _11569_/C _11569_/Y vdd gnd OAI21X1
XFILL_2__9665_ vdd gnd FILL
XFILL_0__11113_ vdd gnd FILL
XFILL_1__10664_ vdd gnd FILL
XFILL_0__7700_ vdd gnd FILL
XFILL_0__12093_ vdd gnd FILL
X_13308_ _13308_/A _13308_/B _13308_/Y vdd gnd NOR2X1
X_14288_ _14288_/A _14288_/B _14288_/Y vdd gnd NAND2X1
XFILL_1__12403_ vdd gnd FILL
XFILL_0__8680_ vdd gnd FILL
XFILL_2__9596_ vdd gnd FILL
XFILL_1__13383_ vdd gnd FILL
XFILL_0__11044_ vdd gnd FILL
XFILL_1__10595_ vdd gnd FILL
XFILL_0__7631_ vdd gnd FILL
X_13239_ _13239_/A _13239_/B _13239_/C _13239_/Y vdd gnd OAI21X1
XFILL_1__12334_ vdd gnd FILL
XFILL_2__10905_ vdd gnd FILL
XFILL_0__7562_ vdd gnd FILL
XFILL_0__14803_ vdd gnd FILL
XFILL_1__12265_ vdd gnd FILL
XFILL_2__10836_ vdd gnd FILL
XFILL_0__9301_ vdd gnd FILL
XFILL_0__12995_ vdd gnd FILL
XFILL_0__7493_ vdd gnd FILL
XFILL_1__14004_ vdd gnd FILL
XFILL_2__7429_ vdd gnd FILL
XFILL_1__11216_ vdd gnd FILL
XFILL_0__14734_ vdd gnd FILL
XFILL_0__11946_ vdd gnd FILL
XFILL_1__12196_ vdd gnd FILL
XFILL_0__9232_ vdd gnd FILL
X_9860_ _9860_/A _9860_/B _9860_/C _9860_/Y vdd gnd OAI21X1
XFILL_2__12506_ vdd gnd FILL
XFILL_1__11147_ vdd gnd FILL
XFILL_0__14665_ vdd gnd FILL
XFILL_0__9163_ vdd gnd FILL
XFILL_0__11877_ vdd gnd FILL
X_8811_ _8811_/A _8811_/B _8811_/C _8811_/Y vdd gnd OAI21X1
X_9791_ _9791_/D _9791_/CLK _9791_/Q vdd gnd DFFPOSX1
XFILL_0__13616_ vdd gnd FILL
XFILL_2__12437_ vdd gnd FILL
XFILL_1__11078_ vdd gnd FILL
XFILL_0__10828_ vdd gnd FILL
XFILL_0__14596_ vdd gnd FILL
XFILL_0__8114_ vdd gnd FILL
XFILL_0__9094_ vdd gnd FILL
X_8742_ _8742_/A _8742_/B _8742_/C _8742_/Y vdd gnd OAI21X1
XFILL_1__10029_ vdd gnd FILL
XFILL_0__13547_ vdd gnd FILL
XFILL_0__8045_ vdd gnd FILL
X_8673_ _8673_/A _8673_/Y vdd gnd INVX1
XFILL_1__14837_ vdd gnd FILL
X_7624_ _7624_/A _7624_/Y vdd gnd INVX1
XFILL_0__12429_ vdd gnd FILL
XFILL_1__14768_ vdd gnd FILL
X_7555_ _7555_/A _7555_/B _7555_/C _7555_/Y vdd gnd AOI21X1
XFILL_0__9996_ vdd gnd FILL
XFILL_1__13719_ vdd gnd FILL
XFILL_1__14699_ vdd gnd FILL
XFILL_0__8947_ vdd gnd FILL
XFILL_1__7740_ vdd gnd FILL
X_7486_ _7486_/A _7486_/B _7486_/C _7486_/Y vdd gnd AOI21X1
X_9225_ _9225_/A _9225_/B _9225_/C _9225_/Y vdd gnd AOI21X1
XFILL_1__7671_ vdd gnd FILL
XFILL_1__9410_ vdd gnd FILL
X_9156_ _9156_/A _9156_/B _9156_/Y vdd gnd NAND2X1
XFILL_0__7829_ vdd gnd FILL
X_8107_ _8107_/A _8107_/B _8107_/Y vdd gnd NAND2X1
XFILL_1__9341_ vdd gnd FILL
X_9087_ _9087_/A _9087_/B _9087_/C _9087_/Y vdd gnd OAI21X1
X_8038_ _8038_/A _8038_/Y vdd gnd INVX1
XFILL_1__9272_ vdd gnd FILL
XFILL_1__8223_ vdd gnd FILL
X_10940_ _10940_/A _10940_/B _10940_/C _10940_/D _10940_/Y vdd gnd AOI22X1
XFILL_1__8154_ vdd gnd FILL
X_9989_ _9989_/A _9989_/Y vdd gnd INVX1
XFILL_1__7105_ vdd gnd FILL
XFILL_1__8085_ vdd gnd FILL
X_10871_ _10871_/A _10871_/Y vdd gnd INVX1
X_12610_ _12610_/D _12610_/CLK _12610_/Q vdd gnd DFFPOSX1
X_13590_ _13590_/A _13590_/B _13590_/Y vdd gnd NAND2X1
X_12541_ _12541_/D _12541_/CLK _12541_/Q vdd gnd DFFPOSX1
X_12472_ _12472_/A _12472_/B _12472_/Y vdd gnd NAND2X1
XFILL_1__8987_ vdd gnd FILL
X_14211_ _14211_/D _14211_/CLK _14211_/Q vdd gnd DFFPOSX1
X_11423_ _11423_/A _11423_/B _11423_/C _11423_/Y vdd gnd OAI21X1
X_11354_ _11354_/A _11354_/B _11354_/C _11354_/Y vdd gnd NAND3X1
X_14142_ _14142_/A _14142_/B _14142_/C _14142_/Y vdd gnd OAI21X1
XFILL_2__9450_ vdd gnd FILL
XFILL_1__7869_ vdd gnd FILL
X_10305_ _10305_/A _10305_/B _10305_/C _10305_/Y vdd gnd OAI21X1
XFILL_1__9608_ vdd gnd FILL
X_14073_ _14073_/A _14073_/B _14073_/C _14073_/Y vdd gnd OAI21X1
X_11285_ _11285_/A _11285_/B _11285_/Y vdd gnd NOR2X1
XCLKBUF1_insert107 CLKBUF1_insert107/A CLKBUF1_insert107/Y vdd gnd CLKBUF1
XFILL_2__9381_ vdd gnd FILL
XFILL_1__10380_ vdd gnd FILL
X_13024_ _13024_/A _13024_/B _13024_/Y vdd gnd NAND2X1
X_10236_ _10236_/A _10236_/B _10236_/Y vdd gnd NAND2X1
XFILL_1__9539_ vdd gnd FILL
X_10167_ _10167_/A _10167_/B _10167_/C _10167_/Y vdd gnd OAI21X1
XFILL_1__12050_ vdd gnd FILL
XFILL_0__11800_ vdd gnd FILL
XFILL_0__12780_ vdd gnd FILL
XFILL_1__11001_ vdd gnd FILL
X_10098_ _10098_/A _10098_/B _10098_/C _10098_/Y vdd gnd OAI21X1
XFILL_0__11731_ vdd gnd FILL
X_13926_ _13926_/A _13926_/B _13926_/S _13926_/Y vdd gnd MUX2X1
XFILL_0__14450_ vdd gnd FILL
XFILL_2__12222_ vdd gnd FILL
X_13857_ _13857_/A _13857_/B _13857_/Y vdd gnd NAND2X1
XFILL_2__7076_ vdd gnd FILL
XFILL_0__13401_ vdd gnd FILL
XFILL_0__10613_ vdd gnd FILL
XFILL_1__12952_ vdd gnd FILL
XFILL_0__14381_ vdd gnd FILL
XFILL_1_BUFX2_insert240 vdd gnd FILL
XFILL_0__11593_ vdd gnd FILL
X_12808_ _12808_/A _12808_/B _12808_/C _12808_/Y vdd gnd NAND3X1
XFILL_1_BUFX2_insert251 vdd gnd FILL
XFILL_1_BUFX2_insert262 vdd gnd FILL
XFILL_2__12153_ vdd gnd FILL
X_13788_ _13788_/A _13788_/B _13788_/C _13788_/Y vdd gnd NAND3X1
XFILL_1__11903_ vdd gnd FILL
XFILL_0__13332_ vdd gnd FILL
XFILL_1_BUFX2_insert273 vdd gnd FILL
XFILL_0__10544_ vdd gnd FILL
XCLKBUF1_insert33 CLKBUF1_insert33/A CLKBUF1_insert33/Y vdd gnd CLKBUF1
XFILL_1__12883_ vdd gnd FILL
XFILL_1_BUFX2_insert284 vdd gnd FILL
XCLKBUF1_insert44 CLKBUF1_insert44/A CLKBUF1_insert44/Y vdd gnd CLKBUF1
XFILL_1_BUFX2_insert295 vdd gnd FILL
X_12739_ _12739_/A _12739_/B _12739_/C _12739_/Y vdd gnd AOI21X1
XCLKBUF1_insert55 CLKBUF1_insert55/A CLKBUF1_insert55/Y vdd gnd CLKBUF1
XCLKBUF1_insert66 CLKBUF1_insert66/A CLKBUF1_insert66/Y vdd gnd CLKBUF1
XFILL_1__14622_ vdd gnd FILL
XFILL_1__11834_ vdd gnd FILL
XFILL_2__12084_ vdd gnd FILL
XCLKBUF1_insert77 CLKBUF1_insert77/A CLKBUF1_insert77/Y vdd gnd CLKBUF1
XFILL_0__13263_ vdd gnd FILL
XFILL_0__10475_ vdd gnd FILL
XCLKBUF1_insert88 CLKBUF1_insert88/A CLKBUF1_insert88/Y vdd gnd CLKBUF1
XFILL_0__9850_ vdd gnd FILL
XCLKBUF1_insert99 CLKBUF1_insert99/A CLKBUF1_insert99/Y vdd gnd CLKBUF1
XFILL_0__12214_ vdd gnd FILL
XFILL_1__11765_ vdd gnd FILL
XFILL_0__13194_ vdd gnd FILL
X_14409_ _14409_/A _14409_/B _14409_/C _14409_/Y vdd gnd AOI21X1
XFILL_0__8801_ vdd gnd FILL
X_7340_ _7340_/A _7340_/B _7340_/Y vdd gnd NAND2X1
XFILL_2__9717_ vdd gnd FILL
XFILL_1__13504_ vdd gnd FILL
XFILL_1__14484_ vdd gnd FILL
XFILL_0__12145_ vdd gnd FILL
XFILL_1__11696_ vdd gnd FILL
XFILL_0__8732_ vdd gnd FILL
X_7271_ _7271_/A _7271_/B _7271_/C _7271_/Y vdd gnd NAND3X1
XFILL_2__9648_ vdd gnd FILL
XFILL_1__10647_ vdd gnd FILL
X_9010_ _9010_/A _9010_/B _9010_/S _9010_/Y vdd gnd MUX2X1
XFILL_2__12986_ vdd gnd FILL
XFILL_0__12076_ vdd gnd FILL
XFILL_0__8663_ vdd gnd FILL
XFILL_0__11027_ vdd gnd FILL
XFILL_2__9579_ vdd gnd FILL
XFILL_1__13366_ vdd gnd FILL
XFILL_1__10578_ vdd gnd FILL
XFILL_0__7614_ vdd gnd FILL
XFILL_0__8594_ vdd gnd FILL
XFILL_1__12317_ vdd gnd FILL
XFILL_1__13297_ vdd gnd FILL
XFILL_0__7545_ vdd gnd FILL
XFILL_1__12248_ vdd gnd FILL
XFILL_2__10819_ vdd gnd FILL
XFILL_0__12978_ vdd gnd FILL
X_9912_ _9912_/A _9912_/B _9912_/S _9912_/Y vdd gnd MUX2X1
XFILL_0__7476_ vdd gnd FILL
XFILL_0__14717_ vdd gnd FILL
XFILL_0__11929_ vdd gnd FILL
XFILL_1__12179_ vdd gnd FILL
XFILL_0__9215_ vdd gnd FILL
X_9843_ _9843_/D _9843_/CLK _9843_/Q vdd gnd DFFPOSX1
XFILL_0__14648_ vdd gnd FILL
XFILL_0__9146_ vdd gnd FILL
X_9774_ _9774_/D _9774_/CLK _9774_/Q vdd gnd DFFPOSX1
XFILL_0__14579_ vdd gnd FILL
XFILL_0__9077_ vdd gnd FILL
X_8725_ _8725_/A _8725_/B _8725_/C _8725_/Y vdd gnd OAI21X1
XFILL_0__8028_ vdd gnd FILL
X_8656_ _8656_/A _8656_/B _8656_/Y vdd gnd NOR2X1
XFILL_1__9890_ vdd gnd FILL
X_7607_ _7607_/A _7607_/B _7607_/C _7607_/Y vdd gnd OAI21X1
X_8587_ _8587_/A _8587_/B _8587_/C _8587_/Y vdd gnd OAI21X1
X_7538_ _7538_/A _7538_/B _7538_/C _7538_/Y vdd gnd OAI21X1
XFILL_0__9979_ vdd gnd FILL
XFILL_1__8772_ vdd gnd FILL
XFILL_1__7723_ vdd gnd FILL
X_7469_ _7469_/A _7469_/B _7469_/C _7469_/Y vdd gnd OAI21X1
X_9208_ _9208_/A _9208_/Y vdd gnd INVX1
XFILL_1__7654_ vdd gnd FILL
X_11070_ _11070_/A _11070_/B _11070_/C _11070_/Y vdd gnd NAND3X1
X_9139_ _9139_/A _9139_/B _9139_/C _9139_/Y vdd gnd NAND3X1
XFILL_1__7585_ vdd gnd FILL
X_10021_ _10021_/A _10021_/B _10021_/C _10021_/Y vdd gnd OAI21X1
XFILL_1__9324_ vdd gnd FILL
XFILL_1__9255_ vdd gnd FILL
XFILL257550x165750 vdd gnd FILL
X_14760_ _14760_/A _14760_/B _14760_/C _14760_/Y vdd gnd OAI21X1
XFILL_1__8206_ vdd gnd FILL
X_11972_ _11972_/A _11972_/B _11972_/C _11972_/Y vdd gnd OAI21X1
XFILL_1__9186_ vdd gnd FILL
X_13711_ _13711_/A _13711_/B _13711_/C _13711_/Y vdd gnd OAI21X1
XFILL257250x36150 vdd gnd FILL
X_10923_ _10923_/A _10923_/B _10923_/C _10923_/Y vdd gnd AOI21X1
X_14691_ _14691_/A _14691_/B _14691_/C _14691_/Y vdd gnd AOI21X1
XFILL_1__8137_ vdd gnd FILL
X_13642_ _13642_/A _13642_/Y vdd gnd INVX2
X_10854_ _10854_/A _10854_/B _10854_/Y vdd gnd NAND2X1
XFILL_2__8950_ vdd gnd FILL
XFILL_1__8068_ vdd gnd FILL
XFILL_2__7901_ vdd gnd FILL
XFILL_0_BUFX2_insert203 vdd gnd FILL
X_13573_ _13573_/A _13573_/B _13573_/Y vdd gnd NOR2X1
XFILL_0_BUFX2_insert214 vdd gnd FILL
X_10785_ _10785_/A _10785_/B _10785_/C _10785_/Y vdd gnd AOI21X1
XFILL_0_BUFX2_insert225 vdd gnd FILL
XFILL_0_BUFX2_insert236 vdd gnd FILL
X_12524_ _12524_/A _12524_/B _12524_/Y vdd gnd NAND2X1
XFILL_0_BUFX2_insert247 vdd gnd FILL
XFILL_2__7832_ vdd gnd FILL
XFILL_0_BUFX2_insert258 vdd gnd FILL
XFILL_0_BUFX2_insert269 vdd gnd FILL
XFILL_0__10260_ vdd gnd FILL
X_12455_ _12455_/A _12455_/B _12455_/Y vdd gnd NAND2X1
XFILL_2__7763_ vdd gnd FILL
XFILL_1__11550_ vdd gnd FILL
XFILL_0__10191_ vdd gnd FILL
X_11406_ _11406_/A _11406_/B _11406_/C _11406_/Y vdd gnd OAI21X1
XFILL_1__10501_ vdd gnd FILL
X_12386_ _12386_/A _12386_/Y vdd gnd INVX1
XFILL_2__7694_ vdd gnd FILL
XFILL_1__11481_ vdd gnd FILL
X_14125_ _14125_/A _14125_/B _14125_/C _14125_/Y vdd gnd OAI21X1
X_11337_ _11337_/A _11337_/B _11337_/Y vdd gnd NOR2X1
XFILL_1__13220_ vdd gnd FILL
XFILL_1__10432_ vdd gnd FILL
XFILL_0__13950_ vdd gnd FILL
X_14056_ _14056_/A _14056_/B _14056_/C _14056_/Y vdd gnd OAI21X1
X_11268_ _11268_/A _11268_/Y vdd gnd INVX1
XFILL_1__13151_ vdd gnd FILL
XFILL_2__11722_ vdd gnd FILL
XFILL_0__12901_ vdd gnd FILL
XFILL_1__10363_ vdd gnd FILL
XFILL_0__13881_ vdd gnd FILL
X_13007_ _13007_/A _13007_/B _13007_/Y vdd gnd NAND2X1
X_10219_ _10219_/A _10219_/B _10219_/S _10219_/Y vdd gnd MUX2X1
XFILL_2__8315_ vdd gnd FILL
XFILL_1__12102_ vdd gnd FILL
X_11199_ _11199_/A _11199_/B _11199_/Y vdd gnd NOR2X1
XFILL_1__13082_ vdd gnd FILL
XFILL_2__9295_ vdd gnd FILL
XFILL_0__12832_ vdd gnd FILL
XFILL_1__10294_ vdd gnd FILL
XFILL_0__7330_ vdd gnd FILL
XFILL_2__10604_ vdd gnd FILL
XFILL_1__12033_ vdd gnd FILL
XFILL_2__8246_ vdd gnd FILL
XFILL_2__11584_ vdd gnd FILL
XFILL_0__12763_ vdd gnd FILL
XFILL_0__7261_ vdd gnd FILL
XFILL_2__10535_ vdd gnd FILL
XFILL_0__11714_ vdd gnd FILL
XFILL_0__9000_ vdd gnd FILL
X_13909_ _13909_/A _13909_/B _13909_/C _13909_/Y vdd gnd AOI21X1
XFILL_0__12694_ vdd gnd FILL
XFILL_0__7192_ vdd gnd FILL
X_14889_ _14889_/D _14889_/CLK _14889_/Q vdd gnd DFFPOSX1
XFILL_0__14433_ vdd gnd FILL
XFILL_1__13984_ vdd gnd FILL
XFILL_2__12205_ vdd gnd FILL
XFILL_1__12935_ vdd gnd FILL
XFILL_0__14364_ vdd gnd FILL
X_8510_ _8510_/A _8510_/B _8510_/Y vdd gnd NOR2X1
XFILL_0__11576_ vdd gnd FILL
X_9490_ _9490_/A _9490_/B _9490_/C _9490_/Y vdd gnd OAI21X1
XFILL_2__12136_ vdd gnd FILL
XFILL_0__13315_ vdd gnd FILL
XFILL_0__10527_ vdd gnd FILL
XFILL_0__9902_ vdd gnd FILL
XFILL_0__14295_ vdd gnd FILL
XFILL_1__12866_ vdd gnd FILL
X_8441_ _8441_/A _8441_/B _8441_/Y vdd gnd OR2X2
XFILL_1__14605_ vdd gnd FILL
XFILL_2__12067_ vdd gnd FILL
XFILL_1__11817_ vdd gnd FILL
XFILL_0__13246_ vdd gnd FILL
XFILL_0__10458_ vdd gnd FILL
XFILL_1__12797_ vdd gnd FILL
X_8372_ _8372_/A _8372_/B _8372_/Y vdd gnd NAND2X1
XFILL257550x230550 vdd gnd FILL
XFILL_0__13177_ vdd gnd FILL
XFILL_1__11748_ vdd gnd FILL
XFILL_0__10389_ vdd gnd FILL
X_7323_ _7323_/A _7323_/B _7323_/Y vdd gnd AND2X2
XFILL_0__12128_ vdd gnd FILL
XFILL_1__14467_ vdd gnd FILL
XFILL_0__8715_ vdd gnd FILL
X_7254_ _7254_/A _7254_/B _7254_/C _7254_/Y vdd gnd AOI21X1
XFILL_0__9695_ vdd gnd FILL
XFILL_1__13418_ vdd gnd FILL
XFILL_2__12969_ vdd gnd FILL
XFILL_0__12059_ vdd gnd FILL
XFILL_1__14398_ vdd gnd FILL
XFILL_0__8646_ vdd gnd FILL
X_7185_ _7185_/A _7185_/B _7185_/S _7185_/Y vdd gnd MUX2X1
XFILL_2__14708_ vdd gnd FILL
XFILL_1__13349_ vdd gnd FILL
XFILL_1__7370_ vdd gnd FILL
XFILL_0__8577_ vdd gnd FILL
XFILL_2__14639_ vdd gnd FILL
XFILL_0__7528_ vdd gnd FILL
XFILL_1_BUFX2_insert4 vdd gnd FILL
XFILL_1__9040_ vdd gnd FILL
XFILL_0__7459_ vdd gnd FILL
X_9826_ _9826_/D _9826_/CLK _9826_/Q vdd gnd DFFPOSX1
XFILL_0__9129_ vdd gnd FILL
X_9757_ _9757_/A _9757_/B _9757_/C _9757_/Y vdd gnd OAI21X1
XBUFX2_insert308 BUFX2_insert308/A BUFX2_insert308/Y vdd gnd BUFX2
XFILL_1__9942_ vdd gnd FILL
X_8708_ _8708_/A _8708_/B _8708_/Y vdd gnd NAND2X1
XBUFX2_insert319 BUFX2_insert319/A BUFX2_insert319/Y vdd gnd BUFX2
X_9688_ _9688_/A _9688_/B _9688_/Y vdd gnd OR2X2
X_10570_ _10570_/A _10570_/Y vdd gnd INVX1
XFILL_1__9873_ vdd gnd FILL
X_8639_ _8639_/A _8639_/B _8639_/Y vdd gnd NAND2X1
XFILL_1__8824_ vdd gnd FILL
XFILL257550x140550 vdd gnd FILL
X_12240_ _12240_/A _12240_/B _12240_/Y vdd gnd NOR2X1
XFILL_1__8755_ vdd gnd FILL
X_12171_ _12171_/A _12171_/Y vdd gnd INVX1
XFILL_1__7706_ vdd gnd FILL
XFILL_1__8686_ vdd gnd FILL
X_11122_ _11122_/A _11122_/B _11122_/Y vdd gnd NAND2X1
XFILL_1__7637_ vdd gnd FILL
X_11053_ _11053_/A _11053_/B _11053_/C _11053_/Y vdd gnd OAI21X1
XFILL_1__7568_ vdd gnd FILL
X_10004_ _10004_/A _10004_/Y vdd gnd INVX2
XFILL_1__9307_ vdd gnd FILL
XFILL_2__8100_ vdd gnd FILL
XFILL_1__7499_ vdd gnd FILL
X_14812_ _14812_/A _14812_/B _14812_/Y vdd gnd NOR2X1
XFILL_1__9238_ vdd gnd FILL
XFILL_2__8031_ vdd gnd FILL
X_14743_ _14743_/A _14743_/B _14743_/Y vdd gnd OR2X2
XFILL_2__10320_ vdd gnd FILL
X_11955_ _11955_/A _11955_/Y vdd gnd INVX1
XFILL_1__9169_ vdd gnd FILL
X_10906_ _10906_/A _10906_/B _10906_/S _10906_/Y vdd gnd MUX2X1
X_14674_ _14674_/A _14674_/B _14674_/Y vdd gnd OR2X2
XFILL_2__10251_ vdd gnd FILL
X_11886_ _11886_/A _11886_/Y vdd gnd INVX2
XFILL_0__11430_ vdd gnd FILL
XFILL_1__10981_ vdd gnd FILL
X_13625_ _13625_/A _13625_/B _13625_/S _13625_/Y vdd gnd MUX2X1
X_10837_ _10837_/A _10837_/Y vdd gnd INVX1
XFILL_2__8933_ vdd gnd FILL
XFILL_1__12720_ vdd gnd FILL
XFILL_2__10182_ vdd gnd FILL
XFILL_0__11361_ vdd gnd FILL
X_13556_ _13556_/A _13556_/B _13556_/Y vdd gnd NAND2X1
XFILL_0__13100_ vdd gnd FILL
X_10768_ _10768_/A _10768_/Y vdd gnd INVX1
XFILL_1__12651_ vdd gnd FILL
XFILL_0__10312_ vdd gnd FILL
XFILL_0__14080_ vdd gnd FILL
X_12507_ _12507_/A _12507_/B _12507_/C _12507_/Y vdd gnd OAI21X1
XFILL_0__11292_ vdd gnd FILL
XFILL_2__7815_ vdd gnd FILL
X_13487_ _13487_/D _13487_/CLK _13487_/Q vdd gnd DFFPOSX1
X_10699_ _10699_/D _10699_/CLK _10699_/Q vdd gnd DFFPOSX1
XFILL_1__11602_ vdd gnd FILL
XFILL_0__13031_ vdd gnd FILL
XFILL_0__10243_ vdd gnd FILL
X_12438_ _12438_/A _12438_/B _12438_/C _12438_/Y vdd gnd OAI21X1
XFILL_2__7746_ vdd gnd FILL
XFILL_1__14321_ vdd gnd FILL
XFILL_1__11533_ vdd gnd FILL
XFILL_0__10174_ vdd gnd FILL
X_12369_ _12369_/A _12369_/Y vdd gnd INVX1
XFILL_2__7677_ vdd gnd FILL
XFILL_1__14252_ vdd gnd FILL
XFILL_1__11464_ vdd gnd FILL
XFILL_0__8500_ vdd gnd FILL
X_14108_ _14108_/A _14108_/B _14108_/C _14108_/Y vdd gnd OAI21X1
XFILL_0__9480_ vdd gnd FILL
XFILL_1__13203_ vdd gnd FILL
XFILL_1__10415_ vdd gnd FILL
XFILL_0__13933_ vdd gnd FILL
XFILL_1__11395_ vdd gnd FILL
XFILL_0__8431_ vdd gnd FILL
X_14039_ _14039_/A _14039_/B _14039_/C _14039_/Y vdd gnd OAI21X1
XFILL_1__13134_ vdd gnd FILL
XFILL_2__11705_ vdd gnd FILL
XFILL_1__10346_ vdd gnd FILL
XFILL_0__13864_ vdd gnd FILL
XFILL_0__8362_ vdd gnd FILL
X_8990_ _8990_/A _8990_/B _8990_/Y vdd gnd NAND2X1
XFILL_1__13065_ vdd gnd FILL
XFILL_1__10277_ vdd gnd FILL
XFILL_0__12815_ vdd gnd FILL
XFILL_0__7313_ vdd gnd FILL
XFILL_0__13795_ vdd gnd FILL
X_7941_ _7941_/D _7941_/CLK _7941_/Q vdd gnd DFFPOSX1
XFILL_0__8293_ vdd gnd FILL
XFILL_1__12016_ vdd gnd FILL
XFILL_2__8229_ vdd gnd FILL
XFILL_0__12746_ vdd gnd FILL
XFILL_0__7244_ vdd gnd FILL
X_7872_ _7872_/A _7872_/B _7872_/C _7872_/Y vdd gnd OAI21X1
XFILL_2__10518_ vdd gnd FILL
XFILL_0__12677_ vdd gnd FILL
XFILL_0__7175_ vdd gnd FILL
X_9611_ _9611_/A _9611_/Y vdd gnd INVX1
XFILL_2__10449_ vdd gnd FILL
XFILL_0__14416_ vdd gnd FILL
XFILL_1__13967_ vdd gnd FILL
X_9542_ _9542_/A _9542_/Y vdd gnd INVX1
XFILL_0__14347_ vdd gnd FILL
XFILL_1__12918_ vdd gnd FILL
XFILL_0__11559_ vdd gnd FILL
XFILL_1__13898_ vdd gnd FILL
X_9473_ _9473_/A _9473_/B _9473_/C _9473_/Y vdd gnd OAI21X1
XFILL_0__14278_ vdd gnd FILL
XFILL_1__12849_ vdd gnd FILL
X_8424_ _8424_/A _8424_/B _8424_/C _8424_/Y vdd gnd NAND3X1
XFILL_0__13229_ vdd gnd FILL
X_8355_ _8355_/A _8355_/B _8355_/C _8355_/Y vdd gnd OAI21X1
X_7306_ _7306_/A _7306_/Y vdd gnd INVX1
XFILL_0__9747_ vdd gnd FILL
XFILL_1__8540_ vdd gnd FILL
X_8286_ _8286_/A _8286_/B _8286_/C _8286_/Y vdd gnd NAND3X1
X_7237_ _7237_/A _7237_/Y vdd gnd INVX1
XFILL_0__9678_ vdd gnd FILL
XFILL_1__8471_ vdd gnd FILL
XFILL_1__7422_ vdd gnd FILL
XFILL_0__8629_ vdd gnd FILL
X_7168_ _7168_/A _7168_/B _7168_/C _7168_/Y vdd gnd NAND3X1
XFILL_1__7353_ vdd gnd FILL
X_7099_ _7099_/A _7099_/Y vdd gnd INVX1
XFILL_2_BUFX2_insert117 vdd gnd FILL
XFILL_2_BUFX2_insert139 vdd gnd FILL
XFILL_1__7284_ vdd gnd FILL
XFILL_1__9023_ vdd gnd FILL
X_11740_ _11740_/A _11740_/B _11740_/C _11740_/Y vdd gnd OAI21X1
X_9809_ _9809_/D _9809_/CLK _9809_/Q vdd gnd DFFPOSX1
X_11671_ _11671_/D _11671_/CLK _11671_/Q vdd gnd DFFPOSX1
XBUFX2_insert116 BUFX2_insert116/A BUFX2_insert116/Y vdd gnd BUFX2
XBUFX2_insert127 BUFX2_insert127/A BUFX2_insert127/Y vdd gnd BUFX2
X_13410_ _13410_/A _13410_/B _13410_/C _13410_/Y vdd gnd OAI21X1
X_10622_ _10622_/A _10622_/B _10622_/C _10622_/Y vdd gnd OAI21X1
XBUFX2_insert138 BUFX2_insert138/A BUFX2_insert138/Y vdd gnd BUFX2
XFILL_1__9925_ vdd gnd FILL
X_14390_ _14390_/A _14390_/B _14390_/C _14390_/Y vdd gnd NAND3X1
XBUFX2_insert149 BUFX2_insert149/A BUFX2_insert149/Y vdd gnd BUFX2
X_13341_ _13341_/A _13341_/B _13341_/Y vdd gnd NAND2X1
X_10553_ _10553_/A _10553_/Y vdd gnd INVX1
XFILL_1__9856_ vdd gnd FILL
XFILL_1__8807_ vdd gnd FILL
X_13272_ _13272_/A _13272_/B _13272_/C _13272_/Y vdd gnd AOI21X1
X_10484_ _10484_/A _10484_/B _10484_/S _10484_/Y vdd gnd MUX2X1
X_12223_ _12223_/A _12223_/Y vdd gnd INVX1
XFILL_1__8738_ vdd gnd FILL
X_12154_ _12154_/A _12154_/B _12154_/Y vdd gnd NAND2X1
XFILL_1__8669_ vdd gnd FILL
X_11105_ _11105_/A _11105_/B _11105_/C _11105_/Y vdd gnd AOI21X1
XFILL_1__10200_ vdd gnd FILL
X_12085_ _12085_/A _12085_/B _12085_/Y vdd gnd NAND2X1
XFILL_2__7393_ vdd gnd FILL
XFILL_1__11180_ vdd gnd FILL
XFILL_0__10930_ vdd gnd FILL
X_11036_ _11036_/A _11036_/B _11036_/Y vdd gnd NAND2X1
XFILL_1__10131_ vdd gnd FILL
XFILL_2__12470_ vdd gnd FILL
XFILL_0__10861_ vdd gnd FILL
XFILL_1__10062_ vdd gnd FILL
XFILL_0__13580_ vdd gnd FILL
XFILL_0__10792_ vdd gnd FILL
XFILL_2__8014_ vdd gnd FILL
XFILL_2__14140_ vdd gnd FILL
X_12987_ _12987_/A _12987_/B _12987_/Y vdd gnd NOR2X1
XFILL_0__12531_ vdd gnd FILL
X_14726_ _14726_/A _14726_/B _14726_/Y vdd gnd AND2X2
X_11938_ _11938_/A _11938_/B _11938_/C _11938_/Y vdd gnd AOI21X1
XFILL_2__10303_ vdd gnd FILL
XFILL_1__13821_ vdd gnd FILL
XFILL_0__12462_ vdd gnd FILL
X_14657_ _14657_/A _14657_/Y vdd gnd INVX1
XFILL_2__10234_ vdd gnd FILL
X_11869_ _11869_/A _11869_/B _11869_/C _11869_/Y vdd gnd OAI21X1
XFILL_2__13022_ vdd gnd FILL
XFILL_0__11413_ vdd gnd FILL
XFILL_1__13752_ vdd gnd FILL
XFILL_1__10964_ vdd gnd FILL
XFILL_0__12393_ vdd gnd FILL
X_13608_ _13608_/A _13608_/B _13608_/S _13608_/Y vdd gnd MUX2X1
XFILL_0__8980_ vdd gnd FILL
X_14588_ _14588_/A _14588_/Y vdd gnd INVX1
XFILL_2__10165_ vdd gnd FILL
XFILL_1__12703_ vdd gnd FILL
XFILL_0__14132_ vdd gnd FILL
XFILL_0__11344_ vdd gnd FILL
XFILL_1__10895_ vdd gnd FILL
XFILL_1__13683_ vdd gnd FILL
X_13539_ _13539_/A _13539_/B _13539_/C _13539_/Y vdd gnd OAI21X1
XFILL_1__12634_ vdd gnd FILL
XFILL_2__10096_ vdd gnd FILL
XFILL_0__14063_ vdd gnd FILL
XFILL_0__11275_ vdd gnd FILL
XFILL_0__7862_ vdd gnd FILL
XFILL_0__13014_ vdd gnd FILL
XFILL_0__10226_ vdd gnd FILL
XFILL_0__9601_ vdd gnd FILL
X_8140_ _8140_/A _8140_/B _8140_/Y vdd gnd NAND2X1
XFILL_2__7729_ vdd gnd FILL
XFILL_0__7793_ vdd gnd FILL
XFILL_1__14304_ vdd gnd FILL
XFILL_1__11516_ vdd gnd FILL
XFILL_0__10157_ vdd gnd FILL
XFILL_1__12496_ vdd gnd FILL
XFILL_0__9532_ vdd gnd FILL
X_8071_ _8071_/A _8071_/B _8071_/S _8071_/Y vdd gnd MUX2X1
XFILL_1__14235_ vdd gnd FILL
XFILL_1__11447_ vdd gnd FILL
XFILL_2__10998_ vdd gnd FILL
XFILL_0__10088_ vdd gnd FILL
XFILL_0__9463_ vdd gnd FILL
XFILL_0__13916_ vdd gnd FILL
XFILL_1__11378_ vdd gnd FILL
XFILL_0__8414_ vdd gnd FILL
XFILL_0__9394_ vdd gnd FILL
XFILL_1__13117_ vdd gnd FILL
XFILL_1__10329_ vdd gnd FILL
XFILL_1__14097_ vdd gnd FILL
XFILL_0__13847_ vdd gnd FILL
XFILL_0__8345_ vdd gnd FILL
XFILL_1__13048_ vdd gnd FILL
X_8973_ _8973_/A _8973_/B _8973_/C _8973_/Y vdd gnd OAI21X1
XFILL_0__13778_ vdd gnd FILL
X_7924_ _7924_/D _7924_/CLK _7924_/Q vdd gnd DFFPOSX1
XFILL_0__8276_ vdd gnd FILL
XFILL_0__12729_ vdd gnd FILL
XFILL_0__7227_ vdd gnd FILL
X_7855_ _7855_/A _7855_/B _7855_/C _7855_/Y vdd gnd OAI21X1
XFILL_0__7158_ vdd gnd FILL
X_7786_ _7786_/A _7786_/B _7786_/Y vdd gnd NAND2X1
X_9525_ _9525_/A _9525_/B _9525_/C _9525_/Y vdd gnd AOI21X1
XFILL_0__7089_ vdd gnd FILL
XFILL_1__9710_ vdd gnd FILL
X_9456_ _9456_/A _9456_/B _9456_/Y vdd gnd NAND2X1
XFILL_1__9641_ vdd gnd FILL
X_8407_ _8407_/A _8407_/B _8407_/C _8407_/Y vdd gnd AOI21X1
X_9387_ _9387_/A _9387_/B _9387_/Y vdd gnd OR2X2
XFILL_1__9572_ vdd gnd FILL
X_8338_ _8338_/A _8338_/B _8338_/C _8338_/Y vdd gnd OAI21X1
XFILL_1__8523_ vdd gnd FILL
X_8269_ _8269_/A _8269_/B _8269_/C _8269_/Y vdd gnd OAI21X1
XFILL_1__8454_ vdd gnd FILL
XFILL_1__7405_ vdd gnd FILL
XFILL_1__8385_ vdd gnd FILL
X_12910_ _12910_/A _12910_/B _12910_/Y vdd gnd AND2X2
X_13890_ _13890_/A _13890_/B _13890_/C _13890_/Y vdd gnd OAI21X1
XFILL_1__7336_ vdd gnd FILL
X_12841_ _12841_/A _12841_/B _12841_/C _12841_/Y vdd gnd OAI21X1
XFILL_1__7267_ vdd gnd FILL
XFILL_1__9006_ vdd gnd FILL
X_12772_ _12772_/A _12772_/Y vdd gnd INVX1
XFILL_1__7198_ vdd gnd FILL
X_14511_ _14511_/D _14511_/CLK _14511_/Q vdd gnd DFFPOSX1
X_11723_ _11723_/A _11723_/B _11723_/C _11723_/D _11723_/Y vdd gnd AOI22X1
X_14442_ _14442_/A _14442_/B _14442_/Y vdd gnd NAND2X1
X_11654_ _11654_/D _11654_/CLK _11654_/Q vdd gnd DFFPOSX1
X_10605_ _10605_/A _10605_/B _10605_/Y vdd gnd NAND2X1
X_14373_ _14373_/A _14373_/B _14373_/Y vdd gnd AND2X2
XFILL_2__8701_ vdd gnd FILL
XFILL_1__9908_ vdd gnd FILL
X_11585_ _11585_/A _11585_/B _11585_/C _11585_/Y vdd gnd OAI21X1
XFILL_1__10680_ vdd gnd FILL
X_13324_ _13324_/A _13324_/B _13324_/C _13324_/Y vdd gnd NAND3X1
X_10536_ _10536_/A _10536_/B _10536_/Y vdd gnd NAND2X1
XFILL_2__8632_ vdd gnd FILL
XFILL_0__11060_ vdd gnd FILL
X_13255_ _13255_/A _13255_/B _13255_/C _13255_/Y vdd gnd OAI21X1
X_10467_ _10467_/A _10467_/B _10467_/Y vdd gnd NOR2X1
XFILL_0__10011_ vdd gnd FILL
XFILL_2__8563_ vdd gnd FILL
XFILL_1__12350_ vdd gnd FILL
X_12206_ _12206_/A _12206_/B _12206_/Y vdd gnd NOR2X1
X_13186_ _13186_/A _13186_/B _13186_/Y vdd gnd NAND2X1
XFILL_1__11301_ vdd gnd FILL
X_10398_ _10398_/A _10398_/Y vdd gnd INVX1
XFILL_1__12281_ vdd gnd FILL
X_12137_ _12137_/A _12137_/B _12137_/Y vdd gnd OR2X2
XFILL_1__11232_ vdd gnd FILL
XFILL_1__14020_ vdd gnd FILL
XFILL_0__14750_ vdd gnd FILL
XFILL_0__11962_ vdd gnd FILL
X_12068_ _12068_/A _12068_/B _12068_/Y vdd gnd NAND2X1
XFILL_2__12522_ vdd gnd FILL
XFILL_1__11163_ vdd gnd FILL
XFILL_0__10913_ vdd gnd FILL
XFILL_0__13701_ vdd gnd FILL
X_11019_ _11019_/A _11019_/B _11019_/Y vdd gnd AND2X2
XFILL_0__14681_ vdd gnd FILL
XFILL_0__11893_ vdd gnd FILL
XFILL_1__10114_ vdd gnd FILL
XFILL_2__12453_ vdd gnd FILL
XFILL_0__13632_ vdd gnd FILL
XFILL_1__11094_ vdd gnd FILL
XFILL_0__10844_ vdd gnd FILL
XFILL_0__8130_ vdd gnd FILL
XFILL256350x201750 vdd gnd FILL
XBUFX2_insert5 BUFX2_insert5/A BUFX2_insert5/Y vdd gnd BUFX2
XFILL_1__10045_ vdd gnd FILL
XFILL_2__12384_ vdd gnd FILL
XFILL_0__13563_ vdd gnd FILL
XFILL_0__10775_ vdd gnd FILL
XFILL_0__8061_ vdd gnd FILL
XFILL_2__14123_ vdd gnd FILL
XFILL_0__12514_ vdd gnd FILL
XFILL_1__14853_ vdd gnd FILL
X_14709_ _14709_/A _14709_/B _14709_/C _14709_/Y vdd gnd OAI21X1
X_7640_ _7640_/A _7640_/B _7640_/Y vdd gnd NOR2X1
XFILL_2__14054_ vdd gnd FILL
XFILL_1__13804_ vdd gnd FILL
XFILL_0__12445_ vdd gnd FILL
XFILL_1__14784_ vdd gnd FILL
XFILL_1__11996_ vdd gnd FILL
X_7571_ _7571_/A _7571_/B _7571_/C _7571_/Y vdd gnd OAI21X1
XFILL_2__13005_ vdd gnd FILL
XFILL_1__13735_ vdd gnd FILL
XFILL_0__12376_ vdd gnd FILL
XFILL_1__10947_ vdd gnd FILL
X_9310_ _9310_/A _9310_/B _9310_/C _9310_/Y vdd gnd OAI21X1
XFILL_0__8963_ vdd gnd FILL
XFILL_0__14115_ vdd gnd FILL
XFILL_2__10148_ vdd gnd FILL
XFILL_0__11327_ vdd gnd FILL
XFILL_1__13666_ vdd gnd FILL
XFILL_0__7914_ vdd gnd FILL
XFILL_1__10878_ vdd gnd FILL
X_9241_ _9241_/A _9241_/B _9241_/C _9241_/Y vdd gnd OAI21X1
XFILL_2__10079_ vdd gnd FILL
XFILL_0__14046_ vdd gnd FILL
XFILL_1__12617_ vdd gnd FILL
XFILL_0__11258_ vdd gnd FILL
XFILL_1__13597_ vdd gnd FILL
XFILL_0__7845_ vdd gnd FILL
X_9172_ _9172_/A _9172_/B _9172_/C _9172_/Y vdd gnd NAND3X1
XFILL_0__10209_ vdd gnd FILL
X_8123_ _8123_/A _8123_/B _8123_/Y vdd gnd AND2X2
XFILL_0__11189_ vdd gnd FILL
XFILL_0__7776_ vdd gnd FILL
XFILL_0__9515_ vdd gnd FILL
XFILL_1__12479_ vdd gnd FILL
X_8054_ _8054_/A _8054_/Y vdd gnd INVX1
XFILL_1__14218_ vdd gnd FILL
XFILL_1_BUFX2_insert20 vdd gnd FILL
XFILL_0__9446_ vdd gnd FILL
XFILL_1__14149_ vdd gnd FILL
XFILL_0__9377_ vdd gnd FILL
XFILL_1__8170_ vdd gnd FILL
XFILL_1__7121_ vdd gnd FILL
XFILL_0__8328_ vdd gnd FILL
X_8956_ _8956_/A _8956_/Y vdd gnd INVX1
X_7907_ _7907_/A _7907_/B _7907_/C _7907_/Y vdd gnd OAI21X1
XFILL_0__8259_ vdd gnd FILL
X_8887_ _8887_/D _8887_/CLK _8887_/Q vdd gnd DFFPOSX1
XFILL_1_CLKBUF1_insert32 vdd gnd FILL
X_7838_ _7838_/A _7838_/B _7838_/C _7838_/Y vdd gnd OAI21X1
XFILL_1_CLKBUF1_insert43 vdd gnd FILL
XFILL_1_CLKBUF1_insert54 vdd gnd FILL
XFILL_1_CLKBUF1_insert65 vdd gnd FILL
XFILL_1_CLKBUF1_insert76 vdd gnd FILL
XFILL_1_CLKBUF1_insert87 vdd gnd FILL
X_7769_ _7769_/A _7769_/B _7769_/Y vdd gnd NOR2X1
XFILL_1_CLKBUF1_insert98 vdd gnd FILL
X_9508_ _9508_/A _9508_/B _9508_/C _9508_/Y vdd gnd OAI21X1
X_11370_ _11370_/A _11370_/B _11370_/C _11370_/D _11370_/Y vdd gnd AOI22X1
X_9439_ _9439_/A _9439_/B _9439_/Y vdd gnd AND2X2
XFILL_1__7885_ vdd gnd FILL
X_10321_ _10321_/A _10321_/B _10321_/Y vdd gnd NAND2X1
XFILL_1__9624_ vdd gnd FILL
X_13040_ _13040_/A _13040_/B _13040_/Y vdd gnd NOR2X1
X_10252_ _10252_/A _10252_/B _10252_/Y vdd gnd AND2X2
XFILL_1__9555_ vdd gnd FILL
X_10183_ _10183_/A _10183_/B _10183_/C _10183_/Y vdd gnd AOI21X1
XFILL_1__8506_ vdd gnd FILL
XFILL257250x176550 vdd gnd FILL
XFILL_1__9486_ vdd gnd FILL
XFILL_1__8437_ vdd gnd FILL
X_13942_ _13942_/A _13942_/B _13942_/C _13942_/D _13942_/Y vdd gnd AOI22X1
XFILL_1__8368_ vdd gnd FILL
X_13873_ _13873_/A _13873_/B _13873_/Y vdd gnd NAND2X1
XFILL_1__7319_ vdd gnd FILL
XFILL_1__8299_ vdd gnd FILL
X_12824_ _12824_/A _12824_/B _12824_/C _12824_/Y vdd gnd NAND3X1
XFILL_0__10560_ vdd gnd FILL
X_12755_ _12755_/A _12755_/B _12755_/C _12755_/Y vdd gnd OAI21X1
XFILL_2__11120_ vdd gnd FILL
XFILL_1__11850_ vdd gnd FILL
XFILL_0__10491_ vdd gnd FILL
X_11706_ _11706_/A _11706_/B _11706_/C _11706_/Y vdd gnd OAI21X1
XFILL_2__11051_ vdd gnd FILL
X_12686_ _12686_/A _12686_/B _12686_/Y vdd gnd NOR2X1
XFILL_0__12230_ vdd gnd FILL
XFILL_1__10801_ vdd gnd FILL
X_14425_ _14425_/A _14425_/Y vdd gnd INVX1
XFILL_1__11781_ vdd gnd FILL
X_11637_ _11637_/D _11637_/CLK _11637_/Q vdd gnd DFFPOSX1
XFILL_1__13520_ vdd gnd FILL
XFILL_0__12161_ vdd gnd FILL
X_14356_ _14356_/A _14356_/Y vdd gnd INVX1
XFILL_2__14810_ vdd gnd FILL
X_11568_ _11568_/A _11568_/B _11568_/C _11568_/Y vdd gnd OAI21X1
XFILL_0__11112_ vdd gnd FILL
XFILL_1__10663_ vdd gnd FILL
XFILL_0__12092_ vdd gnd FILL
X_13307_ _13307_/A _13307_/B _13307_/Y vdd gnd NAND2X1
X_10519_ _10519_/A _10519_/B _10519_/C _10519_/Y vdd gnd OAI21X1
XFILL_2__8615_ vdd gnd FILL
X_14287_ _14287_/A _14287_/B _14287_/C _14287_/Y vdd gnd OAI21X1
XFILL_2__14741_ vdd gnd FILL
XFILL_1__12402_ vdd gnd FILL
X_11499_ _11499_/A _11499_/B _11499_/C _11499_/Y vdd gnd AOI21X1
XFILL_2__11953_ vdd gnd FILL
XFILL_0__11043_ vdd gnd FILL
XFILL_1__10594_ vdd gnd FILL
XFILL_1__13382_ vdd gnd FILL
XFILL_0__7630_ vdd gnd FILL
X_13238_ _13238_/A _13238_/B _13238_/Y vdd gnd NAND2X1
XFILL_2__8546_ vdd gnd FILL
XFILL_2__14672_ vdd gnd FILL
XFILL_1__12333_ vdd gnd FILL
XFILL_2__11884_ vdd gnd FILL
X_13169_ _13169_/A _13169_/B _13169_/Y vdd gnd NAND2X1
XFILL_0__7561_ vdd gnd FILL
XFILL_0__14802_ vdd gnd FILL
XFILL_1__12264_ vdd gnd FILL
XFILL_2__8477_ vdd gnd FILL
XFILL_0__9300_ vdd gnd FILL
XFILL_0__12994_ vdd gnd FILL
XFILL_0__7492_ vdd gnd FILL
XFILL_1__14003_ vdd gnd FILL
XFILL_1__11215_ vdd gnd FILL
XFILL_0__14733_ vdd gnd FILL
XFILL_1__12195_ vdd gnd FILL
XFILL_0__9231_ vdd gnd FILL
XFILL_0__11945_ vdd gnd FILL
XFILL_1__11146_ vdd gnd FILL
XFILL_0__14664_ vdd gnd FILL
XFILL_0__11876_ vdd gnd FILL
XFILL_0__9162_ vdd gnd FILL
X_8810_ _8810_/A _8810_/B _8810_/Y vdd gnd NAND2X1
X_9790_ _9790_/D _9790_/CLK _9790_/Q vdd gnd DFFPOSX1
XFILL_1__11077_ vdd gnd FILL
XFILL_0__13615_ vdd gnd FILL
XFILL_0__8113_ vdd gnd FILL
XFILL_0__10827_ vdd gnd FILL
XFILL_0__14595_ vdd gnd FILL
XFILL_2__9029_ vdd gnd FILL
XFILL_0__9093_ vdd gnd FILL
X_8741_ _8741_/A _8741_/B _8741_/Y vdd gnd NAND2X1
XFILL_1__10028_ vdd gnd FILL
XFILL_2__12367_ vdd gnd FILL
XFILL_0__13546_ vdd gnd FILL
XFILL_0__8044_ vdd gnd FILL
XFILL_2__14106_ vdd gnd FILL
X_8672_ _8672_/A _8672_/B _8672_/C _8672_/Y vdd gnd OAI21X1
XFILL_2__11318_ vdd gnd FILL
XFILL_1__14836_ vdd gnd FILL
XFILL_2__12298_ vdd gnd FILL
XFILL257250x241350 vdd gnd FILL
X_7623_ _7623_/A _7623_/B _7623_/C _7623_/Y vdd gnd NAND3X1
XFILL_2__14037_ vdd gnd FILL
XFILL_1__14767_ vdd gnd FILL
XFILL_0__12428_ vdd gnd FILL
XFILL_1__11979_ vdd gnd FILL
X_7554_ _7554_/A _7554_/B _7554_/Y vdd gnd NOR2X1
XFILL_0__9995_ vdd gnd FILL
XFILL_1__13718_ vdd gnd FILL
XFILL_0__12359_ vdd gnd FILL
XFILL_1__14698_ vdd gnd FILL
XFILL_0__8946_ vdd gnd FILL
X_7485_ _7485_/A _7485_/B _7485_/Y vdd gnd NAND2X1
XFILL_1__13649_ vdd gnd FILL
X_9224_ _9224_/A _9224_/Y vdd gnd INVX1
XFILL_1__7670_ vdd gnd FILL
XFILL_0__14029_ vdd gnd FILL
XFILL_0__7828_ vdd gnd FILL
X_9155_ _9155_/A _9155_/B _9155_/C _9155_/Y vdd gnd OAI21X1
XFILL_1__9340_ vdd gnd FILL
X_8106_ _8106_/A _8106_/Y vdd gnd INVX1
XFILL_0__7759_ vdd gnd FILL
X_9086_ _9086_/A _9086_/B _9086_/Y vdd gnd NAND2X1
XFILL_1__9271_ vdd gnd FILL
X_8037_ _8037_/A _8037_/B _8037_/Y vdd gnd NAND2X1
XFILL_0__9429_ vdd gnd FILL
XFILL257250x108150 vdd gnd FILL
XFILL_1__8222_ vdd gnd FILL
XFILL_1__8153_ vdd gnd FILL
X_9988_ _9988_/A _9988_/B _9988_/Y vdd gnd NAND2X1
XFILL_1__7104_ vdd gnd FILL
X_10870_ _10870_/A _10870_/B _10870_/C _10870_/Y vdd gnd OAI21X1
X_8939_ _8939_/A _8939_/B _8939_/Y vdd gnd NAND2X1
XFILL_1__8084_ vdd gnd FILL
X_12540_ _12540_/D _12540_/CLK _12540_/Q vdd gnd DFFPOSX1
X_12471_ _12471_/A _12471_/B _12471_/Y vdd gnd AND2X2
XFILL_1__8986_ vdd gnd FILL
X_14210_ _14210_/D _14210_/CLK _14210_/Q vdd gnd DFFPOSX1
X_11422_ _11422_/A _11422_/B _11422_/C _11422_/Y vdd gnd OAI21X1
X_14141_ _14141_/A _14141_/B _14141_/Y vdd gnd NAND2X1
X_11353_ _11353_/A _11353_/B _11353_/Y vdd gnd NOR2X1
XFILL_1__7868_ vdd gnd FILL
X_10304_ _10304_/A _10304_/B _10304_/Y vdd gnd NAND2X1
XFILL_2__8400_ vdd gnd FILL
X_14072_ _14072_/A _14072_/B _14072_/C _14072_/Y vdd gnd NAND3X1
XFILL_1__9607_ vdd gnd FILL
X_11284_ _11284_/A _11284_/B _11284_/Y vdd gnd NAND2X1
XFILL_1__7799_ vdd gnd FILL
X_13023_ _13023_/A _13023_/B _13023_/C _13023_/Y vdd gnd AOI21X1
X_10235_ _10235_/A _10235_/B _10235_/S _10235_/Y vdd gnd MUX2X1
XFILL_1__9538_ vdd gnd FILL
XFILL_2__8331_ vdd gnd FILL
X_10166_ _10166_/A _10166_/Y vdd gnd INVX1
XFILL_1__9469_ vdd gnd FILL
XFILL_2__10620_ vdd gnd FILL
XFILL_2__8262_ vdd gnd FILL
XFILL_1__11000_ vdd gnd FILL
X_10097_ _10097_/A _10097_/B _10097_/C _10097_/Y vdd gnd AOI21X1
XFILL_2__10551_ vdd gnd FILL
XFILL_0__11730_ vdd gnd FILL
XFILL_2__8193_ vdd gnd FILL
X_13925_ _13925_/A _13925_/B _13925_/C _13925_/Y vdd gnd OAI21X1
XFILL_2__13270_ vdd gnd FILL
XFILL_2__10482_ vdd gnd FILL
X_13856_ _13856_/A _13856_/B _13856_/C _13856_/Y vdd gnd NAND3X1
XFILL_0__10612_ vdd gnd FILL
XFILL_0__13400_ vdd gnd FILL
XFILL_1__12951_ vdd gnd FILL
XFILL_0__14380_ vdd gnd FILL
XFILL_0__11592_ vdd gnd FILL
X_12807_ _12807_/A _12807_/B _12807_/C _12807_/Y vdd gnd OAI21X1
XFILL_1_BUFX2_insert230 vdd gnd FILL
XFILL_1_BUFX2_insert241 vdd gnd FILL
X_13787_ _13787_/A _13787_/B _13787_/Y vdd gnd AND2X2
XFILL_1__11902_ vdd gnd FILL
X_10999_ _10999_/A _10999_/B _10999_/Y vdd gnd NAND2X1
XFILL_1_BUFX2_insert252 vdd gnd FILL
XFILL_0__10543_ vdd gnd FILL
XFILL_0__13331_ vdd gnd FILL
XFILL_1_BUFX2_insert263 vdd gnd FILL
XFILL_1_BUFX2_insert274 vdd gnd FILL
XFILL_1__12882_ vdd gnd FILL
XCLKBUF1_insert34 CLKBUF1_insert34/A CLKBUF1_insert34/Y vdd gnd CLKBUF1
XFILL_1_BUFX2_insert285 vdd gnd FILL
X_12738_ _12738_/A _12738_/B _12738_/Y vdd gnd OR2X2
XCLKBUF1_insert45 CLKBUF1_insert45/A CLKBUF1_insert45/Y vdd gnd CLKBUF1
XFILL_2__11103_ vdd gnd FILL
XFILL_1__14621_ vdd gnd FILL
XCLKBUF1_insert56 CLKBUF1_insert56/A CLKBUF1_insert56/Y vdd gnd CLKBUF1
XFILL_1_BUFX2_insert296 vdd gnd FILL
XFILL_1__11833_ vdd gnd FILL
XFILL_0__13262_ vdd gnd FILL
XCLKBUF1_insert67 CLKBUF1_insert67/A CLKBUF1_insert67/Y vdd gnd CLKBUF1
XFILL_0__10474_ vdd gnd FILL
XCLKBUF1_insert78 CLKBUF1_insert78/A CLKBUF1_insert78/Y vdd gnd CLKBUF1
XCLKBUF1_insert89 CLKBUF1_insert89/A CLKBUF1_insert89/Y vdd gnd CLKBUF1
X_12669_ _12669_/A _12669_/Y vdd gnd INVX8
XFILL_2__11034_ vdd gnd FILL
XFILL_0__12213_ vdd gnd FILL
XFILL_0__13193_ vdd gnd FILL
X_14408_ _14408_/A _14408_/B _14408_/Y vdd gnd OR2X2
XFILL_0__8800_ vdd gnd FILL
XFILL_1__11764_ vdd gnd FILL
XFILL_1__13503_ vdd gnd FILL
XFILL_0__12144_ vdd gnd FILL
XFILL_1__14483_ vdd gnd FILL
XFILL_0__8731_ vdd gnd FILL
XFILL_1__11695_ vdd gnd FILL
X_14339_ _14339_/A _14339_/B _14339_/Y vdd gnd NAND2X1
X_7270_ _7270_/A _7270_/B _7270_/C _7270_/Y vdd gnd OAI21X1
XFILL_1__10646_ vdd gnd FILL
XFILL_0__12075_ vdd gnd FILL
XFILL_0__8662_ vdd gnd FILL
XFILL_2__14724_ vdd gnd FILL
XFILL_2__11936_ vdd gnd FILL
XFILL_0__11026_ vdd gnd FILL
XFILL_1__13365_ vdd gnd FILL
XFILL_0__7613_ vdd gnd FILL
XFILL_1__10577_ vdd gnd FILL
XFILL_0__8593_ vdd gnd FILL
XFILL_2__8529_ vdd gnd FILL
XFILL_2__14655_ vdd gnd FILL
XFILL_1__12316_ vdd gnd FILL
XFILL_2__11867_ vdd gnd FILL
XFILL_1__13296_ vdd gnd FILL
XFILL_0__7544_ vdd gnd FILL
XFILL_2__13606_ vdd gnd FILL
XFILL_2__14586_ vdd gnd FILL
XFILL_1__12247_ vdd gnd FILL
XFILL_2__11798_ vdd gnd FILL
X_9911_ _9911_/A _9911_/B _9911_/C _9911_/Y vdd gnd OAI21X1
XFILL_0__12977_ vdd gnd FILL
XFILL_0__7475_ vdd gnd FILL
XFILL_2__13537_ vdd gnd FILL
XFILL_0__14716_ vdd gnd FILL
XFILL_0__9214_ vdd gnd FILL
XFILL_0__11928_ vdd gnd FILL
XFILL_1__12178_ vdd gnd FILL
X_9842_ _9842_/D _9842_/CLK _9842_/Q vdd gnd DFFPOSX1
XFILL_1__11129_ vdd gnd FILL
XFILL_0__14647_ vdd gnd FILL
XFILL_0__9145_ vdd gnd FILL
XFILL_0__11859_ vdd gnd FILL
X_9773_ _9773_/D _9773_/CLK _9773_/Q vdd gnd DFFPOSX1
XFILL_0__14578_ vdd gnd FILL
XFILL_0__9076_ vdd gnd FILL
X_8724_ _8724_/A _8724_/B _8724_/Y vdd gnd NOR2X1
XFILL_0__13529_ vdd gnd FILL
XFILL_0__8027_ vdd gnd FILL
X_8655_ _8655_/A _8655_/Y vdd gnd INVX1
XFILL_1__14819_ vdd gnd FILL
X_7606_ _7606_/A _7606_/Y vdd gnd INVX1
X_8586_ _8586_/A _8586_/B _8586_/Y vdd gnd OR2X2
X_7537_ _7537_/A _7537_/B _7537_/C _7537_/Y vdd gnd NAND3X1
XFILL_1__8771_ vdd gnd FILL
XFILL_0__9978_ vdd gnd FILL
XFILL_1__7722_ vdd gnd FILL
XFILL_0__8929_ vdd gnd FILL
X_7468_ _7468_/A _7468_/B _7468_/Y vdd gnd NAND2X1
X_9207_ _9207_/A _9207_/B _9207_/Y vdd gnd NOR2X1
XFILL_1__7653_ vdd gnd FILL
X_7399_ _7399_/A _7399_/B _7399_/Y vdd gnd NAND2X1
X_9138_ _9138_/A _9138_/B _9138_/C _9138_/Y vdd gnd OAI21X1
XFILL_1__7584_ vdd gnd FILL
X_10020_ _10020_/A _10020_/Y vdd gnd INVX1
XFILL_1__9323_ vdd gnd FILL
X_9069_ _9069_/A _9069_/B _9069_/C _9069_/Y vdd gnd NAND3X1
XFILL_1__9254_ vdd gnd FILL
XFILL_1__8205_ vdd gnd FILL
X_11971_ _11971_/A _11971_/Y vdd gnd INVX1
XFILL_1__9185_ vdd gnd FILL
X_13710_ _13710_/A _13710_/B _13710_/C _13710_/Y vdd gnd OAI21X1
X_10922_ _10922_/A _10922_/B _10922_/C _10922_/Y vdd gnd OAI21X1
X_14690_ _14690_/A _14690_/B _14690_/C _14690_/Y vdd gnd OAI21X1
XFILL_1__8136_ vdd gnd FILL
X_13641_ _13641_/A _13641_/B _13641_/C _13641_/Y vdd gnd AOI21X1
X_10853_ _10853_/A _10853_/Y vdd gnd INVX8
XFILL_1__8067_ vdd gnd FILL
X_13572_ _13572_/A _13572_/B _13572_/Y vdd gnd NAND2X1
X_10784_ _10784_/A _10784_/B _10784_/C _10784_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert204 vdd gnd FILL
XFILL_0_BUFX2_insert215 vdd gnd FILL
X_12523_ _12523_/A _12523_/B _12523_/C _12523_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert226 vdd gnd FILL
XFILL_0_BUFX2_insert237 vdd gnd FILL
XFILL_0_BUFX2_insert248 vdd gnd FILL
XFILL_0_BUFX2_insert259 vdd gnd FILL
X_12454_ _12454_/A _12454_/B _12454_/Y vdd gnd NOR2X1
XFILL_1__8969_ vdd gnd FILL
XFILL_0__10190_ vdd gnd FILL
X_11405_ _11405_/A _11405_/B _11405_/C _11405_/Y vdd gnd OAI21X1
X_12385_ _12385_/A _12385_/B _12385_/C _12385_/Y vdd gnd OAI21X1
XFILL_1__10500_ vdd gnd FILL
XFILL_1__11480_ vdd gnd FILL
X_14124_ _14124_/A _14124_/B _14124_/C _14124_/Y vdd gnd OAI21X1
X_11336_ _11336_/A _11336_/B _11336_/Y vdd gnd NOR2X1
XFILL_1__10431_ vdd gnd FILL
X_14055_ _14055_/A _14055_/B _14055_/Y vdd gnd NOR2X1
X_11267_ _11267_/A _11267_/B _11267_/C _11267_/Y vdd gnd OAI21X1
XFILL_1__13150_ vdd gnd FILL
XFILL_1__10362_ vdd gnd FILL
XFILL_0__12900_ vdd gnd FILL
X_13006_ _13006_/A _13006_/B _13006_/C _13006_/Y vdd gnd OAI21X1
X_10218_ _10218_/A _10218_/B _10218_/C _10218_/Y vdd gnd OAI21X1
XFILL_0__13880_ vdd gnd FILL
XFILL_2__14440_ vdd gnd FILL
XFILL_1__12101_ vdd gnd FILL
X_11198_ _11198_/A _11198_/B _11198_/C _11198_/Y vdd gnd AOI21X1
XFILL_1__13081_ vdd gnd FILL
XFILL_1__10293_ vdd gnd FILL
XFILL_0__12831_ vdd gnd FILL
X_10149_ _10149_/A _10149_/B _10149_/C _10149_/Y vdd gnd AOI21X1
XFILL_1__12032_ vdd gnd FILL
XFILL_2__14371_ vdd gnd FILL
XFILL_0__12762_ vdd gnd FILL
XFILL_0__7260_ vdd gnd FILL
XFILL_2__13322_ vdd gnd FILL
XFILL_2__8176_ vdd gnd FILL
XFILL_0__11713_ vdd gnd FILL
X_13908_ _13908_/A _13908_/B _13908_/Y vdd gnd NAND2X1
XFILL_0__12693_ vdd gnd FILL
XFILL_0__7191_ vdd gnd FILL
XFILL_2__7127_ vdd gnd FILL
X_14888_ _14888_/D _14888_/CLK _14888_/Q vdd gnd DFFPOSX1
XFILL_2__13253_ vdd gnd FILL
XFILL_2__10465_ vdd gnd FILL
XFILL_0__14432_ vdd gnd FILL
XFILL_1__13983_ vdd gnd FILL
X_13839_ _13839_/A _13839_/B _13839_/Y vdd gnd NAND2X1
XFILL_2__13184_ vdd gnd FILL
XFILL_1__12934_ vdd gnd FILL
XFILL_2__10396_ vdd gnd FILL
XFILL_0__14363_ vdd gnd FILL
XFILL_0__11575_ vdd gnd FILL
XFILL_0__10526_ vdd gnd FILL
XFILL_0__13314_ vdd gnd FILL
XFILL_1__12865_ vdd gnd FILL
XFILL_0__9901_ vdd gnd FILL
XFILL_0__14294_ vdd gnd FILL
X_8440_ _8440_/A _8440_/B _8440_/Y vdd gnd NAND2X1
XFILL_1__14604_ vdd gnd FILL
XFILL_1__11816_ vdd gnd FILL
XFILL_0__10457_ vdd gnd FILL
XFILL_0__13245_ vdd gnd FILL
XFILL_1__12796_ vdd gnd FILL
X_8371_ _8371_/A _8371_/B _8371_/S _8371_/Y vdd gnd MUX2X1
XFILL_2__11017_ vdd gnd FILL
XFILL_0__13176_ vdd gnd FILL
XFILL_1__11747_ vdd gnd FILL
XFILL_0__10388_ vdd gnd FILL
X_7322_ _7322_/A _7322_/B _7322_/C _7322_/Y vdd gnd AOI21X1
XFILL_0__9763_ vdd gnd FILL
XFILL_0__12127_ vdd gnd FILL
XFILL_1__14466_ vdd gnd FILL
XFILL_0__8714_ vdd gnd FILL
X_7253_ _7253_/A _7253_/B _7253_/Y vdd gnd NAND2X1
XFILL_0__9694_ vdd gnd FILL
XFILL_1__13417_ vdd gnd FILL
XFILL_1__10629_ vdd gnd FILL
XFILL_0__12058_ vdd gnd FILL
XFILL_1__14397_ vdd gnd FILL
XFILL_0__8645_ vdd gnd FILL
X_7184_ _7184_/A _7184_/B _7184_/C _7184_/Y vdd gnd OAI21X1
XFILL_0__11009_ vdd gnd FILL
XFILL_2__11919_ vdd gnd FILL
XFILL_1__13348_ vdd gnd FILL
XFILL_0__8576_ vdd gnd FILL
XFILL_1__13279_ vdd gnd FILL
XFILL_0__7527_ vdd gnd FILL
XFILL_1_BUFX2_insert5 vdd gnd FILL
XFILL_0__7458_ vdd gnd FILL
X_9825_ _9825_/D _9825_/CLK _9825_/Q vdd gnd DFFPOSX1
XFILL_0__7389_ vdd gnd FILL
XFILL_0__9128_ vdd gnd FILL
X_9756_ _9756_/A _9756_/B _9756_/C _9756_/Y vdd gnd OAI21X1
XFILL_0__9059_ vdd gnd FILL
X_8707_ _8707_/A _8707_/Y vdd gnd INVX1
XFILL_1__9941_ vdd gnd FILL
XBUFX2_insert309 BUFX2_insert309/A BUFX2_insert309/Y vdd gnd BUFX2
X_9687_ _9687_/A _9687_/Y vdd gnd INVX1
X_8638_ _8638_/A _8638_/B _8638_/Y vdd gnd OR2X2
XFILL_1__9872_ vdd gnd FILL
XFILL_1__8823_ vdd gnd FILL
X_8569_ _8569_/A _8569_/B _8569_/Y vdd gnd NAND2X1
XFILL_1__8754_ vdd gnd FILL
XFILL_1__7705_ vdd gnd FILL
X_12170_ _12170_/A _12170_/B _12170_/C _12170_/D _12170_/Y vdd gnd AOI22X1
XFILL_1__8685_ vdd gnd FILL
X_11121_ _11121_/A _11121_/B _11121_/Y vdd gnd NAND2X1
XFILL_1__7636_ vdd gnd FILL
X_11052_ _11052_/A _11052_/B _11052_/Y vdd gnd OR2X2
XFILL_1__7567_ vdd gnd FILL
X_10003_ _10003_/A _10003_/Y vdd gnd INVX1
XFILL_1__9306_ vdd gnd FILL
XFILL_1__7498_ vdd gnd FILL
X_14811_ _14811_/A _14811_/B _14811_/Y vdd gnd NOR2X1
XFILL_1__9237_ vdd gnd FILL
X_14742_ _14742_/A _14742_/B _14742_/Y vdd gnd NAND2X1
X_11954_ _11954_/A _11954_/B _11954_/C _11954_/Y vdd gnd NAND3X1
XFILL_1__9168_ vdd gnd FILL
X_10905_ _10905_/A _10905_/B _10905_/S _10905_/Y vdd gnd MUX2X1
X_14673_ _14673_/A _14673_/B _14673_/Y vdd gnd NAND2X1
XFILL_1__8119_ vdd gnd FILL
X_11885_ _11885_/A _11885_/B _11885_/C _11885_/Y vdd gnd OAI21X1
XFILL_1__9099_ vdd gnd FILL
XFILL_2__9981_ vdd gnd FILL
XFILL_1__10980_ vdd gnd FILL
X_13624_ _13624_/A _13624_/B _13624_/S _13624_/Y vdd gnd MUX2X1
X_10836_ _10836_/A _10836_/B _10836_/S _10836_/Y vdd gnd MUX2X1
XFILL_0__11360_ vdd gnd FILL
X_13555_ _13555_/A _13555_/Y vdd gnd INVX1
X_10767_ _10767_/D _10767_/CLK _10767_/Q vdd gnd DFFPOSX1
XFILL_0__10311_ vdd gnd FILL
XFILL_1__12650_ vdd gnd FILL
X_12506_ _12506_/A _12506_/B _12506_/Y vdd gnd NAND2X1
XFILL_0__11291_ vdd gnd FILL
X_13486_ _13486_/D _13486_/CLK _13486_/Q vdd gnd DFFPOSX1
X_10698_ _10698_/D _10698_/CLK _10698_/Q vdd gnd DFFPOSX1
XFILL_1__11601_ vdd gnd FILL
XFILL_0__13030_ vdd gnd FILL
XFILL_0__10242_ vdd gnd FILL
XFILL_2__8794_ vdd gnd FILL
X_12437_ _12437_/A _12437_/B _12437_/Y vdd gnd NAND2X1
XFILL_1__14320_ vdd gnd FILL
XFILL_1__11532_ vdd gnd FILL
XFILL_0__10173_ vdd gnd FILL
X_12368_ _12368_/A _12368_/B _12368_/C _12368_/Y vdd gnd OAI21X1
XFILL_2__12822_ vdd gnd FILL
XFILL_1__14251_ vdd gnd FILL
XFILL_1__11463_ vdd gnd FILL
X_14107_ _14107_/A _14107_/B _14107_/Y vdd gnd OR2X2
X_11319_ _11319_/A _11319_/B _11319_/C _11319_/Y vdd gnd NAND3X1
XFILL_1__13202_ vdd gnd FILL
XFILL_2__9415_ vdd gnd FILL
X_12299_ _12299_/A _12299_/B _12299_/Y vdd gnd NOR2X1
XFILL_1__10414_ vdd gnd FILL
XFILL_0__13932_ vdd gnd FILL
XFILL_0__8430_ vdd gnd FILL
XFILL_1__11394_ vdd gnd FILL
X_14038_ _14038_/A _14038_/Y vdd gnd INVX1
XFILL_2__9346_ vdd gnd FILL
XFILL_1__13133_ vdd gnd FILL
XFILL_1__10345_ vdd gnd FILL
XFILL_0__13863_ vdd gnd FILL
XFILL_0__8361_ vdd gnd FILL
XFILL_2__14423_ vdd gnd FILL
XFILL_1__10276_ vdd gnd FILL
XFILL_0__12814_ vdd gnd FILL
XFILL_1__13064_ vdd gnd FILL
XFILL_0__7312_ vdd gnd FILL
XFILL_0__13794_ vdd gnd FILL
X_7940_ _7940_/D _7940_/CLK _7940_/Q vdd gnd DFFPOSX1
XFILL_0__8292_ vdd gnd FILL
XFILL_2__14354_ vdd gnd FILL
XFILL_1__12015_ vdd gnd FILL
XFILL_0__12745_ vdd gnd FILL
XFILL_0__7243_ vdd gnd FILL
XFILL_2__13305_ vdd gnd FILL
X_7871_ _7871_/A _7871_/Y vdd gnd INVX1
XFILL_2__14285_ vdd gnd FILL
X_9610_ _9610_/A _9610_/B _9610_/Y vdd gnd NAND2X1
XFILL_0__12676_ vdd gnd FILL
XFILL_0__7174_ vdd gnd FILL
XFILL_2__13236_ vdd gnd FILL
XFILL_0__14415_ vdd gnd FILL
XFILL_1__13966_ vdd gnd FILL
X_9541_ _9541_/A _9541_/B _9541_/Y vdd gnd NAND2X1
XFILL_2__13167_ vdd gnd FILL
XFILL_1__12917_ vdd gnd FILL
XFILL_0__14346_ vdd gnd FILL
XFILL_1__13897_ vdd gnd FILL
XFILL_0__11558_ vdd gnd FILL
X_9472_ _9472_/A _9472_/Y vdd gnd INVX1
XFILL_0__10509_ vdd gnd FILL
XFILL_1__12848_ vdd gnd FILL
XFILL_2__13098_ vdd gnd FILL
XFILL_0__14277_ vdd gnd FILL
XFILL_0__11489_ vdd gnd FILL
X_8423_ _8423_/A _8423_/B _8423_/C _8423_/Y vdd gnd OAI21X1
XFILL_0__13228_ vdd gnd FILL
XFILL_1__12779_ vdd gnd FILL
X_8354_ _8354_/A _8354_/B _8354_/C _8354_/Y vdd gnd AOI21X1
XFILL_0__13159_ vdd gnd FILL
X_7305_ _7305_/A _7305_/B _7305_/C _7305_/Y vdd gnd NAND3X1
XFILL_0__9746_ vdd gnd FILL
X_8285_ _8285_/A _8285_/B _8285_/C _8285_/Y vdd gnd OAI21X1
XFILL_1__14449_ vdd gnd FILL
X_7236_ _7236_/A _7236_/B _7236_/C _7236_/Y vdd gnd NAND3X1
XFILL_0__9677_ vdd gnd FILL
XFILL_1__8470_ vdd gnd FILL
XFILL_1__7421_ vdd gnd FILL
XFILL_0__8628_ vdd gnd FILL
X_7167_ _7167_/A _7167_/B _7167_/C _7167_/Y vdd gnd NAND3X1
XFILL_1__7352_ vdd gnd FILL
XFILL_0__8559_ vdd gnd FILL
X_7098_ _7098_/A _7098_/B _7098_/C _7098_/Y vdd gnd AOI21X1
XFILL_2_BUFX2_insert129 vdd gnd FILL
XFILL_1__7283_ vdd gnd FILL
XFILL_1__9022_ vdd gnd FILL
X_9808_ _9808_/D _9808_/CLK _9808_/Q vdd gnd DFFPOSX1
XFILL256950x150 vdd gnd FILL
X_11670_ _11670_/D _11670_/CLK _11670_/Q vdd gnd DFFPOSX1
X_9739_ _9739_/A _9739_/B _9739_/C _9739_/Y vdd gnd OAI21X1
X_10621_ _10621_/A _10621_/B _10621_/Y vdd gnd NAND2X1
XBUFX2_insert117 BUFX2_insert117/A BUFX2_insert117/Y vdd gnd BUFX2
XBUFX2_insert128 BUFX2_insert128/A BUFX2_insert128/Y vdd gnd BUFX2
XBUFX2_insert139 BUFX2_insert139/A BUFX2_insert139/Y vdd gnd BUFX2
XFILL_1__9924_ vdd gnd FILL
X_13340_ _13340_/A _13340_/B _13340_/Y vdd gnd NAND2X1
X_10552_ _10552_/A _10552_/B _10552_/C _10552_/Y vdd gnd OAI21X1
XFILL_1__9855_ vdd gnd FILL
X_13271_ _13271_/A _13271_/B _13271_/Y vdd gnd NAND2X1
X_10483_ _10483_/A _10483_/B _10483_/C _10483_/Y vdd gnd OAI21X1
XFILL_1__8806_ vdd gnd FILL
X_12222_ _12222_/A _12222_/B _12222_/Y vdd gnd NOR2X1
XFILL_1__8737_ vdd gnd FILL
X_12153_ _12153_/A _12153_/B _12153_/C _12153_/Y vdd gnd OAI21X1
XFILL_1__8668_ vdd gnd FILL
X_11104_ _11104_/A _11104_/B _11104_/C _11104_/Y vdd gnd AOI21X1
XFILL_2__9200_ vdd gnd FILL
X_12084_ _12084_/A _12084_/B _12084_/Y vdd gnd NAND2X1
XFILL_1__7619_ vdd gnd FILL
XFILL_1__8599_ vdd gnd FILL
X_11035_ _11035_/A _11035_/B _11035_/C _11035_/Y vdd gnd NAND3X1
XFILL_2__9131_ vdd gnd FILL
XFILL_1__10130_ vdd gnd FILL
XFILL_2_CLKBUF1_insert387 vdd gnd FILL
XFILL_0__10860_ vdd gnd FILL
XFILL_2__9062_ vdd gnd FILL
XFILL_2__11420_ vdd gnd FILL
XFILL_1__10061_ vdd gnd FILL
XFILL_0__10791_ vdd gnd FILL
X_12986_ _12986_/A _12986_/B _12986_/Y vdd gnd AND2X2
XFILL_2__11351_ vdd gnd FILL
XFILL_0__12530_ vdd gnd FILL
X_14725_ _14725_/A _14725_/B _14725_/Y vdd gnd NAND2X1
X_11937_ _11937_/A _11937_/B _11937_/Y vdd gnd NAND2X1
XFILL_2__14070_ vdd gnd FILL
XFILL_1__13820_ vdd gnd FILL
XFILL_2__11282_ vdd gnd FILL
XFILL_0__12461_ vdd gnd FILL
X_14656_ _14656_/A _14656_/B _14656_/C _14656_/Y vdd gnd AOI21X1
X_11868_ _11868_/A _11868_/Y vdd gnd INVX1
XFILL_2__9964_ vdd gnd FILL
XFILL_0__11412_ vdd gnd FILL
XFILL_1__13751_ vdd gnd FILL
XFILL_1__10963_ vdd gnd FILL
XFILL_0__12392_ vdd gnd FILL
X_10819_ _10819_/A _10819_/Y vdd gnd INVX1
X_13607_ _13607_/A _13607_/B _13607_/S _13607_/Y vdd gnd MUX2X1
X_14587_ _14587_/A _14587_/Y vdd gnd INVX1
X_11799_ _11799_/A _11799_/Y vdd gnd INVX1
XFILL_1__12702_ vdd gnd FILL
XFILL_0__11343_ vdd gnd FILL
XFILL_0__14131_ vdd gnd FILL
XFILL_2__9895_ vdd gnd FILL
XFILL_1__13682_ vdd gnd FILL
XFILL_1__10894_ vdd gnd FILL
X_13538_ _13538_/A _13538_/B _13538_/Y vdd gnd NOR2X1
XFILL_1__12633_ vdd gnd FILL
XFILL_0__14062_ vdd gnd FILL
XFILL_0__11274_ vdd gnd FILL
XFILL_0__7861_ vdd gnd FILL
X_13469_ _13469_/D _13469_/CLK _13469_/Q vdd gnd DFFPOSX1
XFILL_2__13923_ vdd gnd FILL
XFILL_0__10225_ vdd gnd FILL
XFILL_0__13013_ vdd gnd FILL
XFILL_2__8777_ vdd gnd FILL
XFILL_0__9600_ vdd gnd FILL
XFILL_0__7792_ vdd gnd FILL
XFILL_1__14303_ vdd gnd FILL
XFILL_1__11515_ vdd gnd FILL
XFILL_2__13854_ vdd gnd FILL
XFILL_0__10156_ vdd gnd FILL
XFILL_0__9531_ vdd gnd FILL
XFILL_1__12495_ vdd gnd FILL
X_8070_ _8070_/A _8070_/B _8070_/C _8070_/Y vdd gnd OAI21X1
XFILL_1__14234_ vdd gnd FILL
XFILL_2__12805_ vdd gnd FILL
XFILL_1__11446_ vdd gnd FILL
XFILL_0__10087_ vdd gnd FILL
XFILL_0__9462_ vdd gnd FILL
XFILL_2__12736_ vdd gnd FILL
XFILL_0__13915_ vdd gnd FILL
XFILL_0__8413_ vdd gnd FILL
XFILL_1__11377_ vdd gnd FILL
XFILL_0__9393_ vdd gnd FILL
XFILL_1__13116_ vdd gnd FILL
XFILL_2__9329_ vdd gnd FILL
XFILL_1__10328_ vdd gnd FILL
XFILL_2__12667_ vdd gnd FILL
XFILL_1__14096_ vdd gnd FILL
XFILL_0__13846_ vdd gnd FILL
XFILL_0__8344_ vdd gnd FILL
X_8972_ _8972_/A _8972_/B _8972_/Y vdd gnd NOR2X1
XFILL_2__14406_ vdd gnd FILL
XFILL_1__13047_ vdd gnd FILL
XFILL_1__10259_ vdd gnd FILL
XFILL_0__13777_ vdd gnd FILL
XFILL_0__10989_ vdd gnd FILL
X_7923_ _7923_/D _7923_/CLK _7923_/Q vdd gnd DFFPOSX1
XFILL_0__8275_ vdd gnd FILL
XFILL_2__14337_ vdd gnd FILL
XFILL_2__11549_ vdd gnd FILL
XFILL_0__12728_ vdd gnd FILL
XFILL_0__7226_ vdd gnd FILL
X_7854_ _7854_/A _7854_/B _7854_/Y vdd gnd NAND2X1
XFILL_2__14268_ vdd gnd FILL
XFILL_0__12659_ vdd gnd FILL
XFILL_0__7157_ vdd gnd FILL
X_7785_ _7785_/A _7785_/B _7785_/Y vdd gnd OR2X2
XFILL_1__13949_ vdd gnd FILL
X_9524_ _9524_/A _9524_/Y vdd gnd INVX1
XFILL_0__7088_ vdd gnd FILL
XFILL_0__14329_ vdd gnd FILL
X_9455_ _9455_/A _9455_/B _9455_/C _9455_/Y vdd gnd OAI21X1
X_8406_ _8406_/A _8406_/B _8406_/Y vdd gnd OR2X2
XFILL_1__9640_ vdd gnd FILL
X_9386_ _9386_/A _9386_/B _9386_/C _9386_/Y vdd gnd OAI21X1
XFILL_1__9571_ vdd gnd FILL
X_8337_ _8337_/A _8337_/B _8337_/C _8337_/Y vdd gnd NAND3X1
XFILL_1__8522_ vdd gnd FILL
XFILL_0__9729_ vdd gnd FILL
X_8268_ _8268_/A _8268_/B _8268_/Y vdd gnd NOR2X1
X_7219_ _7219_/A _7219_/B _7219_/Y vdd gnd NAND2X1
XFILL_1__8453_ vdd gnd FILL
X_8199_ _8199_/A _8199_/B _8199_/Y vdd gnd NAND2X1
XFILL_1__7404_ vdd gnd FILL
XFILL_1__8384_ vdd gnd FILL
XFILL_1__7335_ vdd gnd FILL
X_12840_ _12840_/A _12840_/B _12840_/Y vdd gnd NAND2X1
XFILL_1__7266_ vdd gnd FILL
XFILL_1__9005_ vdd gnd FILL
X_12771_ _12771_/A _12771_/Y vdd gnd INVX1
XFILL_1__7197_ vdd gnd FILL
X_14510_ _14510_/D _14510_/CLK _14510_/Q vdd gnd DFFPOSX1
X_11722_ _11722_/A _11722_/B _11722_/C _11722_/Y vdd gnd OAI21X1
X_14441_ _14441_/A _14441_/B _14441_/C _14441_/Y vdd gnd OAI21X1
X_11653_ _11653_/D _11653_/CLK _11653_/Q vdd gnd DFFPOSX1
X_10604_ _10604_/A _10604_/B _10604_/Y vdd gnd NAND2X1
X_14372_ _14372_/A _14372_/B _14372_/Y vdd gnd OR2X2
XFILL_1__9907_ vdd gnd FILL
X_11584_ _11584_/A _11584_/B _11584_/Y vdd gnd NAND2X1
X_13323_ _13323_/A _13323_/B _13323_/C _13323_/Y vdd gnd AOI21X1
X_10535_ _10535_/A _10535_/Y vdd gnd INVX1
X_13254_ _13254_/A _13254_/B _13254_/Y vdd gnd NOR2X1
X_10466_ _10466_/A _10466_/Y vdd gnd INVX1
XFILL_0__10010_ vdd gnd FILL
XFILL_2__10920_ vdd gnd FILL
X_12205_ _12205_/A _12205_/B _12205_/C _12205_/Y vdd gnd AOI21X1
X_13185_ _13185_/A _13185_/B _13185_/Y vdd gnd NAND2X1
XFILL_1__11300_ vdd gnd FILL
X_10397_ _10397_/A _10397_/B _10397_/C _10397_/Y vdd gnd OAI21X1
XFILL_2__7513_ vdd gnd FILL
XFILL_2__8493_ vdd gnd FILL
XFILL_1__12280_ vdd gnd FILL
X_12136_ _12136_/A _12136_/B _12136_/Y vdd gnd NAND2X1
XFILL_1__11231_ vdd gnd FILL
XFILL_2__13570_ vdd gnd FILL
XFILL_0__11961_ vdd gnd FILL
X_12067_ _12067_/A _12067_/B _12067_/S _12067_/Y vdd gnd MUX2X1
XFILL_0__13700_ vdd gnd FILL
XFILL_1__11162_ vdd gnd FILL
XFILL_0__10912_ vdd gnd FILL
X_11018_ _11018_/A _11018_/B _11018_/C _11018_/Y vdd gnd AOI21X1
XFILL_0__14680_ vdd gnd FILL
XFILL_0__11892_ vdd gnd FILL
XFILL_2__9114_ vdd gnd FILL
XFILL_1__10113_ vdd gnd FILL
XFILL_0__13631_ vdd gnd FILL
XFILL_1__11093_ vdd gnd FILL
XFILL_0__10843_ vdd gnd FILL
XFILL_2__9045_ vdd gnd FILL
XFILL_2__11403_ vdd gnd FILL
XFILL_1__10044_ vdd gnd FILL
XBUFX2_insert6 BUFX2_insert6/A BUFX2_insert6/Y vdd gnd BUFX2
XFILL_0__13562_ vdd gnd FILL
XFILL_0__8060_ vdd gnd FILL
XFILL_0__10774_ vdd gnd FILL
X_12969_ _12969_/A _12969_/B _12969_/C _12969_/Y vdd gnd OAI21X1
XFILL_2__11334_ vdd gnd FILL
XFILL_1__14852_ vdd gnd FILL
XFILL_0__12513_ vdd gnd FILL
X_14708_ _14708_/A _14708_/B _14708_/Y vdd gnd NOR2X1
XFILL_1__13803_ vdd gnd FILL
XFILL_2__11265_ vdd gnd FILL
XFILL_1__14783_ vdd gnd FILL
XFILL_0__12444_ vdd gnd FILL
XFILL_1__11995_ vdd gnd FILL
X_14639_ _14639_/A _14639_/B _14639_/Y vdd gnd AND2X2
X_7570_ _7570_/A _7570_/B _7570_/C _7570_/Y vdd gnd OAI21X1
XFILL_2__9947_ vdd gnd FILL
XFILL_1__13734_ vdd gnd FILL
XFILL_2__11196_ vdd gnd FILL
XFILL_1__10946_ vdd gnd FILL
XFILL_0__12375_ vdd gnd FILL
XFILL_0__8962_ vdd gnd FILL
XFILL_0__14114_ vdd gnd FILL
XFILL_1__13665_ vdd gnd FILL
XFILL_2__9878_ vdd gnd FILL
XFILL_0__11326_ vdd gnd FILL
XFILL_1__10877_ vdd gnd FILL
X_9240_ _9240_/A _9240_/B _9240_/C _9240_/Y vdd gnd OAI21X1
XFILL_0__7913_ vdd gnd FILL
XFILL_2__8829_ vdd gnd FILL
XFILL_1__12616_ vdd gnd FILL
XFILL_0__14045_ vdd gnd FILL
XFILL_0__11257_ vdd gnd FILL
XFILL_1__13596_ vdd gnd FILL
XFILL_0__7844_ vdd gnd FILL
X_9171_ _9171_/A _9171_/B _9171_/Y vdd gnd AND2X2
XFILL_2__13906_ vdd gnd FILL
XFILL_0__10208_ vdd gnd FILL
XFILL_0__11188_ vdd gnd FILL
X_8122_ _8122_/A _8122_/B _8122_/C _8122_/Y vdd gnd NAND3X1
XFILL_0__7775_ vdd gnd FILL
XFILL_0__10139_ vdd gnd FILL
XFILL_2__13837_ vdd gnd FILL
XFILL_1__12478_ vdd gnd FILL
XFILL_0__9514_ vdd gnd FILL
X_8053_ _8053_/A _8053_/B _8053_/C _8053_/Y vdd gnd OAI21X1
XFILL_1__14217_ vdd gnd FILL
XFILL_1_BUFX2_insert10 vdd gnd FILL
XFILL_1__11429_ vdd gnd FILL
XFILL_2__13768_ vdd gnd FILL
XFILL_1_BUFX2_insert21 vdd gnd FILL
XFILL_0__9445_ vdd gnd FILL
XFILL_2__12719_ vdd gnd FILL
XFILL_1__14148_ vdd gnd FILL
XFILL_2__13699_ vdd gnd FILL
XFILL_0__9376_ vdd gnd FILL
XFILL_1__14079_ vdd gnd FILL
XFILL_0__13829_ vdd gnd FILL
XFILL_1__7120_ vdd gnd FILL
XFILL_0__8327_ vdd gnd FILL
X_8955_ _8955_/A _8955_/B _8955_/C _8955_/Y vdd gnd AOI21X1
X_7906_ _7906_/A _7906_/B _7906_/Y vdd gnd NAND2X1
XFILL_0__8258_ vdd gnd FILL
X_8886_ _8886_/D _8886_/CLK _8886_/Q vdd gnd DFFPOSX1
XFILL_0__7209_ vdd gnd FILL
X_7837_ _7837_/A _7837_/B _7837_/Y vdd gnd NAND2X1
XFILL_0__8189_ vdd gnd FILL
XFILL_1_CLKBUF1_insert33 vdd gnd FILL
XFILL_1_CLKBUF1_insert44 vdd gnd FILL
XFILL_1_CLKBUF1_insert55 vdd gnd FILL
XFILL_1_CLKBUF1_insert66 vdd gnd FILL
X_7768_ _7768_/A _7768_/B _7768_/C _7768_/Y vdd gnd OAI21X1
XFILL_1_CLKBUF1_insert77 vdd gnd FILL
XFILL_1_CLKBUF1_insert88 vdd gnd FILL
XFILL_1_CLKBUF1_insert99 vdd gnd FILL
X_9507_ _9507_/A _9507_/B _9507_/C _9507_/Y vdd gnd OAI21X1
X_7699_ _7699_/A _7699_/B _7699_/Y vdd gnd AND2X2
X_9438_ _9438_/A _9438_/B _9438_/Y vdd gnd AND2X2
XFILL_1__7884_ vdd gnd FILL
X_10320_ _10320_/A _10320_/B _10320_/Y vdd gnd NAND2X1
XFILL_1__9623_ vdd gnd FILL
X_9369_ _9369_/A _9369_/B _9369_/C _9369_/Y vdd gnd AOI21X1
X_10251_ _10251_/A _10251_/B _10251_/C _10251_/Y vdd gnd NAND3X1
XFILL256950x165750 vdd gnd FILL
XFILL_1__9554_ vdd gnd FILL
X_10182_ _10182_/A _10182_/B _10182_/C _10182_/Y vdd gnd NAND3X1
XFILL_1__8505_ vdd gnd FILL
XFILL_1__9485_ vdd gnd FILL
XFILL_1__8436_ vdd gnd FILL
X_13941_ _13941_/A _13941_/B _13941_/Y vdd gnd NAND2X1
XFILL_2__7160_ vdd gnd FILL
XFILL_1__8367_ vdd gnd FILL
XFILL_1__7318_ vdd gnd FILL
X_13872_ _13872_/A _13872_/B _13872_/Y vdd gnd NOR2X1
XFILL_2__7091_ vdd gnd FILL
XFILL_1__8298_ vdd gnd FILL
X_12823_ _12823_/A _12823_/B _12823_/C _12823_/Y vdd gnd OAI21X1
XFILL_1__7249_ vdd gnd FILL
XFILL257250x64950 vdd gnd FILL
X_12754_ _12754_/A _12754_/Y vdd gnd INVX1
XFILL_0__10490_ vdd gnd FILL
X_11705_ _11705_/A _11705_/B _11705_/C _11705_/D _11705_/Y vdd gnd AOI22X1
X_12685_ _12685_/A _12685_/B _12685_/S _12685_/Y vdd gnd MUX2X1
XFILL_1__10800_ vdd gnd FILL
XFILL_1__11780_ vdd gnd FILL
X_14424_ _14424_/A _14424_/B _14424_/Y vdd gnd NAND2X1
X_11636_ _11636_/D _11636_/CLK _11636_/Q vdd gnd DFFPOSX1
XFILL_2__10001_ vdd gnd FILL
XFILL_2__9732_ vdd gnd FILL
XFILL_0__12160_ vdd gnd FILL
X_14355_ _14355_/A _14355_/B _14355_/C _14355_/Y vdd gnd OAI21X1
X_11567_ _11567_/A _11567_/Y vdd gnd INVX1
XFILL_0__11111_ vdd gnd FILL
XFILL_1__10662_ vdd gnd FILL
XFILL_0__12091_ vdd gnd FILL
X_10518_ _10518_/A _10518_/B _10518_/C _10518_/Y vdd gnd OAI21X1
X_13306_ _13306_/A _13306_/B _13306_/Y vdd gnd OR2X2
X_14286_ _14286_/A _14286_/Y vdd gnd INVX1
XFILL_1__12401_ vdd gnd FILL
X_11498_ _11498_/A _11498_/B _11498_/Y vdd gnd NOR2X1
XFILL_0__11042_ vdd gnd FILL
XFILL_1__13381_ vdd gnd FILL
XFILL_1__10593_ vdd gnd FILL
X_13237_ _13237_/A _13237_/B _13237_/Y vdd gnd NAND2X1
X_10449_ _10449_/A _10449_/B _10449_/C _10449_/Y vdd gnd AOI21X1
XFILL_2__10903_ vdd gnd FILL
XFILL_1__12332_ vdd gnd FILL
X_13168_ _13168_/A _13168_/B _13168_/C _13168_/Y vdd gnd NAND3X1
XFILL_0__7560_ vdd gnd FILL
XFILL_2__13622_ vdd gnd FILL
XFILL_0__14801_ vdd gnd FILL
XFILL_2__10834_ vdd gnd FILL
XFILL_1__12263_ vdd gnd FILL
X_12119_ _12119_/A _12119_/B _12119_/C _12119_/Y vdd gnd OAI21X1
XFILL_0__12993_ vdd gnd FILL
XFILL_1__14002_ vdd gnd FILL
X_13099_ _13099_/A _13099_/B _13099_/C _13099_/Y vdd gnd OAI21X1
XFILL_0__7491_ vdd gnd FILL
XFILL_2__7427_ vdd gnd FILL
XFILL_1__11214_ vdd gnd FILL
XFILL_2__13553_ vdd gnd FILL
XFILL_0__14732_ vdd gnd FILL
XFILL_0__9230_ vdd gnd FILL
XFILL_0__11944_ vdd gnd FILL
XFILL_1__12194_ vdd gnd FILL
XFILL_2__7358_ vdd gnd FILL
XFILL_1__11145_ vdd gnd FILL
XFILL_0__14663_ vdd gnd FILL
XFILL_0__9161_ vdd gnd FILL
XFILL_0__11875_ vdd gnd FILL
XFILL_0__13614_ vdd gnd FILL
XFILL_2__7289_ vdd gnd FILL
XFILL_1__11076_ vdd gnd FILL
XFILL_0__8112_ vdd gnd FILL
XFILL_0__10826_ vdd gnd FILL
XFILL_0__14594_ vdd gnd FILL
XFILL_0__9092_ vdd gnd FILL
X_8740_ _8740_/A _8740_/B _8740_/C _8740_/D _8740_/Y vdd gnd OAI22X1
XFILL_1__10027_ vdd gnd FILL
XFILL_0__13545_ vdd gnd FILL
XFILL256950x230550 vdd gnd FILL
XFILL_0__8043_ vdd gnd FILL
X_8671_ _8671_/A _8671_/B _8671_/C _8671_/Y vdd gnd OAI21X1
XFILL_1__14835_ vdd gnd FILL
X_7622_ _7622_/A _7622_/Y vdd gnd INVX1
XFILL_2__11248_ vdd gnd FILL
XFILL_1__14766_ vdd gnd FILL
XFILL_0__12427_ vdd gnd FILL
XFILL_1__11978_ vdd gnd FILL
X_7553_ _7553_/A _7553_/B _7553_/Y vdd gnd NAND2X1
XFILL_0__9994_ vdd gnd FILL
XFILL_1__13717_ vdd gnd FILL
XFILL_2__11179_ vdd gnd FILL
XFILL_1__10929_ vdd gnd FILL
XFILL_1__14697_ vdd gnd FILL
XFILL_0__12358_ vdd gnd FILL
XFILL_0__8945_ vdd gnd FILL
X_7484_ _7484_/A _7484_/B _7484_/C _7484_/Y vdd gnd OAI21X1
XFILL_1__13648_ vdd gnd FILL
XFILL_0__11309_ vdd gnd FILL
X_9223_ _9223_/A _9223_/B _9223_/C _9223_/Y vdd gnd OAI21X1
XFILL_0__12289_ vdd gnd FILL
XFILL_0__14028_ vdd gnd FILL
XFILL_1__13579_ vdd gnd FILL
X_9154_ _9154_/A _9154_/Y vdd gnd INVX1
XFILL_0__7827_ vdd gnd FILL
X_8105_ _8105_/A _8105_/B _8105_/C _8105_/Y vdd gnd OAI21X1
X_9085_ _9085_/A _9085_/Y vdd gnd INVX1
XFILL_0__7758_ vdd gnd FILL
XFILL_1__9270_ vdd gnd FILL
X_8036_ _8036_/A _8036_/B _8036_/C _8036_/D _8036_/Y vdd gnd AOI22X1
XFILL_0__7689_ vdd gnd FILL
XFILL_1__8221_ vdd gnd FILL
XFILL_0__9428_ vdd gnd FILL
XFILL_1__8152_ vdd gnd FILL
XFILL_0__9359_ vdd gnd FILL
X_9987_ _9987_/A _9987_/B _9987_/C _9987_/Y vdd gnd AOI21X1
XFILL_1__7103_ vdd gnd FILL
X_8938_ _8938_/A _8938_/Y vdd gnd INVX1
XFILL_1__8083_ vdd gnd FILL
XFILL256950x140550 vdd gnd FILL
X_8869_ _8869_/D _8869_/CLK _8869_/Q vdd gnd DFFPOSX1
X_12470_ _12470_/A _12470_/B _12470_/C _12470_/Y vdd gnd OAI21X1
XFILL_1__8985_ vdd gnd FILL
X_11421_ _11421_/A _11421_/B _11421_/Y vdd gnd NOR2X1
X_14140_ _14140_/A _14140_/B _14140_/C _14140_/Y vdd gnd OAI21X1
X_11352_ _11352_/A _11352_/B _11352_/C _11352_/Y vdd gnd AOI21X1
XFILL_1__7867_ vdd gnd FILL
X_10303_ _10303_/A _10303_/B _10303_/C _10303_/Y vdd gnd OAI21X1
X_14071_ _14071_/A _14071_/B _14071_/Y vdd gnd NOR2X1
XFILL_1__9606_ vdd gnd FILL
X_11283_ _11283_/A _11283_/B _11283_/C _11283_/Y vdd gnd OAI21X1
XFILL_1__7798_ vdd gnd FILL
X_13022_ _13022_/A _13022_/B _13022_/Y vdd gnd NAND2X1
X_10234_ _10234_/A _10234_/B _10234_/C _10234_/Y vdd gnd OAI21X1
XFILL_1__9537_ vdd gnd FILL
X_10165_ _10165_/A _10165_/B _10165_/C _10165_/Y vdd gnd OAI21X1
XFILL_1__9468_ vdd gnd FILL
XFILL_2__7212_ vdd gnd FILL
X_10096_ _10096_/A _10096_/B _10096_/C _10096_/Y vdd gnd NAND3X1
XFILL_1__8419_ vdd gnd FILL
XFILL_1__9399_ vdd gnd FILL
X_13924_ _13924_/A _13924_/B _13924_/Y vdd gnd NAND2X1
XFILL_2__7143_ vdd gnd FILL
X_13855_ _13855_/A _13855_/B _13855_/C _13855_/D _13855_/Y vdd gnd AOI22X1
XFILL_2__12220_ vdd gnd FILL
XFILL_2__7074_ vdd gnd FILL
XFILL_1__12950_ vdd gnd FILL
XFILL_0__10611_ vdd gnd FILL
XFILL_1_BUFX2_insert220 vdd gnd FILL
XFILL_0__11591_ vdd gnd FILL
X_12806_ _12806_/A _12806_/B _12806_/Y vdd gnd NOR2X1
XFILL_1_BUFX2_insert231 vdd gnd FILL
X_10998_ _10998_/A _10998_/B _10998_/C _10998_/Y vdd gnd AOI21X1
XFILL_1__11901_ vdd gnd FILL
XFILL_2__12151_ vdd gnd FILL
XFILL_1_BUFX2_insert242 vdd gnd FILL
X_13786_ _13786_/A _13786_/B _13786_/Y vdd gnd AND2X2
XFILL_1_BUFX2_insert253 vdd gnd FILL
XFILL_0__13330_ vdd gnd FILL
XFILL_0__10542_ vdd gnd FILL
XFILL_1__12881_ vdd gnd FILL
XFILL_1_BUFX2_insert264 vdd gnd FILL
XFILL_1_BUFX2_insert275 vdd gnd FILL
X_12737_ _12737_/A _12737_/B _12737_/C _12737_/Y vdd gnd OAI21X1
XCLKBUF1_insert35 CLKBUF1_insert35/A CLKBUF1_insert35/Y vdd gnd CLKBUF1
XFILL_1__14620_ vdd gnd FILL
XFILL_1_BUFX2_insert286 vdd gnd FILL
XCLKBUF1_insert46 CLKBUF1_insert46/A CLKBUF1_insert46/Y vdd gnd CLKBUF1
XFILL_1__11832_ vdd gnd FILL
XFILL_1_BUFX2_insert297 vdd gnd FILL
XCLKBUF1_insert57 CLKBUF1_insert57/A CLKBUF1_insert57/Y vdd gnd CLKBUF1
XFILL_0__13261_ vdd gnd FILL
XFILL_0__10473_ vdd gnd FILL
XCLKBUF1_insert68 CLKBUF1_insert68/A CLKBUF1_insert68/Y vdd gnd CLKBUF1
XCLKBUF1_insert79 CLKBUF1_insert79/A CLKBUF1_insert79/Y vdd gnd CLKBUF1
X_12668_ _12668_/A _12668_/Y vdd gnd INVX1
XFILL_0__12212_ vdd gnd FILL
XFILL_1__11763_ vdd gnd FILL
XFILL_0__13192_ vdd gnd FILL
XFILL_0_CLKBUF1_insert390 vdd gnd FILL
X_14407_ _14407_/A _14407_/B _14407_/C _14407_/Y vdd gnd OAI21X1
X_11619_ _11619_/D _11619_/CLK _11619_/Q vdd gnd DFFPOSX1
XFILL_2__9715_ vdd gnd FILL
XFILL_1__13502_ vdd gnd FILL
X_12599_ _12599_/D _12599_/CLK _12599_/Q vdd gnd DFFPOSX1
XFILL_1__14482_ vdd gnd FILL
XFILL_0__12143_ vdd gnd FILL
XFILL_1__11694_ vdd gnd FILL
XFILL_0__8730_ vdd gnd FILL
X_14338_ _14338_/A _14338_/B _14338_/Y vdd gnd NAND2X1
XFILL_2__9646_ vdd gnd FILL
XFILL_1__10645_ vdd gnd FILL
XFILL_0__12074_ vdd gnd FILL
XFILL_2__12984_ vdd gnd FILL
X_14269_ _14269_/A _14269_/B _14269_/Y vdd gnd NAND2X1
XFILL_0__8661_ vdd gnd FILL
XFILL_0__11025_ vdd gnd FILL
XFILL_2__9577_ vdd gnd FILL
XFILL_1__13364_ vdd gnd FILL
XFILL_1__10576_ vdd gnd FILL
XFILL_0__7612_ vdd gnd FILL
XFILL_0__8592_ vdd gnd FILL
XFILL_1__12315_ vdd gnd FILL
XFILL_1__13295_ vdd gnd FILL
XFILL_0__7543_ vdd gnd FILL
XFILL_1__12246_ vdd gnd FILL
XFILL_2__10817_ vdd gnd FILL
XFILL_0__12976_ vdd gnd FILL
XFILL_0__7474_ vdd gnd FILL
X_9910_ _9910_/A _9910_/B _9910_/Y vdd gnd NAND2X1
XFILL_0__14715_ vdd gnd FILL
XFILL_0__11927_ vdd gnd FILL
XFILL_1__12177_ vdd gnd FILL
XFILL_0__9213_ vdd gnd FILL
X_9841_ _9841_/D _9841_/CLK _9841_/Q vdd gnd DFFPOSX1
XFILL_1__11128_ vdd gnd FILL
XFILL_0__14646_ vdd gnd FILL
XFILL_0__9144_ vdd gnd FILL
XFILL_0__11858_ vdd gnd FILL
X_9772_ _9772_/D _9772_/CLK _9772_/Q vdd gnd DFFPOSX1
XFILL_1__11059_ vdd gnd FILL
XFILL_2__13398_ vdd gnd FILL
XFILL_0__10809_ vdd gnd FILL
XFILL_0__14577_ vdd gnd FILL
XFILL_0__9075_ vdd gnd FILL
X_8723_ _8723_/A _8723_/B _8723_/C _8723_/Y vdd gnd AOI21X1
XFILL_0__11789_ vdd gnd FILL
XFILL_0__13528_ vdd gnd FILL
XFILL_0__8026_ vdd gnd FILL
X_8654_ _8654_/A _8654_/B _8654_/Y vdd gnd NAND2X1
XFILL_1__14818_ vdd gnd FILL
X_7605_ _7605_/A _7605_/B _7605_/C _7605_/Y vdd gnd NAND3X1
X_8585_ _8585_/A _8585_/Y vdd gnd INVX1
XFILL_1__14749_ vdd gnd FILL
X_7536_ _7536_/A _7536_/Y vdd gnd INVX1
XFILL_0__9977_ vdd gnd FILL
XFILL_1__8770_ vdd gnd FILL
XFILL_0__8928_ vdd gnd FILL
XFILL_1__7721_ vdd gnd FILL
X_7467_ _7467_/A _7467_/Y vdd gnd INVX1
X_9206_ _9206_/A _9206_/B _9206_/C _9206_/Y vdd gnd NAND3X1
XFILL_1__7652_ vdd gnd FILL
X_7398_ _7398_/A _7398_/B _7398_/C _7398_/Y vdd gnd NAND3X1
XFILL257550x100950 vdd gnd FILL
X_9137_ _9137_/A _9137_/Y vdd gnd INVX1
XFILL_1__7583_ vdd gnd FILL
XFILL_1__9322_ vdd gnd FILL
X_9068_ _9068_/A _9068_/B _9068_/C _9068_/Y vdd gnd AOI21X1
X_8019_ _8019_/A _8019_/B _8019_/Y vdd gnd NAND2X1
XFILL_1__9253_ vdd gnd FILL
XFILL_1__8204_ vdd gnd FILL
XFILL_1__9184_ vdd gnd FILL
X_11970_ _11970_/A _11970_/B _11970_/C _11970_/Y vdd gnd OAI21X1
XFILL_1__8135_ vdd gnd FILL
X_10921_ _10921_/A _10921_/Y vdd gnd INVX1
X_13640_ _13640_/A _13640_/B _13640_/C _13640_/Y vdd gnd OAI21X1
X_10852_ _10852_/A _10852_/B _10852_/C _10852_/Y vdd gnd OAI21X1
XFILL_1__8066_ vdd gnd FILL
X_10783_ _10783_/A _10783_/Y vdd gnd INVX1
X_13571_ _13571_/A _13571_/Y vdd gnd INVX4
XFILL_0_BUFX2_insert205 vdd gnd FILL
XFILL_0_BUFX2_insert216 vdd gnd FILL
X_12522_ _12522_/A _12522_/B _12522_/Y vdd gnd NAND2X1
XFILL_0_BUFX2_insert227 vdd gnd FILL
XFILL_2__7830_ vdd gnd FILL
XFILL_0_BUFX2_insert238 vdd gnd FILL
XFILL_0_BUFX2_insert249 vdd gnd FILL
X_12453_ _12453_/A _12453_/B _12453_/Y vdd gnd NAND2X1
XFILL_1__8968_ vdd gnd FILL
X_11404_ _11404_/A _11404_/Y vdd gnd INVX1
XFILL_2__9500_ vdd gnd FILL
X_12384_ _12384_/A _12384_/B _12384_/Y vdd gnd NAND2X1
X_11335_ _11335_/A _11335_/B _11335_/Y vdd gnd NAND2X1
X_14123_ _14123_/A _14123_/B _14123_/C _14123_/Y vdd gnd OAI21X1
XFILL_2__9431_ vdd gnd FILL
XFILL_1__10430_ vdd gnd FILL
X_14054_ _14054_/A _14054_/B _14054_/Y vdd gnd NOR2X1
X_11266_ _11266_/A _11266_/B _11266_/C _11266_/Y vdd gnd OAI21X1
XFILL_2__9362_ vdd gnd FILL
XFILL_1__10361_ vdd gnd FILL
X_10217_ _10217_/A _10217_/B _10217_/Y vdd gnd NAND2X1
X_13005_ _13005_/A _13005_/B _13005_/Y vdd gnd NAND2X1
XFILL_1__12100_ vdd gnd FILL
X_11197_ _11197_/A _11197_/Y vdd gnd INVX1
XFILL_1__13080_ vdd gnd FILL
XFILL_2__9293_ vdd gnd FILL
XFILL_0__12830_ vdd gnd FILL
XFILL_1__10292_ vdd gnd FILL
X_10148_ _10148_/A _10148_/Y vdd gnd INVX1
XFILL_1__12031_ vdd gnd FILL
XFILL_2__11582_ vdd gnd FILL
XFILL_0__12761_ vdd gnd FILL
X_10079_ _10079_/A _10079_/B _10079_/C _10079_/Y vdd gnd OAI21X1
XFILL_0__11712_ vdd gnd FILL
X_13907_ _13907_/A _13907_/B _13907_/Y vdd gnd NAND2X1
XFILL_0__12692_ vdd gnd FILL
XFILL_0__7190_ vdd gnd FILL
X_14887_ _14887_/D _14887_/CLK _14887_/Q vdd gnd DFFPOSX1
XFILL_0__14431_ vdd gnd FILL
XFILL_1__13982_ vdd gnd FILL
XFILL_2__12203_ vdd gnd FILL
X_13838_ _13838_/A _13838_/Y vdd gnd INVX1
XFILL_1__12933_ vdd gnd FILL
XFILL_0__14362_ vdd gnd FILL
XFILL_0__11574_ vdd gnd FILL
XFILL_2__12134_ vdd gnd FILL
X_13769_ _13769_/A _13769_/Y vdd gnd INVX1
XFILL_0__13313_ vdd gnd FILL
XFILL_0__10525_ vdd gnd FILL
XFILL_1__12864_ vdd gnd FILL
XFILL_0__9900_ vdd gnd FILL
XFILL_0__14293_ vdd gnd FILL
XFILL_1__14603_ vdd gnd FILL
XFILL_1__11815_ vdd gnd FILL
XFILL_2__12065_ vdd gnd FILL
XFILL_0__13244_ vdd gnd FILL
XFILL_0__10456_ vdd gnd FILL
XFILL_1__12795_ vdd gnd FILL
X_8370_ _8370_/A _8370_/B _8370_/C _8370_/Y vdd gnd OAI21X1
XFILL_1__11746_ vdd gnd FILL
XFILL_0__13175_ vdd gnd FILL
X_7321_ _7321_/A _7321_/Y vdd gnd INVX1
XFILL_0__10387_ vdd gnd FILL
XFILL_0__9762_ vdd gnd FILL
XFILL_1__14465_ vdd gnd FILL
XFILL_0__12126_ vdd gnd FILL
XFILL_0__8713_ vdd gnd FILL
X_7252_ _7252_/A _7252_/Y vdd gnd INVX1
XFILL_0__9693_ vdd gnd FILL
XFILL_2__9629_ vdd gnd FILL
XFILL_1__13416_ vdd gnd FILL
XFILL_1__10628_ vdd gnd FILL
XFILL_2__12967_ vdd gnd FILL
XFILL_1__14396_ vdd gnd FILL
XFILL_0__12057_ vdd gnd FILL
XFILL_0__8644_ vdd gnd FILL
X_7183_ _7183_/A _7183_/B _7183_/Y vdd gnd NAND2X1
XFILL_0__11008_ vdd gnd FILL
XFILL_1__13347_ vdd gnd FILL
XFILL_1__10559_ vdd gnd FILL
XFILL_2__12898_ vdd gnd FILL
XFILL_0__8575_ vdd gnd FILL
XFILL_1__13278_ vdd gnd FILL
XFILL_0__7526_ vdd gnd FILL
XFILL_1__12229_ vdd gnd FILL
XFILL_1_BUFX2_insert6 vdd gnd FILL
XFILL_0__12959_ vdd gnd FILL
XFILL_0__7457_ vdd gnd FILL
XFILL_2__14499_ vdd gnd FILL
XFILL_0__7388_ vdd gnd FILL
X_9824_ _9824_/D _9824_/CLK _9824_/Q vdd gnd DFFPOSX1
XFILL_0__14629_ vdd gnd FILL
XFILL_0__9127_ vdd gnd FILL
X_9755_ _9755_/A _9755_/B _9755_/C _9755_/Y vdd gnd OAI21X1
XFILL_0__9058_ vdd gnd FILL
XFILL_1__9940_ vdd gnd FILL
X_8706_ _8706_/A _8706_/B _8706_/Y vdd gnd NAND2X1
X_9686_ _9686_/A _9686_/B _9686_/C _9686_/Y vdd gnd OAI21X1
XFILL_0__8009_ vdd gnd FILL
X_8637_ _8637_/A _8637_/B _8637_/Y vdd gnd NAND2X1
XFILL_1__9871_ vdd gnd FILL
XFILL_1__8822_ vdd gnd FILL
X_8568_ _8568_/A _8568_/B _8568_/C _8568_/Y vdd gnd OAI21X1
X_7519_ _7519_/A _7519_/B _7519_/Y vdd gnd OR2X2
XFILL_1__8753_ vdd gnd FILL
X_8499_ _8499_/A _8499_/B _8499_/Y vdd gnd NAND2X1
XFILL_1__7704_ vdd gnd FILL
XFILL_1__8684_ vdd gnd FILL
X_11120_ _11120_/A _11120_/Y vdd gnd INVX1
XFILL_1__7635_ vdd gnd FILL
X_11051_ _11051_/A _11051_/Y vdd gnd INVX1
XFILL_1__7566_ vdd gnd FILL
X_10002_ _10002_/A _10002_/B _10002_/C _10002_/Y vdd gnd OAI21X1
XFILL_1__9305_ vdd gnd FILL
XFILL_1__7497_ vdd gnd FILL
X_14810_ _14810_/A _14810_/B _14810_/Y vdd gnd AND2X2
XFILL_1__9236_ vdd gnd FILL
X_14741_ _14741_/A _14741_/B _14741_/C _14741_/Y vdd gnd OAI21X1
X_11953_ _11953_/A _11953_/B _11953_/C _11953_/Y vdd gnd OAI21X1
XFILL_1__9167_ vdd gnd FILL
X_10904_ _10904_/A _10904_/B _10904_/C _10904_/Y vdd gnd AOI21X1
X_14672_ _14672_/A _14672_/B _14672_/C _14672_/Y vdd gnd OAI21X1
XFILL_1__8118_ vdd gnd FILL
X_11884_ _11884_/A _11884_/B _11884_/Y vdd gnd NAND2X1
XFILL_1__9098_ vdd gnd FILL
X_13623_ _13623_/A _13623_/B _13623_/S _13623_/Y vdd gnd MUX2X1
X_10835_ _10835_/A _10835_/B _10835_/C _10835_/Y vdd gnd OAI21X1
XFILL_2__8931_ vdd gnd FILL
XFILL_1__8049_ vdd gnd FILL
X_13554_ _13554_/A _13554_/B _13554_/S _13554_/Y vdd gnd MUX2X1
X_10766_ _10766_/D _10766_/CLK _10766_/Q vdd gnd DFFPOSX1
XFILL_0__10310_ vdd gnd FILL
X_12505_ _12505_/A _12505_/B _12505_/C _12505_/Y vdd gnd OAI21X1
XFILL_0__11290_ vdd gnd FILL
XFILL_2__7813_ vdd gnd FILL
X_10697_ _10697_/D _10697_/CLK _10697_/Q vdd gnd DFFPOSX1
XFILL_1__11600_ vdd gnd FILL
X_13485_ _13485_/D _13485_/CLK _13485_/Q vdd gnd DFFPOSX1
XFILL_0__10241_ vdd gnd FILL
X_12436_ _12436_/A _12436_/B _12436_/C _12436_/D _12436_/Y vdd gnd OAI22X1
XFILL_2__7744_ vdd gnd FILL
XFILL_1__11531_ vdd gnd FILL
XFILL_2__13870_ vdd gnd FILL
XFILL_0__10172_ vdd gnd FILL
X_12367_ _12367_/A _12367_/B _12367_/C _12367_/Y vdd gnd OAI21X1
XFILL_1__14250_ vdd gnd FILL
XFILL_2__7675_ vdd gnd FILL
XFILL_1__11462_ vdd gnd FILL
X_14106_ _14106_/A _14106_/Y vdd gnd INVX1
X_11318_ _11318_/A _11318_/Y vdd gnd INVX1
XFILL_1__13201_ vdd gnd FILL
X_12298_ _12298_/A _12298_/B _12298_/Y vdd gnd NAND2X1
XFILL_1__10413_ vdd gnd FILL
XFILL_0__13931_ vdd gnd FILL
XFILL_2__12752_ vdd gnd FILL
XFILL_1__11393_ vdd gnd FILL
X_11249_ _11249_/A _11249_/B _11249_/Y vdd gnd NAND2X1
X_14037_ _14037_/A _14037_/B _14037_/C _14037_/Y vdd gnd NAND3X1
XFILL_1__13132_ vdd gnd FILL
XFILL_2__11703_ vdd gnd FILL
XFILL_1__10344_ vdd gnd FILL
XFILL_0__13862_ vdd gnd FILL
XFILL_2__12683_ vdd gnd FILL
XFILL_0__8360_ vdd gnd FILL
XFILL_2__9276_ vdd gnd FILL
XFILL_0__12813_ vdd gnd FILL
XFILL_1__13063_ vdd gnd FILL
XFILL_1__10275_ vdd gnd FILL
XFILL_0__7311_ vdd gnd FILL
XFILL_0__13793_ vdd gnd FILL
XFILL_0__8291_ vdd gnd FILL
XFILL_1__12014_ vdd gnd FILL
XFILL_2__11565_ vdd gnd FILL
XFILL_0__12744_ vdd gnd FILL
XFILL_0__7242_ vdd gnd FILL
X_7870_ _7870_/A _7870_/B _7870_/C _7870_/Y vdd gnd OAI21X1
XFILL_2__11496_ vdd gnd FILL
XFILL_0__12675_ vdd gnd FILL
XFILL_0__7173_ vdd gnd FILL
XFILL_0__14414_ vdd gnd FILL
XFILL_1__13965_ vdd gnd FILL
X_9540_ _9540_/A _9540_/B _9540_/C _9540_/Y vdd gnd OAI21X1
XFILL_0__14345_ vdd gnd FILL
XFILL_1__12916_ vdd gnd FILL
XFILL_0__11557_ vdd gnd FILL
XFILL_1__13896_ vdd gnd FILL
X_9471_ _9471_/A _9471_/B _9471_/C _9471_/Y vdd gnd NAND3X1
XFILL_2__12117_ vdd gnd FILL
XFILL_0__10508_ vdd gnd FILL
XFILL_0__14276_ vdd gnd FILL
XFILL_1__12847_ vdd gnd FILL
X_8422_ _8422_/A _8422_/B _8422_/C _8422_/Y vdd gnd AOI21X1
XFILL_0__11488_ vdd gnd FILL
XFILL_2__12048_ vdd gnd FILL
XFILL_0__13227_ vdd gnd FILL
XFILL_0__10439_ vdd gnd FILL
XFILL_1__12778_ vdd gnd FILL
X_8353_ _8353_/A _8353_/B _8353_/C _8353_/Y vdd gnd NOR3X1
XFILL_1__11729_ vdd gnd FILL
XFILL_0__13158_ vdd gnd FILL
X_7304_ _7304_/A _7304_/B _7304_/C _7304_/Y vdd gnd OAI21X1
XFILL_0__9745_ vdd gnd FILL
X_8284_ _8284_/A _8284_/Y vdd gnd INVX1
XFILL_0__12109_ vdd gnd FILL
XFILL_1__14448_ vdd gnd FILL
XFILL_0__13089_ vdd gnd FILL
XFILL_2__13999_ vdd gnd FILL
X_7235_ _7235_/A _7235_/Y vdd gnd INVX1
XFILL_0__9676_ vdd gnd FILL
XFILL_1__14379_ vdd gnd FILL
XFILL_1__7420_ vdd gnd FILL
XFILL_0__8627_ vdd gnd FILL
X_7166_ _7166_/A _7166_/B _7166_/C _7166_/Y vdd gnd NAND3X1
XFILL_1__7351_ vdd gnd FILL
XFILL_0__8558_ vdd gnd FILL
X_7097_ _7097_/A _7097_/B _7097_/C _7097_/Y vdd gnd OAI21X1
XFILL_2_BUFX2_insert108 vdd gnd FILL
XFILL_0__7509_ vdd gnd FILL
XFILL_1__7282_ vdd gnd FILL
XFILL_0__8489_ vdd gnd FILL
XFILL_1__9021_ vdd gnd FILL
X_9807_ _9807_/D _9807_/CLK _9807_/Q vdd gnd DFFPOSX1
X_7999_ _7999_/A _7999_/Y vdd gnd INVX2
X_9738_ _9738_/A _9738_/B _9738_/Y vdd gnd NAND2X1
X_10620_ _10620_/A _10620_/B _10620_/C _10620_/Y vdd gnd OAI21X1
XBUFX2_insert118 BUFX2_insert118/A BUFX2_insert118/Y vdd gnd BUFX2
XFILL_1__9923_ vdd gnd FILL
XBUFX2_insert129 BUFX2_insert129/A BUFX2_insert129/Y vdd gnd BUFX2
X_9669_ _9669_/A _9669_/B _9669_/C _9669_/Y vdd gnd AOI21X1
X_10551_ _10551_/A _10551_/B _10551_/Y vdd gnd NAND2X1
XFILL_1__9854_ vdd gnd FILL
X_10482_ _10482_/A _10482_/B _10482_/C _10482_/Y vdd gnd OAI21X1
XFILL_1__8805_ vdd gnd FILL
X_13270_ _13270_/A _13270_/B _13270_/Y vdd gnd NAND2X1
X_12221_ _12221_/A _12221_/B _12221_/Y vdd gnd NAND2X1
XFILL_1__8736_ vdd gnd FILL
X_12152_ _12152_/A _12152_/B _12152_/Y vdd gnd NAND2X1
XFILL_2__7460_ vdd gnd FILL
XFILL_1__8667_ vdd gnd FILL
X_11103_ _11103_/A _11103_/B _11103_/Y vdd gnd NAND2X1
X_12083_ _12083_/A _12083_/B _12083_/S _12083_/Y vdd gnd MUX2X1
XFILL_1__7618_ vdd gnd FILL
XFILL_2__7391_ vdd gnd FILL
XFILL_1__8598_ vdd gnd FILL
X_11034_ _11034_/A _11034_/B _11034_/C _11034_/Y vdd gnd NAND3X1
XFILL_1__7549_ vdd gnd FILL
XFILL_1__10060_ vdd gnd FILL
XFILL_0__10790_ vdd gnd FILL
XFILL_1__9219_ vdd gnd FILL
XFILL_2__8012_ vdd gnd FILL
X_12985_ _12985_/A _12985_/B _12985_/Y vdd gnd NAND2X1
X_14724_ _14724_/A _14724_/B _14724_/Y vdd gnd NAND2X1
XFILL_2__10301_ vdd gnd FILL
X_11936_ _11936_/A _11936_/B _11936_/C _11936_/Y vdd gnd OAI21X1
XFILL_0__12460_ vdd gnd FILL
X_14655_ _14655_/A _14655_/B _14655_/C _14655_/Y vdd gnd OAI21X1
XFILL_2__10232_ vdd gnd FILL
X_11867_ _11867_/A _11867_/Y vdd gnd INVX1
XFILL_0__11411_ vdd gnd FILL
XFILL_1__10962_ vdd gnd FILL
XFILL_1__13750_ vdd gnd FILL
XFILL_0__12391_ vdd gnd FILL
X_13606_ _13606_/A _13606_/B _13606_/S _13606_/Y vdd gnd MUX2X1
X_10818_ _10818_/A _10818_/B _10818_/Y vdd gnd NAND2X1
X_14586_ _14586_/A _14586_/B _14586_/Y vdd gnd NAND2X1
XFILL_2__10163_ vdd gnd FILL
X_11798_ _11798_/A _11798_/B _11798_/S _11798_/Y vdd gnd MUX2X1
XFILL_1__12701_ vdd gnd FILL
XFILL_0__14130_ vdd gnd FILL
XFILL_0__11342_ vdd gnd FILL
XFILL_1__13681_ vdd gnd FILL
XFILL_1__10893_ vdd gnd FILL
X_13537_ _13537_/A _13537_/Y vdd gnd INVX1
X_10749_ _10749_/D _10749_/CLK _10749_/Q vdd gnd DFFPOSX1
XFILL_1__12632_ vdd gnd FILL
XFILL_2__10094_ vdd gnd FILL
XFILL_0__14061_ vdd gnd FILL
XFILL_0__11273_ vdd gnd FILL
XFILL_0__7860_ vdd gnd FILL
X_13468_ _13468_/D _13468_/CLK _13468_/Q vdd gnd DFFPOSX1
XFILL_0__13012_ vdd gnd FILL
XFILL_0__10224_ vdd gnd FILL
X_12419_ _12419_/A _12419_/B _12419_/C _12419_/Y vdd gnd AOI21X1
XFILL_2__7727_ vdd gnd FILL
XFILL_0__7791_ vdd gnd FILL
XFILL_1__14302_ vdd gnd FILL
XFILL_1__11514_ vdd gnd FILL
X_13399_ _13399_/A _13399_/B _13399_/C _13399_/Y vdd gnd OAI21X1
XFILL_0__10155_ vdd gnd FILL
XFILL_1__12494_ vdd gnd FILL
XFILL_0__9530_ vdd gnd FILL
XFILL_1__14233_ vdd gnd FILL
XFILL_2__7658_ vdd gnd FILL
XFILL_1__11445_ vdd gnd FILL
XFILL_2__13784_ vdd gnd FILL
XFILL_2__10996_ vdd gnd FILL
XFILL_0__10086_ vdd gnd FILL
XFILL_0__9461_ vdd gnd FILL
XFILL_0__13914_ vdd gnd FILL
XFILL_2__7589_ vdd gnd FILL
XFILL_1__11376_ vdd gnd FILL
XFILL_0__8412_ vdd gnd FILL
XFILL_1__13115_ vdd gnd FILL
XFILL_0__9392_ vdd gnd FILL
XFILL_1__10327_ vdd gnd FILL
XFILL_1__14095_ vdd gnd FILL
XFILL_0__13845_ vdd gnd FILL
XFILL_0__8343_ vdd gnd FILL
X_8971_ _8971_/A _8971_/Y vdd gnd INVX1
XFILL257250x226950 vdd gnd FILL
XFILL_1__13046_ vdd gnd FILL
XFILL_1__10258_ vdd gnd FILL
XFILL_0__13776_ vdd gnd FILL
XFILL_0__10988_ vdd gnd FILL
X_7922_ _7922_/D _7922_/CLK _7922_/Q vdd gnd DFFPOSX1
XFILL_0__8274_ vdd gnd FILL
XFILL_0__12727_ vdd gnd FILL
XFILL_1__10189_ vdd gnd FILL
XFILL_0__7225_ vdd gnd FILL
X_7853_ _7853_/A _7853_/B _7853_/C _7853_/Y vdd gnd OAI21X1
XFILL_0__12658_ vdd gnd FILL
XFILL_0__7156_ vdd gnd FILL
X_7784_ _7784_/A _7784_/B _7784_/Y vdd gnd NAND2X1
XFILL_0__11609_ vdd gnd FILL
XFILL_1__13948_ vdd gnd FILL
X_9523_ _9523_/A _9523_/B _9523_/Y vdd gnd NAND2X1
XFILL_0__7087_ vdd gnd FILL
XFILL_0__14328_ vdd gnd FILL
XFILL_1__13879_ vdd gnd FILL
X_9454_ _9454_/A _9454_/Y vdd gnd INVX1
XFILL_0__14259_ vdd gnd FILL
X_8405_ _8405_/A _8405_/B _8405_/Y vdd gnd NAND2X1
X_9385_ _9385_/A _9385_/B _9385_/C _9385_/Y vdd gnd NAND3X1
X_8336_ _8336_/A _8336_/B _8336_/Y vdd gnd AND2X2
XFILL_1__9570_ vdd gnd FILL
XFILL256650x108150 vdd gnd FILL
XFILL_0__9728_ vdd gnd FILL
XFILL_1__8521_ vdd gnd FILL
X_8267_ _8267_/A _8267_/Y vdd gnd INVX1
X_7218_ _7218_/A _7218_/B _7218_/C _7218_/Y vdd gnd OAI21X1
XFILL_0__9659_ vdd gnd FILL
XFILL_1__8452_ vdd gnd FILL
X_8198_ _8198_/A _8198_/B _8198_/C _8198_/Y vdd gnd OAI21X1
XFILL_1__7403_ vdd gnd FILL
X_7149_ _7149_/A _7149_/B _7149_/Y vdd gnd NOR2X1
XFILL_1__8383_ vdd gnd FILL
XFILL_1__7334_ vdd gnd FILL
XFILL257250x136950 vdd gnd FILL
XFILL_1__7265_ vdd gnd FILL
XFILL_1__9004_ vdd gnd FILL
X_12770_ _12770_/A _12770_/B _12770_/C _12770_/Y vdd gnd OAI21X1
XFILL_1__7196_ vdd gnd FILL
X_11721_ _11721_/A _11721_/B _11721_/C _11721_/Y vdd gnd OAI21X1
X_14440_ _14440_/A _14440_/B _14440_/Y vdd gnd NAND2X1
X_11652_ _11652_/D _11652_/CLK _11652_/Q vdd gnd DFFPOSX1
X_10603_ _10603_/A _10603_/B _10603_/C _10603_/Y vdd gnd OAI21X1
XFILL_1__9906_ vdd gnd FILL
X_14371_ _14371_/A _14371_/B _14371_/Y vdd gnd NAND2X1
X_11583_ _11583_/A _11583_/B _11583_/C _11583_/Y vdd gnd OAI21X1
X_13322_ _13322_/A _13322_/B _13322_/Y vdd gnd NOR2X1
X_10534_ _10534_/A _10534_/B _10534_/Y vdd gnd NAND2X1
X_10465_ _10465_/A _10465_/B _10465_/Y vdd gnd NAND2X1
X_13253_ _13253_/A _13253_/Y vdd gnd INVX1
X_12204_ _12204_/A _12204_/B _12204_/Y vdd gnd NAND2X1
X_13184_ _13184_/A _13184_/B _13184_/C _13184_/Y vdd gnd NAND3X1
X_10396_ _10396_/A _10396_/Y vdd gnd INVX1
XFILL_1__8719_ vdd gnd FILL
XFILL_1__9699_ vdd gnd FILL
XFILL_2__10850_ vdd gnd FILL
X_12135_ _12135_/A _12135_/B _12135_/Y vdd gnd NAND2X1
XFILL_1__11230_ vdd gnd FILL
XFILL_2__7443_ vdd gnd FILL
XFILL_2__10781_ vdd gnd FILL
XFILL_0__11960_ vdd gnd FILL
X_12066_ _12066_/A _12066_/B _12066_/C _12066_/Y vdd gnd OAI21X1
XFILL_2__12520_ vdd gnd FILL
XFILL_1__11161_ vdd gnd FILL
XFILL_2__7374_ vdd gnd FILL
XFILL_0__10911_ vdd gnd FILL
XFILL_0__11891_ vdd gnd FILL
X_11017_ _11017_/A _11017_/Y vdd gnd INVX1
XFILL_1__10112_ vdd gnd FILL
XFILL_0__13630_ vdd gnd FILL
XFILL_2__12451_ vdd gnd FILL
XFILL_1__11092_ vdd gnd FILL
XFILL_0__10842_ vdd gnd FILL
XFILL_1__14920_ vdd gnd FILL
XFILL_1__10043_ vdd gnd FILL
XFILL_2__12382_ vdd gnd FILL
XBUFX2_insert7 BUFX2_insert7/A BUFX2_insert7/Y vdd gnd BUFX2
XFILL_0__13561_ vdd gnd FILL
XFILL_0__10773_ vdd gnd FILL
X_12968_ _12968_/A _12968_/B _12968_/C _12968_/Y vdd gnd OAI21X1
XFILL_2__14121_ vdd gnd FILL
XFILL_0__12512_ vdd gnd FILL
XFILL_1__14851_ vdd gnd FILL
X_14707_ _14707_/A _14707_/B _14707_/Y vdd gnd NOR2X1
X_11919_ _11919_/A _11919_/Y vdd gnd INVX1
XFILL_1__13802_ vdd gnd FILL
X_12899_ _12899_/A _12899_/B _12899_/C _12899_/Y vdd gnd NAND3X1
XFILL_0__12443_ vdd gnd FILL
XFILL_1__14782_ vdd gnd FILL
XFILL_1__11994_ vdd gnd FILL
X_14638_ _14638_/A _14638_/B _14638_/Y vdd gnd AND2X2
XFILL_2__10215_ vdd gnd FILL
XFILL_2__13003_ vdd gnd FILL
XFILL_1__13733_ vdd gnd FILL
XFILL_0__12374_ vdd gnd FILL
XFILL_1__10945_ vdd gnd FILL
XFILL_0__8961_ vdd gnd FILL
X_14569_ _14569_/A _14569_/B _14569_/Y vdd gnd NAND2X1
XFILL_2__10146_ vdd gnd FILL
XFILL_0__14113_ vdd gnd FILL
XFILL_0__11325_ vdd gnd FILL
XFILL_1__13664_ vdd gnd FILL
XFILL_1__10876_ vdd gnd FILL
XFILL_0__7912_ vdd gnd FILL
XFILL257250x201750 vdd gnd FILL
XFILL_2__10077_ vdd gnd FILL
XFILL_0__14044_ vdd gnd FILL
XFILL_1__13595_ vdd gnd FILL
XFILL_0__11256_ vdd gnd FILL
XFILL_0__7843_ vdd gnd FILL
X_9170_ _9170_/A _9170_/B _9170_/C _9170_/Y vdd gnd AOI21X1
XFILL_0__10207_ vdd gnd FILL
XFILL_0__11187_ vdd gnd FILL
X_8121_ _8121_/A _8121_/Y vdd gnd INVX1
XFILL_0__7774_ vdd gnd FILL
XFILL_0__10138_ vdd gnd FILL
XFILL_1__12477_ vdd gnd FILL
XFILL_0__9513_ vdd gnd FILL
X_8052_ _8052_/A _8052_/B _8052_/C _8052_/D _8052_/Y vdd gnd AOI22X1
XFILL_1__14216_ vdd gnd FILL
XFILL_1__11428_ vdd gnd FILL
XFILL_2__10979_ vdd gnd FILL
XFILL_1_BUFX2_insert11 vdd gnd FILL
XFILL_0__10069_ vdd gnd FILL
XFILL_0__9444_ vdd gnd FILL
XFILL_1_BUFX2_insert22 vdd gnd FILL
XFILL_1__11359_ vdd gnd FILL
XFILL_1__14147_ vdd gnd FILL
XFILL_0__9375_ vdd gnd FILL
XFILL_1__14078_ vdd gnd FILL
XFILL_0__13828_ vdd gnd FILL
XFILL_0__8326_ vdd gnd FILL
X_8954_ _8954_/A _8954_/B _8954_/C _8954_/Y vdd gnd OAI21X1
XFILL_1__13029_ vdd gnd FILL
XFILL_0__13759_ vdd gnd FILL
X_7905_ _7905_/A _7905_/B _7905_/C _7905_/Y vdd gnd OAI21X1
XFILL_0__8257_ vdd gnd FILL
X_8885_ _8885_/D _8885_/CLK _8885_/Q vdd gnd DFFPOSX1
XFILL_0__7208_ vdd gnd FILL
X_7836_ _7836_/A _7836_/B _7836_/C _7836_/Y vdd gnd OAI21X1
XFILL_0__8188_ vdd gnd FILL
XFILL_1_CLKBUF1_insert34 vdd gnd FILL
XFILL_1_CLKBUF1_insert45 vdd gnd FILL
XFILL_0__7139_ vdd gnd FILL
XFILL_1_CLKBUF1_insert56 vdd gnd FILL
XFILL_1_CLKBUF1_insert67 vdd gnd FILL
X_7767_ _7767_/A _7767_/B _7767_/C _7767_/Y vdd gnd OAI21X1
XFILL_1_CLKBUF1_insert78 vdd gnd FILL
XFILL_1_CLKBUF1_insert89 vdd gnd FILL
X_9506_ _9506_/A _9506_/B _9506_/C _9506_/Y vdd gnd NAND3X1
X_7698_ _7698_/A _7698_/B _7698_/C _7698_/Y vdd gnd OAI21X1
X_9437_ _9437_/A _9437_/B _9437_/Y vdd gnd NOR2X1
XFILL257250x111750 vdd gnd FILL
XFILL_1__7883_ vdd gnd FILL
XFILL_1__9622_ vdd gnd FILL
X_9368_ _9368_/A _9368_/B _9368_/C _9368_/Y vdd gnd OAI21X1
X_10250_ _10250_/A _10250_/Y vdd gnd INVX1
XFILL_1__9553_ vdd gnd FILL
X_8319_ _8319_/A _8319_/B _8319_/C _8319_/Y vdd gnd OAI21X1
X_9299_ _9299_/A _9299_/B _9299_/Y vdd gnd NAND2X1
X_10181_ _10181_/A _10181_/B _10181_/C _10181_/Y vdd gnd AOI21X1
XFILL_1__8504_ vdd gnd FILL
XFILL_1__9484_ vdd gnd FILL
XFILL_1__8435_ vdd gnd FILL
X_13940_ _13940_/A _13940_/B _13940_/Y vdd gnd NAND2X1
XFILL_1__8366_ vdd gnd FILL
XFILL_1__7317_ vdd gnd FILL
X_13871_ _13871_/A _13871_/B _13871_/Y vdd gnd NAND2X1
XFILL_1__8297_ vdd gnd FILL
X_12822_ _12822_/A _12822_/B _12822_/Y vdd gnd NAND2X1
XFILL_1__7248_ vdd gnd FILL
X_12753_ _12753_/A _12753_/B _12753_/Y vdd gnd NAND2X1
XFILL_1__7179_ vdd gnd FILL
X_11704_ _11704_/A _11704_/B _11704_/Y vdd gnd NOR2X1
X_12684_ _12684_/A _12684_/B _12684_/S _12684_/Y vdd gnd MUX2X1
X_14423_ _14423_/A _14423_/B _14423_/Y vdd gnd NAND2X1
X_11635_ _11635_/D _11635_/CLK _11635_/Q vdd gnd DFFPOSX1
X_14354_ _14354_/A _14354_/B _14354_/C _14354_/Y vdd gnd NAND3X1
X_11566_ _11566_/A _11566_/B _11566_/C _11566_/Y vdd gnd OAI21X1
XFILL_2__9662_ vdd gnd FILL
XFILL_0__11110_ vdd gnd FILL
XFILL_1__10661_ vdd gnd FILL
XFILL_0__12090_ vdd gnd FILL
X_13305_ _13305_/A _13305_/B _13305_/Y vdd gnd NAND2X1
X_10517_ _10517_/A _10517_/B _10517_/Y vdd gnd AND2X2
X_14285_ _14285_/A _14285_/B _14285_/C _14285_/Y vdd gnd OAI21X1
XFILL_2__8613_ vdd gnd FILL
XFILL_1__12400_ vdd gnd FILL
X_11497_ _11497_/A _11497_/B _11497_/C _11497_/Y vdd gnd OAI21X1
XFILL_0__11041_ vdd gnd FILL
XFILL_2__9593_ vdd gnd FILL
XFILL_1__13380_ vdd gnd FILL
XFILL_1__10592_ vdd gnd FILL
X_13236_ _13236_/A _13236_/B _13236_/Y vdd gnd NOR2X1
X_10448_ _10448_/A _10448_/Y vdd gnd INVX1
XFILL_1__12331_ vdd gnd FILL
XFILL_2__14670_ vdd gnd FILL
X_13167_ _13167_/A _13167_/B _13167_/C _13167_/Y vdd gnd AOI21X1
X_10379_ _10379_/A _10379_/B _10379_/C _10379_/Y vdd gnd OAI21X1
XFILL_0__14800_ vdd gnd FILL
XFILL_1__12262_ vdd gnd FILL
X_12118_ _12118_/A _12118_/B _12118_/C _12118_/Y vdd gnd AOI21X1
XFILL_0__12992_ vdd gnd FILL
XFILL_1__14001_ vdd gnd FILL
XFILL_0__7490_ vdd gnd FILL
X_13098_ _13098_/A _13098_/B _13098_/C _13098_/Y vdd gnd NAND3X1
XFILL_1__11213_ vdd gnd FILL
XFILL_0__14731_ vdd gnd FILL
XFILL_0__11943_ vdd gnd FILL
XFILL_1__12193_ vdd gnd FILL
X_12049_ _12049_/A _12049_/B _12049_/C _12049_/Y vdd gnd NOR3X1
XFILL_2__12503_ vdd gnd FILL
XFILL_1__11144_ vdd gnd FILL
XFILL_0__14662_ vdd gnd FILL
XFILL_0__11874_ vdd gnd FILL
XFILL_0__9160_ vdd gnd FILL
XFILL_2__12434_ vdd gnd FILL
XFILL_0__13613_ vdd gnd FILL
XFILL_1__11075_ vdd gnd FILL
XFILL_0__10825_ vdd gnd FILL
XFILL_0__14593_ vdd gnd FILL
XFILL_0__8111_ vdd gnd FILL
XFILL_0__9091_ vdd gnd FILL
XFILL_1__10026_ vdd gnd FILL
XFILL_2__12365_ vdd gnd FILL
XFILL_2_BUFX2_insert291 vdd gnd FILL
XFILL_0__13544_ vdd gnd FILL
XFILL_0__8042_ vdd gnd FILL
X_8670_ _8670_/A _8670_/B _8670_/C _8670_/Y vdd gnd OAI21X1
XFILL_2__14104_ vdd gnd FILL
XFILL_1__14834_ vdd gnd FILL
XFILL_2__12296_ vdd gnd FILL
XFILL_0__10687_ vdd gnd FILL
X_7621_ _7621_/A _7621_/B _7621_/C _7621_/Y vdd gnd AOI21X1
XFILL_2__14035_ vdd gnd FILL
XFILL_0__12426_ vdd gnd FILL
XFILL_1__14765_ vdd gnd FILL
XFILL_1__11977_ vdd gnd FILL
X_7552_ _7552_/A _7552_/B _7552_/C _7552_/Y vdd gnd OAI21X1
XFILL_0__9993_ vdd gnd FILL
XFILL_1__13716_ vdd gnd FILL
XFILL_0__12357_ vdd gnd FILL
XFILL_1__10928_ vdd gnd FILL
XFILL_1__14696_ vdd gnd FILL
XFILL_0__8944_ vdd gnd FILL
X_7483_ _7483_/A _7483_/B _7483_/C _7483_/Y vdd gnd AOI21X1
XFILL_2__10129_ vdd gnd FILL
XBUFX2_insert290 BUFX2_insert290/A BUFX2_insert290/Y vdd gnd BUFX2
XFILL_0__11308_ vdd gnd FILL
XFILL_1__13647_ vdd gnd FILL
XFILL_0__12288_ vdd gnd FILL
XFILL_1__10859_ vdd gnd FILL
X_9222_ _9222_/A _9222_/B _9222_/C _9222_/Y vdd gnd NAND3X1
XFILL_0__14027_ vdd gnd FILL
XFILL_0__11239_ vdd gnd FILL
XFILL_1__13578_ vdd gnd FILL
X_9153_ _9153_/A _9153_/B _9153_/C _9153_/Y vdd gnd NAND3X1
XFILL_0__7826_ vdd gnd FILL
XFILL_1__12529_ vdd gnd FILL
X_8104_ _8104_/A _8104_/B _8104_/Y vdd gnd NAND2X1
X_9084_ _9084_/A _9084_/B _9084_/C _9084_/Y vdd gnd NAND3X1
XFILL_0__7757_ vdd gnd FILL
X_8035_ _8035_/A _8035_/B _8035_/C _8035_/Y vdd gnd OAI21X1
XFILL_0__7688_ vdd gnd FILL
XFILL_0__9427_ vdd gnd FILL
XFILL_1__8220_ vdd gnd FILL
XFILL_0__9358_ vdd gnd FILL
XFILL_1__8151_ vdd gnd FILL
X_9986_ _9986_/A _9986_/B _9986_/C _9986_/Y vdd gnd AOI21X1
XFILL_1__7102_ vdd gnd FILL
XFILL_0__8309_ vdd gnd FILL
XFILL_0__9289_ vdd gnd FILL
X_8937_ _8937_/A _8937_/B _8937_/C _8937_/Y vdd gnd AOI21X1
XFILL_1__8082_ vdd gnd FILL
X_8868_ _8868_/D _8868_/CLK _8868_/Q vdd gnd DFFPOSX1
X_7819_ _7819_/A _7819_/B _7819_/C _7819_/Y vdd gnd NAND3X1
X_8799_ _8799_/A _8799_/B _8799_/C _8799_/Y vdd gnd OAI21X1
XFILL_1__8984_ vdd gnd FILL
X_11420_ _11420_/A _11420_/Y vdd gnd INVX1
X_11351_ _11351_/A _11351_/Y vdd gnd INVX1
XFILL_1__7866_ vdd gnd FILL
X_10302_ _10302_/A _10302_/B _10302_/Y vdd gnd NAND2X1
XFILL_1__9605_ vdd gnd FILL
X_14070_ _14070_/A _14070_/B _14070_/C _14070_/Y vdd gnd AOI21X1
X_11282_ _11282_/A _11282_/B _11282_/Y vdd gnd NOR2X1
XFILL_1__7797_ vdd gnd FILL
X_13021_ _13021_/A _13021_/B _13021_/C _13021_/Y vdd gnd OAI21X1
X_10233_ _10233_/A _10233_/B _10233_/Y vdd gnd NAND2X1
XFILL_1__9536_ vdd gnd FILL
X_10164_ _10164_/A _10164_/B _10164_/C _10164_/Y vdd gnd OAI21X1
XFILL_1__9467_ vdd gnd FILL
XFILL_2__8260_ vdd gnd FILL
X_10095_ _10095_/A _10095_/B _10095_/Y vdd gnd AND2X2
XFILL_1__8418_ vdd gnd FILL
XFILL_1__9398_ vdd gnd FILL
XFILL_2__8191_ vdd gnd FILL
X_13923_ _13923_/A _13923_/Y vdd gnd INVX1
XFILL_1__8349_ vdd gnd FILL
XFILL_2__10480_ vdd gnd FILL
X_13854_ _13854_/A _13854_/B _13854_/Y vdd gnd NOR2X1
XFILL_0__10610_ vdd gnd FILL
XFILL_1_BUFX2_insert210 vdd gnd FILL
XFILL_0__11590_ vdd gnd FILL
X_12805_ _12805_/A _12805_/B _12805_/Y vdd gnd OR2X2
XFILL_1_BUFX2_insert221 vdd gnd FILL
X_13785_ _13785_/A _13785_/B _13785_/Y vdd gnd NAND2X1
X_10997_ _10997_/A _10997_/B _10997_/C _10997_/Y vdd gnd NAND3X1
XFILL_1__11900_ vdd gnd FILL
XFILL_1_BUFX2_insert232 vdd gnd FILL
XFILL_0__10541_ vdd gnd FILL
XFILL_1_BUFX2_insert243 vdd gnd FILL
XFILL_1_BUFX2_insert254 vdd gnd FILL
XFILL_1__12880_ vdd gnd FILL
XFILL_1_BUFX2_insert265 vdd gnd FILL
X_12736_ _12736_/A _12736_/B _12736_/Y vdd gnd AND2X2
XFILL_1_BUFX2_insert276 vdd gnd FILL
XFILL_2__11101_ vdd gnd FILL
XCLKBUF1_insert36 CLKBUF1_insert36/A CLKBUF1_insert36/Y vdd gnd CLKBUF1
XFILL_2__12081_ vdd gnd FILL
XCLKBUF1_insert47 CLKBUF1_insert47/A CLKBUF1_insert47/Y vdd gnd CLKBUF1
XFILL_1_BUFX2_insert287 vdd gnd FILL
XFILL_1__11831_ vdd gnd FILL
XFILL_0__13260_ vdd gnd FILL
XFILL_0__10472_ vdd gnd FILL
XFILL_1_BUFX2_insert298 vdd gnd FILL
XCLKBUF1_insert58 CLKBUF1_insert58/A CLKBUF1_insert58/Y vdd gnd CLKBUF1
XFILL_2__11032_ vdd gnd FILL
XCLKBUF1_insert69 CLKBUF1_insert69/A CLKBUF1_insert69/Y vdd gnd CLKBUF1
X_12667_ _12667_/A _12667_/Y vdd gnd INVX1
XFILL_0__12211_ vdd gnd FILL
XFILL_0__13191_ vdd gnd FILL
X_14406_ _14406_/A _14406_/Y vdd gnd INVX1
XFILL_1__11762_ vdd gnd FILL
X_11618_ _11618_/D _11618_/CLK _11618_/Q vdd gnd DFFPOSX1
XFILL_0_CLKBUF1_insert391 vdd gnd FILL
X_12598_ _12598_/D _12598_/CLK _12598_/Q vdd gnd DFFPOSX1
XFILL_0__12142_ vdd gnd FILL
XFILL_1__11693_ vdd gnd FILL
XFILL_1__14481_ vdd gnd FILL
X_14337_ _14337_/A _14337_/Y vdd gnd INVX1
X_11549_ _11549_/A _11549_/B _11549_/C _11549_/Y vdd gnd OAI21X1
XFILL_1__10644_ vdd gnd FILL
XFILL_0__12073_ vdd gnd FILL
XFILL_0__8660_ vdd gnd FILL
X_14268_ _14268_/A _14268_/B _14268_/Y vdd gnd NAND2X1
XFILL_2__14722_ vdd gnd FILL
XFILL_0__11024_ vdd gnd FILL
XFILL_2__11934_ vdd gnd FILL
XFILL_1__10575_ vdd gnd FILL
XFILL_1__13363_ vdd gnd FILL
X_13219_ _13219_/A _13219_/B _13219_/Y vdd gnd AND2X2
XFILL_0__7611_ vdd gnd FILL
XFILL_0__8591_ vdd gnd FILL
XFILL_2__8527_ vdd gnd FILL
X_14199_ _14199_/D _14199_/CLK _14199_/Q vdd gnd DFFPOSX1
XFILL_2__14653_ vdd gnd FILL
XFILL_1__12314_ vdd gnd FILL
XFILL_2__11865_ vdd gnd FILL
XFILL_1__13294_ vdd gnd FILL
XFILL_0__7542_ vdd gnd FILL
XFILL_2__8458_ vdd gnd FILL
XFILL_1__12245_ vdd gnd FILL
XFILL_2__14584_ vdd gnd FILL
XFILL_2__11796_ vdd gnd FILL
XFILL_0__12975_ vdd gnd FILL
XFILL_0__7473_ vdd gnd FILL
XFILL_0__14714_ vdd gnd FILL
XFILL_2__8389_ vdd gnd FILL
XFILL_1__12176_ vdd gnd FILL
XFILL_0__9212_ vdd gnd FILL
XFILL_0__11926_ vdd gnd FILL
X_9840_ _9840_/D _9840_/CLK _9840_/Q vdd gnd DFFPOSX1
XFILL_1__11127_ vdd gnd FILL
XFILL_0__14645_ vdd gnd FILL
XFILL_2__10678_ vdd gnd FILL
XFILL_0__11857_ vdd gnd FILL
XFILL_0__9143_ vdd gnd FILL
X_9771_ _9771_/D _9771_/CLK _9771_/Q vdd gnd DFFPOSX1
XFILL_2__12417_ vdd gnd FILL
XFILL_1__11058_ vdd gnd FILL
XFILL_0__10808_ vdd gnd FILL
XFILL_0__14576_ vdd gnd FILL
XFILL_0__11788_ vdd gnd FILL
XFILL_0__9074_ vdd gnd FILL
X_8722_ _8722_/A _8722_/Y vdd gnd INVX1
XFILL_1__10009_ vdd gnd FILL
XFILL_2__12348_ vdd gnd FILL
XFILL_0__13527_ vdd gnd FILL
XFILL_0__8025_ vdd gnd FILL
X_8653_ _8653_/A _8653_/B _8653_/Y vdd gnd NOR2X1
XFILL_1__14817_ vdd gnd FILL
XFILL_2__12279_ vdd gnd FILL
X_7604_ _7604_/A _7604_/B _7604_/C _7604_/Y vdd gnd OAI21X1
XFILL_2__14018_ vdd gnd FILL
X_8584_ _8584_/A _8584_/B _8584_/C _8584_/Y vdd gnd OAI21X1
XFILL_1__14748_ vdd gnd FILL
XFILL_0__12409_ vdd gnd FILL
XFILL_0__13389_ vdd gnd FILL
X_7535_ _7535_/A _7535_/B _7535_/C _7535_/Y vdd gnd OAI21X1
XFILL_0__9976_ vdd gnd FILL
XFILL_1__14679_ vdd gnd FILL
XFILL_0__8927_ vdd gnd FILL
XFILL_1__7720_ vdd gnd FILL
X_7466_ _7466_/A _7466_/B _7466_/C _7466_/Y vdd gnd OAI21X1
X_9205_ _9205_/A _9205_/B _9205_/C _9205_/Y vdd gnd OAI21X1
XFILL_1__7651_ vdd gnd FILL
X_7397_ _7397_/A _7397_/B _7397_/C _7397_/Y vdd gnd AOI21X1
XFILL_0__7809_ vdd gnd FILL
X_9136_ _9136_/A _9136_/B _9136_/C _9136_/Y vdd gnd NOR3X1
XFILL_1__7582_ vdd gnd FILL
XFILL_0__8789_ vdd gnd FILL
XFILL_1__9321_ vdd gnd FILL
X_9067_ _9067_/A _9067_/B _9067_/Y vdd gnd NAND2X1
XFILL_1__9252_ vdd gnd FILL
X_8018_ _8018_/A _8018_/B _8018_/C _8018_/D _8018_/Y vdd gnd AOI22X1
XFILL_1__8203_ vdd gnd FILL
XFILL_1__9183_ vdd gnd FILL
X_10920_ _10920_/A _10920_/B _10920_/Y vdd gnd NOR2X1
XFILL_1__8134_ vdd gnd FILL
X_9969_ _9969_/A _9969_/Y vdd gnd INVX1
X_10851_ _10851_/A _10851_/B _10851_/C _10851_/Y vdd gnd OAI21X1
XFILL_1__8065_ vdd gnd FILL
X_13570_ _13570_/A _13570_/B _13570_/C _13570_/Y vdd gnd OAI21X1
X_10782_ _10782_/A _10782_/B _10782_/C _10782_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert206 vdd gnd FILL
X_12521_ _12521_/A _12521_/B _12521_/C _12521_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert217 vdd gnd FILL
XFILL_0_BUFX2_insert228 vdd gnd FILL
XFILL_0_BUFX2_insert239 vdd gnd FILL
X_12452_ _12452_/A _12452_/B _12452_/Y vdd gnd NAND2X1
XFILL_1__8967_ vdd gnd FILL
XFILL_2__7760_ vdd gnd FILL
X_11403_ _11403_/A _11403_/B _11403_/C _11403_/Y vdd gnd OAI21X1
X_12383_ _12383_/A _12383_/Y vdd gnd INVX1
XFILL_2__7691_ vdd gnd FILL
X_14122_ _14122_/A _14122_/B _14122_/C _14122_/Y vdd gnd OAI21X1
X_11334_ _11334_/A _11334_/B _11334_/C _11334_/D _11334_/Y vdd gnd OAI22X1
XFILL_1__7849_ vdd gnd FILL
X_14053_ _14053_/A _14053_/B _14053_/Y vdd gnd NAND2X1
X_11265_ _11265_/A _11265_/B _11265_/Y vdd gnd AND2X2
XFILL_1__10360_ vdd gnd FILL
X_13004_ _13004_/A _13004_/Y vdd gnd INVX1
X_10216_ _10216_/A _10216_/B _10216_/C _10216_/Y vdd gnd OAI21X1
XFILL_1__9519_ vdd gnd FILL
XFILL_2__8312_ vdd gnd FILL
X_11196_ _11196_/A _11196_/B _11196_/C _11196_/Y vdd gnd NAND3X1
XFILL_1__10291_ vdd gnd FILL
X_10147_ _10147_/A _10147_/B _10147_/C _10147_/Y vdd gnd OAI21X1
XFILL_2__10601_ vdd gnd FILL
XFILL_1__12030_ vdd gnd FILL
XFILL_2__8243_ vdd gnd FILL
XFILL_0__12760_ vdd gnd FILL
X_10078_ _10078_/A _10078_/Y vdd gnd INVX1
XFILL_2__13320_ vdd gnd FILL
XFILL_2__10532_ vdd gnd FILL
XFILL_0__11711_ vdd gnd FILL
XFILL_2__8174_ vdd gnd FILL
XFILL_0__12691_ vdd gnd FILL
X_13906_ _13906_/A _13906_/B _13906_/Y vdd gnd NAND2X1
X_14886_ _14886_/D _14886_/CLK _14886_/Q vdd gnd DFFPOSX1
XFILL_2__13251_ vdd gnd FILL
XFILL_2__10463_ vdd gnd FILL
XFILL_0__14430_ vdd gnd FILL
XFILL_1__13981_ vdd gnd FILL
X_13837_ _13837_/A _13837_/B _13837_/Y vdd gnd NAND2X1
XFILL_2__10394_ vdd gnd FILL
XFILL_0__14361_ vdd gnd FILL
XFILL_1__12932_ vdd gnd FILL
XFILL_0__11573_ vdd gnd FILL
X_13768_ _13768_/A _13768_/B _13768_/C _13768_/Y vdd gnd AOI21X1
XFILL_0__13312_ vdd gnd FILL
XFILL_0__10524_ vdd gnd FILL
XFILL_0__14292_ vdd gnd FILL
XFILL_1__12863_ vdd gnd FILL
X_12719_ _12719_/A _12719_/Y vdd gnd INVX1
XFILL_1__14602_ vdd gnd FILL
X_13699_ _13699_/A _13699_/B _13699_/Y vdd gnd NAND2X1
XFILL_1__11814_ vdd gnd FILL
XFILL_0__13243_ vdd gnd FILL
XFILL_0__10455_ vdd gnd FILL
XFILL_1__12794_ vdd gnd FILL
XFILL_2__11015_ vdd gnd FILL
XFILL_0__13174_ vdd gnd FILL
XFILL_1__11745_ vdd gnd FILL
X_7320_ _7320_/A _7320_/B _7320_/C _7320_/D _7320_/Y vdd gnd AOI22X1
XFILL_0__10386_ vdd gnd FILL
XFILL_0__9761_ vdd gnd FILL
XFILL_0__12125_ vdd gnd FILL
XFILL_2__7889_ vdd gnd FILL
XFILL_1__14464_ vdd gnd FILL
XFILL_0__8712_ vdd gnd FILL
X_7251_ _7251_/A _7251_/B _7251_/C _7251_/Y vdd gnd AOI21X1
XFILL_0__9692_ vdd gnd FILL
XFILL_1__13415_ vdd gnd FILL
XFILL_1__10627_ vdd gnd FILL
XFILL_0__12056_ vdd gnd FILL
XFILL_1__14395_ vdd gnd FILL
XFILL_0__8643_ vdd gnd FILL
X_7182_ _7182_/A _7182_/Y vdd gnd INVX1
XFILL_2__14705_ vdd gnd FILL
XFILL_0__11007_ vdd gnd FILL
XFILL_2__11917_ vdd gnd FILL
XFILL256350x252150 vdd gnd FILL
XFILL_1__13346_ vdd gnd FILL
XFILL_1__10558_ vdd gnd FILL
XFILL_0__8574_ vdd gnd FILL
XFILL_2__14636_ vdd gnd FILL
XFILL_2__11848_ vdd gnd FILL
XFILL_1__10489_ vdd gnd FILL
XFILL_1__13277_ vdd gnd FILL
XFILL_0__7525_ vdd gnd FILL
XFILL_2__14567_ vdd gnd FILL
XFILL_1__12228_ vdd gnd FILL
XFILL_2__11779_ vdd gnd FILL
XFILL_1_BUFX2_insert7 vdd gnd FILL
XFILL_0__12958_ vdd gnd FILL
XFILL_0__7456_ vdd gnd FILL
XFILL_2__13518_ vdd gnd FILL
XFILL_0__11909_ vdd gnd FILL
XFILL_1__12159_ vdd gnd FILL
X_9823_ _9823_/D _9823_/CLK _9823_/Q vdd gnd DFFPOSX1
XFILL_0__12889_ vdd gnd FILL
XFILL_0__7387_ vdd gnd FILL
XFILL_0__14628_ vdd gnd FILL
XFILL_0__9126_ vdd gnd FILL
X_9754_ _9754_/A _9754_/B _9754_/Y vdd gnd NAND2X1
XFILL_0__14559_ vdd gnd FILL
XFILL_0__9057_ vdd gnd FILL
X_8705_ _8705_/A _8705_/Y vdd gnd INVX1
X_9685_ _9685_/A _9685_/B _9685_/Y vdd gnd NAND2X1
XFILL_0__8008_ vdd gnd FILL
XFILL_1__9870_ vdd gnd FILL
X_8636_ _8636_/A _8636_/B _8636_/S _8636_/Y vdd gnd MUX2X1
XFILL_1__8821_ vdd gnd FILL
X_8567_ _8567_/A _8567_/Y vdd gnd INVX1
X_7518_ _7518_/A _7518_/B _7518_/C _7518_/Y vdd gnd OAI21X1
XFILL_0__9959_ vdd gnd FILL
XFILL_1__8752_ vdd gnd FILL
X_8498_ _8498_/A _8498_/B _8498_/C _8498_/Y vdd gnd AOI21X1
XFILL_1__7703_ vdd gnd FILL
X_7449_ _7449_/A _7449_/B _7449_/Y vdd gnd AND2X2
XFILL_1__8683_ vdd gnd FILL
XFILL_1__7634_ vdd gnd FILL
X_11050_ _11050_/A _11050_/B _11050_/C _11050_/Y vdd gnd AOI21X1
X_9119_ _9119_/A _9119_/B _9119_/C _9119_/Y vdd gnd NAND3X1
XFILL_1__7565_ vdd gnd FILL
X_10001_ _10001_/A _10001_/B _10001_/C _10001_/Y vdd gnd OAI21X1
XFILL_1__9304_ vdd gnd FILL
XFILL_1__7496_ vdd gnd FILL
XFILL_1__9235_ vdd gnd FILL
X_14740_ _14740_/A _14740_/B _14740_/Y vdd gnd AND2X2
X_11952_ _11952_/A _11952_/Y vdd gnd INVX1
XFILL_1__9166_ vdd gnd FILL
X_10903_ _10903_/A _10903_/B _10903_/Y vdd gnd NAND2X1
X_14671_ _14671_/A _14671_/B _14671_/C _14671_/Y vdd gnd AOI21X1
XFILL_1__8117_ vdd gnd FILL
X_11883_ _11883_/A _11883_/B _11883_/C _11883_/Y vdd gnd OAI21X1
XFILL_1__9097_ vdd gnd FILL
X_13622_ _13622_/A _13622_/B _13622_/C _13622_/Y vdd gnd AOI21X1
X_10834_ _10834_/A _10834_/B _10834_/Y vdd gnd NAND2X1
XFILL_1__8048_ vdd gnd FILL
X_13553_ _13553_/A _13553_/B _13553_/C _13553_/Y vdd gnd OAI21X1
X_10765_ _10765_/D _10765_/CLK _10765_/Q vdd gnd DFFPOSX1
X_12504_ _12504_/A _12504_/B _12504_/C _12504_/Y vdd gnd OAI21X1
X_13484_ _13484_/D _13484_/CLK _13484_/Q vdd gnd DFFPOSX1
X_10696_ _10696_/D _10696_/CLK _10696_/Q vdd gnd DFFPOSX1
XFILL_0__10240_ vdd gnd FILL
XFILL_1__9999_ vdd gnd FILL
X_12435_ _12435_/A _12435_/B _12435_/C _12435_/Y vdd gnd OAI21X1
XFILL_1__11530_ vdd gnd FILL
XFILL_0__10171_ vdd gnd FILL
X_12366_ _12366_/A _12366_/B _12366_/C _12366_/Y vdd gnd OAI21X1
XFILL_1__11461_ vdd gnd FILL
X_14105_ _14105_/A _14105_/B _14105_/C _14105_/Y vdd gnd OAI21X1
X_11317_ _11317_/A _11317_/B _11317_/C _11317_/Y vdd gnd AOI21X1
XFILL_1__13200_ vdd gnd FILL
X_12297_ _12297_/A _12297_/B _12297_/C _12297_/Y vdd gnd AOI21X1
XFILL_1__10412_ vdd gnd FILL
XFILL_0__13930_ vdd gnd FILL
XFILL_1__11392_ vdd gnd FILL
X_14036_ _14036_/A _14036_/Y vdd gnd INVX1
X_11248_ _11248_/A _11248_/B _11248_/C _11248_/Y vdd gnd OAI21X1
XFILL_1__13131_ vdd gnd FILL
XFILL_1__10343_ vdd gnd FILL
XFILL_0__13861_ vdd gnd FILL
XFILL_2__14421_ vdd gnd FILL
X_11179_ _11179_/A _11179_/B _11179_/C _11179_/Y vdd gnd AOI21X1
XFILL_1__10274_ vdd gnd FILL
XFILL_0__12812_ vdd gnd FILL
XFILL_1__13062_ vdd gnd FILL
XFILL_0__7310_ vdd gnd FILL
XFILL_0__13792_ vdd gnd FILL
XFILL_0__8290_ vdd gnd FILL
XFILL_2__8226_ vdd gnd FILL
XFILL_1__12013_ vdd gnd FILL
XFILL_0__12743_ vdd gnd FILL
XFILL_0__7241_ vdd gnd FILL
XFILL_2__13303_ vdd gnd FILL
XFILL_2__10515_ vdd gnd FILL
XFILL_2__8157_ vdd gnd FILL
XFILL256950x68550 vdd gnd FILL
XFILL_0__12674_ vdd gnd FILL
XFILL_0__7172_ vdd gnd FILL
X_14869_ _14869_/D _14869_/CLK _14869_/Q vdd gnd DFFPOSX1
XFILL256350x64950 vdd gnd FILL
XFILL_2__13234_ vdd gnd FILL
XFILL_2__10446_ vdd gnd FILL
XFILL_0__14413_ vdd gnd FILL
XFILL_2__8088_ vdd gnd FILL
XFILL_1__13964_ vdd gnd FILL
XFILL_2__13165_ vdd gnd FILL
XFILL_1__12915_ vdd gnd FILL
XFILL_2__10377_ vdd gnd FILL
XFILL_0__14344_ vdd gnd FILL
XFILL_0__11556_ vdd gnd FILL
XFILL_1__13895_ vdd gnd FILL
X_9470_ _9470_/A _9470_/Y vdd gnd INVX1
XFILL_0__10507_ vdd gnd FILL
XFILL_2__13096_ vdd gnd FILL
XFILL_1__12846_ vdd gnd FILL
XFILL_0__14275_ vdd gnd FILL
XFILL_0__11487_ vdd gnd FILL
X_8421_ _8421_/A _8421_/B _8421_/C _8421_/Y vdd gnd NAND3X1
XFILL_0__10438_ vdd gnd FILL
XFILL_0__13226_ vdd gnd FILL
XFILL_1__12777_ vdd gnd FILL
X_8352_ _8352_/A _8352_/Y vdd gnd INVX1
XFILL_0__13157_ vdd gnd FILL
XFILL_1__11728_ vdd gnd FILL
XFILL_0__10369_ vdd gnd FILL
X_7303_ _7303_/A _7303_/B _7303_/Y vdd gnd NAND2X1
XFILL_0__9744_ vdd gnd FILL
X_8283_ _8283_/A _8283_/B _8283_/Y vdd gnd NOR2X1
XFILL_0__12108_ vdd gnd FILL
XFILL_1__14447_ vdd gnd FILL
XFILL_0__13088_ vdd gnd FILL
X_7234_ _7234_/A _7234_/Y vdd gnd INVX1
XFILL_0__9675_ vdd gnd FILL
XFILL_0__12039_ vdd gnd FILL
XFILL_1__14378_ vdd gnd FILL
XFILL_0__8626_ vdd gnd FILL
X_7165_ _7165_/A _7165_/B _7165_/C _7165_/Y vdd gnd AOI21X1
XFILL_1__13329_ vdd gnd FILL
XFILL_1__7350_ vdd gnd FILL
XFILL_0__8557_ vdd gnd FILL
X_7096_ _7096_/A _7096_/Y vdd gnd INVX1
XFILL_0__7508_ vdd gnd FILL
XFILL_1__7281_ vdd gnd FILL
XFILL_0__8488_ vdd gnd FILL
XFILL_1__9020_ vdd gnd FILL
XFILL_0__7439_ vdd gnd FILL
X_9806_ _9806_/D _9806_/CLK _9806_/Q vdd gnd DFFPOSX1
X_7998_ _7998_/A _7998_/B _7998_/Y vdd gnd NOR2X1
XFILL_0__9109_ vdd gnd FILL
X_9737_ _9737_/A _9737_/B _9737_/C _9737_/Y vdd gnd OAI21X1
XBUFX2_insert108 BUFX2_insert108/A BUFX2_insert108/Y vdd gnd BUFX2
XFILL_1__9922_ vdd gnd FILL
XBUFX2_insert119 BUFX2_insert119/A BUFX2_insert119/Y vdd gnd BUFX2
X_9668_ _9668_/A _9668_/Y vdd gnd INVX1
X_10550_ _10550_/A _10550_/B _10550_/Y vdd gnd NAND2X1
XFILL_1__9853_ vdd gnd FILL
X_8619_ _8619_/A _8619_/B _8619_/Y vdd gnd NOR2X1
X_9599_ _9599_/A _9599_/B _9599_/C _9599_/Y vdd gnd OAI21X1
X_10481_ _10481_/A _10481_/B _10481_/C _10481_/Y vdd gnd OAI21X1
XFILL_1__8804_ vdd gnd FILL
X_12220_ _12220_/A _12220_/Y vdd gnd INVX1
XFILL_1__8735_ vdd gnd FILL
X_12151_ _12151_/A _12151_/B _12151_/C _12151_/Y vdd gnd OAI21X1
XFILL_1__8666_ vdd gnd FILL
X_11102_ _11102_/A _11102_/B _11102_/C _11102_/Y vdd gnd NAND3X1
XFILL_1__7617_ vdd gnd FILL
X_12082_ _12082_/A _12082_/B _12082_/C _12082_/Y vdd gnd OAI21X1
XFILL_1__8597_ vdd gnd FILL
X_11033_ _11033_/A _11033_/B _11033_/Y vdd gnd NAND2X1
XFILL_1__7548_ vdd gnd FILL
XFILL_2_CLKBUF1_insert389 vdd gnd FILL
XFILL_2__9060_ vdd gnd FILL
XFILL_1__7479_ vdd gnd FILL
XFILL_1__9218_ vdd gnd FILL
X_12984_ _12984_/A _12984_/B _12984_/S _12984_/Y vdd gnd MUX2X1
X_14723_ _14723_/A _14723_/B _14723_/C _14723_/Y vdd gnd AOI21X1
X_11935_ _11935_/A _11935_/B _11935_/Y vdd gnd NOR2X1
XFILL_1__9149_ vdd gnd FILL
X_14654_ _14654_/A _14654_/B _14654_/Y vdd gnd NOR2X1
X_11866_ _11866_/A _11866_/B _11866_/C _11866_/Y vdd gnd NAND3X1
XFILL_0__11410_ vdd gnd FILL
XFILL_2__9962_ vdd gnd FILL
XFILL_1__10961_ vdd gnd FILL
XFILL_0__12390_ vdd gnd FILL
X_13605_ _13605_/A _13605_/B _13605_/S _13605_/Y vdd gnd MUX2X1
X_10817_ _10817_/A _10817_/B _10817_/C _10817_/D _10817_/Y vdd gnd AOI22X1
X_14585_ _14585_/A _14585_/Y vdd gnd INVX1
X_11797_ _11797_/A _11797_/B _11797_/C _11797_/Y vdd gnd OAI21X1
XFILL_1__12700_ vdd gnd FILL
XFILL_2__9893_ vdd gnd FILL
XFILL_0__11341_ vdd gnd FILL
XFILL_1__13680_ vdd gnd FILL
X_13536_ _13536_/A _13536_/B _13536_/Y vdd gnd NAND2X1
XFILL_1__10892_ vdd gnd FILL
X_10748_ _10748_/D _10748_/CLK _10748_/Q vdd gnd DFFPOSX1
XFILL_0__14060_ vdd gnd FILL
XFILL_1__12631_ vdd gnd FILL
XFILL_0__11272_ vdd gnd FILL
X_13467_ _13467_/D _13467_/CLK _13467_/Q vdd gnd DFFPOSX1
X_10679_ _10679_/A _10679_/B _10679_/C _10679_/Y vdd gnd OAI21X1
XFILL_0__13011_ vdd gnd FILL
XFILL_0__10223_ vdd gnd FILL
XFILL_2__8775_ vdd gnd FILL
X_12418_ _12418_/A _12418_/Y vdd gnd INVX1
XFILL_0__7790_ vdd gnd FILL
XFILL_1__14301_ vdd gnd FILL
X_13398_ _13398_/A _13398_/B _13398_/Y vdd gnd NAND2X1
XFILL256950x43350 vdd gnd FILL
XFILL_1__11513_ vdd gnd FILL
XFILL_0__10154_ vdd gnd FILL
XFILL_1__12493_ vdd gnd FILL
X_12349_ _12349_/A _12349_/B _12349_/Y vdd gnd NOR2X1
XFILL_2__12803_ vdd gnd FILL
XFILL_1__14232_ vdd gnd FILL
XFILL_1__11444_ vdd gnd FILL
XFILL_0__10085_ vdd gnd FILL
XFILL_0__9460_ vdd gnd FILL
XFILL_0__13913_ vdd gnd FILL
XFILL_0__8411_ vdd gnd FILL
XFILL_1__11375_ vdd gnd FILL
X_14019_ _14019_/A _14019_/B _14019_/C _14019_/Y vdd gnd NAND3X1
XFILL_0__9391_ vdd gnd FILL
XFILL_1__13114_ vdd gnd FILL
XFILL_1__10326_ vdd gnd FILL
XFILL_0__13844_ vdd gnd FILL
XFILL_1__14094_ vdd gnd FILL
XFILL_0__8342_ vdd gnd FILL
XFILL_2__14404_ vdd gnd FILL
X_8970_ _8970_/A _8970_/B _8970_/Y vdd gnd NAND2X1
XFILL_1__10257_ vdd gnd FILL
XFILL_1__13045_ vdd gnd FILL
XFILL_0__13775_ vdd gnd FILL
XFILL_0__10987_ vdd gnd FILL
X_7921_ _7921_/D _7921_/CLK _7921_/Q vdd gnd DFFPOSX1
XFILL_0__8273_ vdd gnd FILL
XFILL_2__14335_ vdd gnd FILL
XFILL_1__10188_ vdd gnd FILL
XFILL_0__12726_ vdd gnd FILL
XFILL_0__7224_ vdd gnd FILL
X_7852_ _7852_/A _7852_/B _7852_/Y vdd gnd NAND2X1
XFILL_2__14266_ vdd gnd FILL
XFILL_0__12657_ vdd gnd FILL
XFILL_0__7155_ vdd gnd FILL
XFILL_2__13217_ vdd gnd FILL
X_7783_ _7783_/A _7783_/Y vdd gnd INVX1
XFILL_0__11608_ vdd gnd FILL
XFILL_1__13947_ vdd gnd FILL
X_9522_ _9522_/A _9522_/B _9522_/C _9522_/D _9522_/Y vdd gnd AOI22X1
XFILL_0__7086_ vdd gnd FILL
XFILL_2__13148_ vdd gnd FILL
XFILL_0__14327_ vdd gnd FILL
XFILL_1__13878_ vdd gnd FILL
XFILL_0__11539_ vdd gnd FILL
X_9453_ _9453_/A _9453_/B _9453_/C _9453_/Y vdd gnd NAND3X1
XFILL_2__13079_ vdd gnd FILL
XFILL_1__12829_ vdd gnd FILL
XFILL_0__14258_ vdd gnd FILL
X_8404_ _8404_/A _8404_/B _8404_/Y vdd gnd AND2X2
X_9384_ _9384_/A _9384_/Y vdd gnd INVX1
XFILL_0__13209_ vdd gnd FILL
X_8335_ _8335_/A _8335_/B _8335_/C _8335_/Y vdd gnd AOI21X1
XFILL_1__8520_ vdd gnd FILL
XFILL_0__9727_ vdd gnd FILL
X_8266_ _8266_/A _8266_/B _8266_/Y vdd gnd NAND2X1
X_7217_ _7217_/A _7217_/Y vdd gnd INVX1
XFILL_0__9658_ vdd gnd FILL
XFILL_1__8451_ vdd gnd FILL
X_8197_ _8197_/A _8197_/B _8197_/Y vdd gnd AND2X2
XFILL_1__7402_ vdd gnd FILL
XFILL_0__8609_ vdd gnd FILL
X_7148_ _7148_/A _7148_/B _7148_/S _7148_/Y vdd gnd MUX2X1
XFILL_0__9589_ vdd gnd FILL
XFILL_1__8382_ vdd gnd FILL
XFILL_1__7333_ vdd gnd FILL
X_7079_ _7079_/A _7079_/B _7079_/C _7079_/Y vdd gnd OAI21X1
XFILL_1__7264_ vdd gnd FILL
XFILL_1__9003_ vdd gnd FILL
XFILL_1__7195_ vdd gnd FILL
X_11720_ _11720_/A _11720_/B _11720_/Y vdd gnd NAND2X1
X_11651_ _11651_/D _11651_/CLK _11651_/Q vdd gnd DFFPOSX1
X_10602_ _10602_/A _10602_/B _10602_/C _10602_/Y vdd gnd OAI21X1
X_14370_ _14370_/A _14370_/B _14370_/Y vdd gnd NAND2X1
XFILL_1__9905_ vdd gnd FILL
X_11582_ _11582_/A _11582_/B _11582_/Y vdd gnd NAND2X1
X_13321_ _13321_/A _13321_/B _13321_/C _13321_/Y vdd gnd OAI21X1
X_10533_ _10533_/A _10533_/B _10533_/C _10533_/D _10533_/Y vdd gnd OAI22X1
X_13252_ _13252_/A _13252_/Y vdd gnd INVX1
X_10464_ _10464_/A _10464_/B _10464_/C _10464_/Y vdd gnd OAI21X1
XFILL_2__8560_ vdd gnd FILL
X_12203_ _12203_/A _12203_/B _12203_/C _12203_/Y vdd gnd NAND3X1
X_13183_ _13183_/A _13183_/B _13183_/Y vdd gnd OR2X2
X_10395_ _10395_/A _10395_/B _10395_/C _10395_/Y vdd gnd NAND3X1
XFILL_1__8718_ vdd gnd FILL
XFILL_1__9698_ vdd gnd FILL
XFILL_2__8491_ vdd gnd FILL
X_12134_ _12134_/A _12134_/B _12134_/Y vdd gnd NAND2X1
XFILL_1__8649_ vdd gnd FILL
X_12065_ _12065_/A _12065_/B _12065_/Y vdd gnd NAND2X1
XFILL_1__11160_ vdd gnd FILL
XFILL_0__10910_ vdd gnd FILL
X_11016_ _11016_/A _11016_/B _11016_/C _11016_/D _11016_/Y vdd gnd AOI22X1
XFILL_2__9112_ vdd gnd FILL
XFILL_0__11890_ vdd gnd FILL
XFILL_1__10111_ vdd gnd FILL
XFILL_1__11091_ vdd gnd FILL
XFILL_0__10841_ vdd gnd FILL
XFILL_2__9043_ vdd gnd FILL
XFILL_2__11401_ vdd gnd FILL
XFILL_1__10042_ vdd gnd FILL
XFILL_0__10772_ vdd gnd FILL
XFILL_0__13560_ vdd gnd FILL
XBUFX2_insert8 BUFX2_insert8/A BUFX2_insert8/Y vdd gnd BUFX2
X_12967_ _12967_/A _12967_/B _12967_/C _12967_/Y vdd gnd AOI21X1
XFILL_2__11332_ vdd gnd FILL
XFILL_1__14850_ vdd gnd FILL
XFILL_0__12511_ vdd gnd FILL
X_14706_ _14706_/A _14706_/B _14706_/Y vdd gnd NAND2X1
X_11918_ _11918_/A _11918_/B _11918_/C _11918_/Y vdd gnd OAI21X1
X_12898_ _12898_/A _12898_/B _12898_/C _12898_/Y vdd gnd OAI21X1
XFILL_2__14051_ vdd gnd FILL
XFILL_1__13801_ vdd gnd FILL
XFILL_2__11263_ vdd gnd FILL
XFILL_1__14781_ vdd gnd FILL
XFILL_0__12442_ vdd gnd FILL
XFILL_1__11993_ vdd gnd FILL
X_14637_ _14637_/A _14637_/B _14637_/C _14637_/Y vdd gnd AOI21X1
X_11849_ _11849_/A _11849_/B _11849_/C _11849_/Y vdd gnd OAI21X1
XFILL_2__9945_ vdd gnd FILL
XFILL_1__13732_ vdd gnd FILL
XFILL_1__10944_ vdd gnd FILL
XFILL_0__12373_ vdd gnd FILL
XFILL_2__11194_ vdd gnd FILL
XFILL_0__8960_ vdd gnd FILL
X_14568_ _14568_/A _14568_/Y vdd gnd INVX1
XFILL_0__14112_ vdd gnd FILL
XFILL_0__11324_ vdd gnd FILL
XFILL_1__13663_ vdd gnd FILL
XFILL_2__9876_ vdd gnd FILL
XFILL_0__7911_ vdd gnd FILL
XFILL_1__10875_ vdd gnd FILL
X_13519_ _13519_/A _13519_/Y vdd gnd INVX1
X_14499_ _14499_/A _14499_/B _14499_/C _14499_/Y vdd gnd OAI21X1
XFILL_2__8827_ vdd gnd FILL
XFILL_0__14043_ vdd gnd FILL
XFILL_0__11255_ vdd gnd FILL
XFILL_1__13594_ vdd gnd FILL
XFILL_0__7842_ vdd gnd FILL
XFILL_0__10206_ vdd gnd FILL
XFILL_2__13904_ vdd gnd FILL
XFILL_2__8758_ vdd gnd FILL
XFILL_0__11186_ vdd gnd FILL
X_8120_ _8120_/A _8120_/B _8120_/C _8120_/Y vdd gnd AOI21X1
XFILL_0__7773_ vdd gnd FILL
XFILL_2__13835_ vdd gnd FILL
XFILL_0__10137_ vdd gnd FILL
XFILL_2__8689_ vdd gnd FILL
XFILL_0__9512_ vdd gnd FILL
XFILL_1__12476_ vdd gnd FILL
X_8051_ _8051_/A _8051_/B _8051_/C _8051_/Y vdd gnd OAI21X1
XFILL_1__11427_ vdd gnd FILL
XFILL_0__10068_ vdd gnd FILL
XFILL_0__9443_ vdd gnd FILL
XFILL_1_BUFX2_insert12 vdd gnd FILL
XFILL_1_BUFX2_insert23 vdd gnd FILL
XFILL_2__12717_ vdd gnd FILL
XFILL_1__14146_ vdd gnd FILL
XFILL_1__11358_ vdd gnd FILL
XFILL_0__9374_ vdd gnd FILL
XFILL_1__10309_ vdd gnd FILL
XFILL_2__12648_ vdd gnd FILL
XFILL_1__14077_ vdd gnd FILL
XFILL_0__13827_ vdd gnd FILL
XFILL_0__8325_ vdd gnd FILL
XFILL_1__11289_ vdd gnd FILL
X_8953_ _8953_/A _8953_/Y vdd gnd INVX1
XFILL_1__13028_ vdd gnd FILL
XFILL_0__13758_ vdd gnd FILL
X_7904_ _7904_/A _7904_/B _7904_/Y vdd gnd NAND2X1
XFILL_0__8256_ vdd gnd FILL
XFILL_2__14318_ vdd gnd FILL
X_8884_ _8884_/D _8884_/CLK _8884_/Q vdd gnd DFFPOSX1
XFILL_0__12709_ vdd gnd FILL
XFILL_0__7207_ vdd gnd FILL
XFILL_0__13689_ vdd gnd FILL
X_7835_ _7835_/A _7835_/B _7835_/Y vdd gnd NAND2X1
XFILL_0__8187_ vdd gnd FILL
XFILL_2__14249_ vdd gnd FILL
XFILL_1_CLKBUF1_insert35 vdd gnd FILL
XFILL_0__7138_ vdd gnd FILL
XFILL_1_CLKBUF1_insert46 vdd gnd FILL
XFILL_1_CLKBUF1_insert57 vdd gnd FILL
X_7766_ _7766_/A _7766_/Y vdd gnd INVX1
XFILL_1_CLKBUF1_insert68 vdd gnd FILL
XFILL_1_CLKBUF1_insert79 vdd gnd FILL
X_9505_ _9505_/A _9505_/B _9505_/Y vdd gnd NOR2X1
X_7697_ _7697_/A _7697_/B _7697_/Y vdd gnd NOR2X1
X_9436_ _9436_/A _9436_/B _9436_/Y vdd gnd NAND2X1
XFILL_1__7882_ vdd gnd FILL
XFILL_1__9621_ vdd gnd FILL
X_9367_ _9367_/A _9367_/B _9367_/Y vdd gnd OR2X2
XFILL_1__9552_ vdd gnd FILL
X_8318_ _8318_/A _8318_/Y vdd gnd INVX1
X_9298_ _9298_/A _9298_/B _9298_/Y vdd gnd NOR2X1
XFILL_1__8503_ vdd gnd FILL
X_10180_ _10180_/A _10180_/B _10180_/C _10180_/Y vdd gnd AOI21X1
XFILL_1__9483_ vdd gnd FILL
X_8249_ _8249_/A _8249_/B _8249_/C _8249_/Y vdd gnd AOI21X1
XFILL_1__8434_ vdd gnd FILL
XFILL_1__8365_ vdd gnd FILL
XFILL_1__7316_ vdd gnd FILL
X_13870_ _13870_/A _13870_/B _13870_/C _13870_/Y vdd gnd OAI21X1
XFILL_1__8296_ vdd gnd FILL
X_12821_ _12821_/A _12821_/B _12821_/C _12821_/Y vdd gnd AOI21X1
XFILL_1__7247_ vdd gnd FILL
X_12752_ _12752_/A _12752_/B _12752_/C _12752_/Y vdd gnd AOI21X1
XFILL_1__7178_ vdd gnd FILL
X_11703_ _11703_/A _11703_/B _11703_/C _11703_/Y vdd gnd OAI21X1
X_12683_ _12683_/A _12683_/B _12683_/C _12683_/Y vdd gnd OAI21X1
X_14422_ _14422_/A _14422_/B _14422_/Y vdd gnd NAND2X1
X_11634_ _11634_/D _11634_/CLK _11634_/Q vdd gnd DFFPOSX1
X_14353_ _14353_/A _14353_/B _14353_/C _14353_/Y vdd gnd OAI21X1
X_11565_ _11565_/A _11565_/B _11565_/C _11565_/Y vdd gnd OAI21X1
XFILL_1__10660_ vdd gnd FILL
X_13304_ _13304_/A _13304_/Y vdd gnd INVX1
X_10516_ _10516_/A _10516_/B _10516_/C _10516_/Y vdd gnd AOI21X1
X_14284_ _14284_/A _14284_/B _14284_/Y vdd gnd NAND2X1
X_11496_ _11496_/A _11496_/B _11496_/Y vdd gnd NOR2X1
XFILL_0__11040_ vdd gnd FILL
XFILL_2__11950_ vdd gnd FILL
XFILL_1__10591_ vdd gnd FILL
X_13235_ _13235_/A _13235_/B _13235_/Y vdd gnd NAND2X1
X_10447_ _10447_/A _10447_/B _10447_/Y vdd gnd NAND2X1
XFILL_2__8543_ vdd gnd FILL
XFILL_1__12330_ vdd gnd FILL
XFILL_2__11881_ vdd gnd FILL
X_13166_ _13166_/A _13166_/B _13166_/Y vdd gnd NAND2X1
X_10378_ _10378_/A _10378_/Y vdd gnd INVX1
XFILL_2__13620_ vdd gnd FILL
XFILL_2__8474_ vdd gnd FILL
XFILL_1__12261_ vdd gnd FILL
X_12117_ _12117_/A _12117_/B _12117_/C _12117_/Y vdd gnd NAND3X1
XFILL_0__12991_ vdd gnd FILL
XFILL_1__14000_ vdd gnd FILL
X_13097_ _13097_/A _13097_/B _13097_/Y vdd gnd NOR2X1
XFILL_2__13551_ vdd gnd FILL
XFILL_1__11212_ vdd gnd FILL
XFILL_0__14730_ vdd gnd FILL
XFILL_0__11942_ vdd gnd FILL
XFILL_1__12192_ vdd gnd FILL
X_12048_ _12048_/A _12048_/Y vdd gnd INVX1
XFILL_1__11143_ vdd gnd FILL
XFILL_0__14661_ vdd gnd FILL
XFILL_0__11873_ vdd gnd FILL
XFILL_0__13612_ vdd gnd FILL
XFILL_1__11074_ vdd gnd FILL
XFILL_0__8110_ vdd gnd FILL
XFILL_0__10824_ vdd gnd FILL
XFILL_0__14592_ vdd gnd FILL
XFILL_2__9026_ vdd gnd FILL
XFILL_0__9090_ vdd gnd FILL
XFILL_2_BUFX2_insert270 vdd gnd FILL
X_13999_ _13999_/A _13999_/B _13999_/C _13999_/Y vdd gnd AOI21X1
XFILL_1__10025_ vdd gnd FILL
XFILL_0__13543_ vdd gnd FILL
XFILL_0__8041_ vdd gnd FILL
XFILL_2__11315_ vdd gnd FILL
XFILL_1__14833_ vdd gnd FILL
XFILL_0__10686_ vdd gnd FILL
X_7620_ _7620_/A _7620_/B _7620_/Y vdd gnd NOR2X1
XFILL_2__11246_ vdd gnd FILL
XFILL_1__14764_ vdd gnd FILL
XFILL_0__12425_ vdd gnd FILL
XFILL_1__11976_ vdd gnd FILL
X_7551_ _7551_/A _7551_/Y vdd gnd INVX1
XFILL_0__9992_ vdd gnd FILL
XFILL_2__9928_ vdd gnd FILL
XFILL_1__13715_ vdd gnd FILL
XFILL_2__11177_ vdd gnd FILL
XFILL_1__10927_ vdd gnd FILL
XFILL_1__14695_ vdd gnd FILL
XFILL_0__12356_ vdd gnd FILL
XFILL_0__8943_ vdd gnd FILL
X_7482_ _7482_/A _7482_/B _7482_/Y vdd gnd OR2X2
XBUFX2_insert280 BUFX2_insert280/A BUFX2_insert280/Y vdd gnd BUFX2
XFILL_2__9859_ vdd gnd FILL
XFILL_1__13646_ vdd gnd FILL
XFILL_0__11307_ vdd gnd FILL
XBUFX2_insert291 BUFX2_insert291/A BUFX2_insert291/Y vdd gnd BUFX2
XFILL_1__10858_ vdd gnd FILL
X_9221_ _9221_/A _9221_/B _9221_/Y vdd gnd AND2X2
XFILL_0__12287_ vdd gnd FILL
XFILL_0__14026_ vdd gnd FILL
XFILL_1__13577_ vdd gnd FILL
XFILL_0__11238_ vdd gnd FILL
XFILL_0__7825_ vdd gnd FILL
XFILL_1__10789_ vdd gnd FILL
X_9152_ _9152_/A _9152_/B _9152_/C _9152_/Y vdd gnd OAI21X1
XFILL_1__12528_ vdd gnd FILL
XFILL_2__14867_ vdd gnd FILL
XFILL_0__11169_ vdd gnd FILL
X_8103_ _8103_/A _8103_/Y vdd gnd INVX1
XFILL_0__7756_ vdd gnd FILL
X_9083_ _9083_/A _9083_/Y vdd gnd INVX1
XFILL_2__13818_ vdd gnd FILL
XFILL_1__12459_ vdd gnd FILL
XFILL_2__14798_ vdd gnd FILL
X_8034_ _8034_/A _8034_/B _8034_/C _8034_/Y vdd gnd OAI21X1
XFILL_0__7687_ vdd gnd FILL
XFILL_2__13749_ vdd gnd FILL
XFILL_0__9426_ vdd gnd FILL
XFILL_1__14129_ vdd gnd FILL
XFILL_0__14859_ vdd gnd FILL
XFILL_0__9357_ vdd gnd FILL
XFILL_1__8150_ vdd gnd FILL
X_9985_ _9985_/A _9985_/B _9985_/C _9985_/D _9985_/Y vdd gnd OAI22X1
XFILL_1__7101_ vdd gnd FILL
XFILL_0__8308_ vdd gnd FILL
XFILL_0__9288_ vdd gnd FILL
X_8936_ _8936_/A _8936_/B _8936_/C _8936_/Y vdd gnd OAI21X1
XFILL_1__8081_ vdd gnd FILL
XFILL_0__8239_ vdd gnd FILL
X_8867_ _8867_/D _8867_/CLK _8867_/Q vdd gnd DFFPOSX1
X_7818_ _7818_/A _7818_/B _7818_/C _7818_/Y vdd gnd OAI21X1
X_8798_ _8798_/A _8798_/B _8798_/Y vdd gnd NAND2X1
X_7749_ _7749_/A _7749_/Y vdd gnd INVX1
XFILL_1__8983_ vdd gnd FILL
X_11350_ _11350_/A _11350_/Y vdd gnd INVX1
X_9419_ _9419_/A _9419_/B _9419_/C _9419_/Y vdd gnd OAI21X1
XFILL_1__7865_ vdd gnd FILL
X_10301_ _10301_/A _10301_/B _10301_/C _10301_/Y vdd gnd AOI21X1
XFILL_1__9604_ vdd gnd FILL
X_11281_ _11281_/A _11281_/B _11281_/C _11281_/Y vdd gnd AOI21X1
XFILL_1__7796_ vdd gnd FILL
X_13020_ _13020_/A _13020_/B _13020_/C _13020_/Y vdd gnd AOI21X1
X_10232_ _10232_/A _10232_/B _10232_/C _10232_/Y vdd gnd OAI21X1
XFILL_1__9535_ vdd gnd FILL
X_10163_ _10163_/A _10163_/B _10163_/C _10163_/Y vdd gnd OAI21X1
XFILL_1__9466_ vdd gnd FILL
XFILL_2__7210_ vdd gnd FILL
X_10094_ _10094_/A _10094_/B _10094_/C _10094_/Y vdd gnd AOI21X1
XFILL_1__8417_ vdd gnd FILL
XFILL_1__9397_ vdd gnd FILL
X_13922_ _13922_/A _13922_/B _13922_/C _13922_/Y vdd gnd OAI21X1
XFILL_2__7141_ vdd gnd FILL
XFILL_1__8348_ vdd gnd FILL
X_13853_ _13853_/A _13853_/B _13853_/Y vdd gnd NOR2X1
XFILL_2__7072_ vdd gnd FILL
XFILL_1__8279_ vdd gnd FILL
XFILL_1_BUFX2_insert200 vdd gnd FILL
X_12804_ _12804_/A _12804_/B _12804_/C _12804_/Y vdd gnd OAI21X1
XFILL_1_BUFX2_insert211 vdd gnd FILL
X_10996_ _10996_/A _10996_/Y vdd gnd INVX1
XFILL_1_BUFX2_insert222 vdd gnd FILL
X_13784_ _13784_/A _13784_/B _13784_/C _13784_/D _13784_/Y vdd gnd AOI22X1
XFILL_1_BUFX2_insert233 vdd gnd FILL
XFILL_0__10540_ vdd gnd FILL
XFILL_1_BUFX2_insert244 vdd gnd FILL
XFILL257550x93750 vdd gnd FILL
XFILL_1_BUFX2_insert255 vdd gnd FILL
X_12735_ _12735_/A _12735_/B _12735_/C _12735_/Y vdd gnd NAND3X1
XFILL_1_BUFX2_insert266 vdd gnd FILL
XFILL_1_BUFX2_insert277 vdd gnd FILL
XFILL_1__11830_ vdd gnd FILL
XFILL_0__10471_ vdd gnd FILL
XFILL_1_BUFX2_insert288 vdd gnd FILL
XCLKBUF1_insert37 CLKBUF1_insert37/A CLKBUF1_insert37/Y vdd gnd CLKBUF1
XCLKBUF1_insert48 CLKBUF1_insert48/A CLKBUF1_insert48/Y vdd gnd CLKBUF1
XFILL_1_BUFX2_insert299 vdd gnd FILL
XCLKBUF1_insert59 CLKBUF1_insert59/A CLKBUF1_insert59/Y vdd gnd CLKBUF1
X_12666_ _12666_/A _12666_/B _12666_/C _12666_/Y vdd gnd OAI21X1
XFILL_0__12210_ vdd gnd FILL
XFILL_0__13190_ vdd gnd FILL
XFILL_1__11761_ vdd gnd FILL
X_14405_ _14405_/A _14405_/B _14405_/C _14405_/Y vdd gnd OAI21X1
X_11617_ _11617_/D _11617_/CLK _11617_/Q vdd gnd DFFPOSX1
XFILL_2__9713_ vdd gnd FILL
X_12597_ _12597_/D _12597_/CLK _12597_/Q vdd gnd DFFPOSX1
XFILL_1__14480_ vdd gnd FILL
XFILL_0__12141_ vdd gnd FILL
XFILL_1__11692_ vdd gnd FILL
X_14336_ _14336_/A _14336_/B _14336_/Y vdd gnd NAND2X1
X_11548_ _11548_/A _11548_/B _11548_/Y vdd gnd NAND2X1
XFILL_1__10643_ vdd gnd FILL
XFILL_0__12072_ vdd gnd FILL
X_14267_ _14267_/A _14267_/B _14267_/C _14267_/Y vdd gnd OAI21X1
X_11479_ _11479_/A _11479_/Y vdd gnd INVX1
XFILL_0__11023_ vdd gnd FILL
XFILL_1__13362_ vdd gnd FILL
X_13218_ _13218_/A _13218_/B _13218_/Y vdd gnd NOR2X1
XFILL_0__7610_ vdd gnd FILL
XFILL_1__10574_ vdd gnd FILL
XFILL_0__8590_ vdd gnd FILL
X_14198_ _14198_/D _14198_/CLK _14198_/Q vdd gnd DFFPOSX1
XFILL_1__12313_ vdd gnd FILL
XFILL_1__13293_ vdd gnd FILL
X_13149_ _13149_/A _13149_/B _13149_/C _13149_/Y vdd gnd NAND3X1
XFILL_0__7541_ vdd gnd FILL
XFILL_2__10815_ vdd gnd FILL
XFILL_2__13603_ vdd gnd FILL
XFILL_1__12244_ vdd gnd FILL
XFILL_0__12974_ vdd gnd FILL
XFILL_0__7472_ vdd gnd FILL
XFILL_2__7408_ vdd gnd FILL
XFILL_2__13534_ vdd gnd FILL
XFILL_0__14713_ vdd gnd FILL
XFILL_0__9211_ vdd gnd FILL
XFILL_0__11925_ vdd gnd FILL
XFILL_1__12175_ vdd gnd FILL
XFILL_2__7339_ vdd gnd FILL
XFILL_1__11126_ vdd gnd FILL
XFILL_0__14644_ vdd gnd FILL
XFILL_0__9142_ vdd gnd FILL
XFILL_0__11856_ vdd gnd FILL
X_9770_ _9770_/D _9770_/CLK _9770_/Q vdd gnd DFFPOSX1
XFILL_1__11057_ vdd gnd FILL
XFILL_2__13396_ vdd gnd FILL
XFILL_0__10807_ vdd gnd FILL
XFILL_0__14575_ vdd gnd FILL
XFILL_0__9073_ vdd gnd FILL
X_8721_ _8721_/A _8721_/B _8721_/C _8721_/Y vdd gnd NAND3X1
XFILL_0__11787_ vdd gnd FILL
XFILL_2__9009_ vdd gnd FILL
XFILL_1__10008_ vdd gnd FILL
XFILL_0__13526_ vdd gnd FILL
XFILL_0__8024_ vdd gnd FILL
X_8652_ _8652_/A _8652_/B _8652_/C _8652_/Y vdd gnd OAI21X1
XFILL_1__14816_ vdd gnd FILL
X_7603_ _7603_/A _7603_/Y vdd gnd INVX1
XFILL_0__10669_ vdd gnd FILL
XFILL_2__11229_ vdd gnd FILL
X_8583_ _8583_/A _8583_/B _8583_/C _8583_/Y vdd gnd OAI21X1
XFILL_1__14747_ vdd gnd FILL
XFILL_0__12408_ vdd gnd FILL
XFILL_1__11959_ vdd gnd FILL
XFILL_0__13388_ vdd gnd FILL
X_7534_ _7534_/A _7534_/B _7534_/Y vdd gnd NAND2X1
XFILL_0__9975_ vdd gnd FILL
XFILL_1__14678_ vdd gnd FILL
XFILL_0__12339_ vdd gnd FILL
XFILL_0__8926_ vdd gnd FILL
X_7465_ _7465_/A _7465_/B _7465_/Y vdd gnd NAND2X1
XFILL_1__13629_ vdd gnd FILL
X_9204_ _9204_/A _9204_/B _9204_/Y vdd gnd OR2X2
XFILL_1__7650_ vdd gnd FILL
X_7396_ _7396_/A _7396_/Y vdd gnd INVX1
XFILL_0__14009_ vdd gnd FILL
X_9135_ _9135_/A _9135_/B _9135_/C _9135_/Y vdd gnd NAND3X1
XFILL_0__7808_ vdd gnd FILL
XFILL_1__7581_ vdd gnd FILL
XFILL_0__8788_ vdd gnd FILL
XFILL_1__9320_ vdd gnd FILL
X_9066_ _9066_/A _9066_/B _9066_/C _9066_/Y vdd gnd OAI21X1
XFILL_0__7739_ vdd gnd FILL
XFILL_1__9251_ vdd gnd FILL
X_8017_ _8017_/A _8017_/B _8017_/C _8017_/Y vdd gnd OAI21X1
XFILL_1__8202_ vdd gnd FILL
XFILL_0__9409_ vdd gnd FILL
XFILL_1__9182_ vdd gnd FILL
XFILL_1__8133_ vdd gnd FILL
X_9968_ _9968_/A _9968_/B _9968_/C _9968_/Y vdd gnd AOI21X1
X_10850_ _10850_/A _10850_/Y vdd gnd INVX2
X_8919_ _8919_/D _8919_/CLK _8919_/Q vdd gnd DFFPOSX1
XFILL_1__8064_ vdd gnd FILL
X_9899_ _9899_/A _9899_/B _9899_/C _9899_/Y vdd gnd OAI21X1
X_10781_ _10781_/A _10781_/B _10781_/C _10781_/D _10781_/Y vdd gnd AOI22X1
X_12520_ _12520_/A _12520_/B _12520_/Y vdd gnd NAND2X1
XFILL_0_BUFX2_insert207 vdd gnd FILL
XFILL_0_BUFX2_insert218 vdd gnd FILL
XFILL_0_BUFX2_insert229 vdd gnd FILL
XFILL257550x25350 vdd gnd FILL
X_12451_ _12451_/A _12451_/B _12451_/C _12451_/Y vdd gnd OAI21X1
XFILL_1__8966_ vdd gnd FILL
X_11402_ _11402_/A _11402_/B _11402_/Y vdd gnd NAND2X1
X_12382_ _12382_/A _12382_/B _12382_/Y vdd gnd NAND2X1
X_14121_ _14121_/A _14121_/B _14121_/Y vdd gnd NAND2X1
X_11333_ _11333_/A _11333_/B _11333_/C _11333_/Y vdd gnd OAI21X1
XFILL_1__7848_ vdd gnd FILL
X_14052_ _14052_/A _14052_/B _14052_/C _14052_/D _14052_/Y vdd gnd OAI22X1
X_11264_ _11264_/A _11264_/B _11264_/Y vdd gnd NOR2X1
XFILL_2__9360_ vdd gnd FILL
XFILL_1__7779_ vdd gnd FILL
X_13003_ _13003_/A _13003_/B _13003_/C _13003_/Y vdd gnd OAI21X1
X_10215_ _10215_/A _10215_/B _10215_/Y vdd gnd NAND2X1
XFILL_1__9518_ vdd gnd FILL
X_11195_ _11195_/A _11195_/B _11195_/C _11195_/Y vdd gnd OAI21X1
XFILL_2__9291_ vdd gnd FILL
XFILL_1__10290_ vdd gnd FILL
X_10146_ _10146_/A _10146_/B _10146_/C _10146_/Y vdd gnd NAND3X1
XFILL_1__9449_ vdd gnd FILL
XFILL_2__11580_ vdd gnd FILL
X_10077_ _10077_/A _10077_/B _10077_/C _10077_/Y vdd gnd NAND3X1
XFILL_0__11710_ vdd gnd FILL
XFILL_0__12690_ vdd gnd FILL
X_13905_ _13905_/A _13905_/B _13905_/C _13905_/Y vdd gnd OAI21X1
XFILL_2__7124_ vdd gnd FILL
X_14885_ _14885_/D _14885_/CLK _14885_/Q vdd gnd DFFPOSX1
XFILL_1__13980_ vdd gnd FILL
XFILL_2__12201_ vdd gnd FILL
X_13836_ _13836_/A _13836_/B _13836_/Y vdd gnd NAND2X1
XFILL_2__13181_ vdd gnd FILL
XFILL_1__12931_ vdd gnd FILL
XFILL_0__14360_ vdd gnd FILL
XFILL_0__11572_ vdd gnd FILL
X_10979_ _10979_/A _10979_/Y vdd gnd INVX1
XFILL_2__12132_ vdd gnd FILL
X_13767_ _13767_/A _13767_/B _13767_/Y vdd gnd NOR2X1
XFILL_0__13311_ vdd gnd FILL
XFILL_0__10523_ vdd gnd FILL
XFILL_1__12862_ vdd gnd FILL
XFILL_0__14291_ vdd gnd FILL
X_12718_ _12718_/A _12718_/B _12718_/C _12718_/Y vdd gnd OAI21X1
XFILL_1__14601_ vdd gnd FILL
XFILL_1__11813_ vdd gnd FILL
X_13698_ _13698_/A _13698_/B _13698_/C _13698_/Y vdd gnd AOI21X1
XFILL_0__13242_ vdd gnd FILL
XFILL_0__10454_ vdd gnd FILL
XFILL_1__12793_ vdd gnd FILL
X_12649_ _12649_/A _12649_/B _12649_/C _12649_/D _12649_/Y vdd gnd AOI22X1
XFILL_1__11744_ vdd gnd FILL
XFILL_0__13173_ vdd gnd FILL
XFILL_0__10385_ vdd gnd FILL
XFILL_0__9760_ vdd gnd FILL
XFILL_1__14463_ vdd gnd FILL
XFILL_0__12124_ vdd gnd FILL
X_14319_ _14319_/A _14319_/Y vdd gnd INVX1
XFILL_0__8711_ vdd gnd FILL
X_7250_ _7250_/A _7250_/B _7250_/C _7250_/Y vdd gnd NAND3X1
XFILL_0__9691_ vdd gnd FILL
XFILL_2__9627_ vdd gnd FILL
XFILL_1__13414_ vdd gnd FILL
XFILL_1__10626_ vdd gnd FILL
XFILL_2__12965_ vdd gnd FILL
XFILL_1__14394_ vdd gnd FILL
XFILL_0__12055_ vdd gnd FILL
XFILL_0__8642_ vdd gnd FILL
X_7181_ _7181_/A _7181_/B _7181_/C _7181_/Y vdd gnd OAI21X1
XFILL_0__11006_ vdd gnd FILL
XFILL_2__9558_ vdd gnd FILL
XFILL_1__13345_ vdd gnd FILL
XFILL_1__10557_ vdd gnd FILL
XFILL_0__8573_ vdd gnd FILL
XFILL_2__9489_ vdd gnd FILL
XFILL_1__13276_ vdd gnd FILL
XFILL_0__7524_ vdd gnd FILL
XFILL_1__10488_ vdd gnd FILL
XFILL_1__12227_ vdd gnd FILL
XFILL_0__12957_ vdd gnd FILL
XFILL_0__7455_ vdd gnd FILL
XFILL_1_BUFX2_insert8 vdd gnd FILL
XFILL_0__11908_ vdd gnd FILL
XFILL_2__14497_ vdd gnd FILL
XFILL_1__12158_ vdd gnd FILL
XFILL_0__12888_ vdd gnd FILL
X_9822_ _9822_/D _9822_/CLK _9822_/Q vdd gnd DFFPOSX1
XFILL_0__7386_ vdd gnd FILL
XFILL_1__11109_ vdd gnd FILL
XFILL_0__14627_ vdd gnd FILL
XFILL_0__9125_ vdd gnd FILL
XFILL_1__12089_ vdd gnd FILL
XFILL_0__11839_ vdd gnd FILL
X_9753_ _9753_/A _9753_/B _9753_/C _9753_/Y vdd gnd OAI21X1
XFILL_2__13379_ vdd gnd FILL
XFILL_0__14558_ vdd gnd FILL
XFILL_0__9056_ vdd gnd FILL
X_8704_ _8704_/A _8704_/B _8704_/C _8704_/Y vdd gnd OAI21X1
X_9684_ _9684_/A _9684_/B _9684_/C _9684_/Y vdd gnd OAI21X1
XFILL_0__13509_ vdd gnd FILL
XFILL_0__8007_ vdd gnd FILL
XFILL_0__14489_ vdd gnd FILL
X_8635_ _8635_/A _8635_/B _8635_/C _8635_/Y vdd gnd OAI21X1
XFILL_1__8820_ vdd gnd FILL
X_8566_ _8566_/A _8566_/B _8566_/C _8566_/Y vdd gnd OAI21X1
X_7517_ _7517_/A _7517_/B _7517_/Y vdd gnd OR2X2
XFILL_0__9958_ vdd gnd FILL
XFILL_1__8751_ vdd gnd FILL
X_8497_ _8497_/A _8497_/B _8497_/C _8497_/Y vdd gnd NAND3X1
XFILL_1__7702_ vdd gnd FILL
X_7448_ _7448_/A _7448_/B _7448_/Y vdd gnd NAND2X1
XFILL_0__9889_ vdd gnd FILL
XFILL_1__8682_ vdd gnd FILL
XFILL256650x136950 vdd gnd FILL
XFILL_1__7633_ vdd gnd FILL
X_7379_ _7379_/A _7379_/B _7379_/C _7379_/Y vdd gnd NOR3X1
X_9118_ _9118_/A _9118_/B _9118_/C _9118_/Y vdd gnd OAI21X1
XFILL_1__7564_ vdd gnd FILL
X_10000_ _10000_/A _10000_/Y vdd gnd INVX2
XFILL_1__9303_ vdd gnd FILL
X_9049_ _9049_/A _9049_/B _9049_/Y vdd gnd OR2X2
XFILL_1__7495_ vdd gnd FILL
XFILL_1__9234_ vdd gnd FILL
XFILL_1__9165_ vdd gnd FILL
X_11951_ _11951_/A _11951_/B _11951_/Y vdd gnd NOR2X1
XFILL_1__8116_ vdd gnd FILL
X_10902_ _10902_/A _10902_/B _10902_/C _10902_/Y vdd gnd OAI21X1
X_14670_ _14670_/A _14670_/B _14670_/C _14670_/Y vdd gnd OAI21X1
X_11882_ _11882_/A _11882_/B _11882_/Y vdd gnd NAND2X1
XFILL_1__9096_ vdd gnd FILL
X_13621_ _13621_/A _13621_/B _13621_/Y vdd gnd NAND2X1
X_10833_ _10833_/A _10833_/Y vdd gnd INVX1
XFILL_1__8047_ vdd gnd FILL
X_10764_ _10764_/D _10764_/CLK _10764_/Q vdd gnd DFFPOSX1
X_13552_ _13552_/A _13552_/B _13552_/Y vdd gnd NAND2X1
X_12503_ _12503_/A _12503_/B _12503_/C _12503_/Y vdd gnd OAI21X1
X_13483_ _13483_/D _13483_/CLK _13483_/Q vdd gnd DFFPOSX1
X_10695_ _10695_/D _10695_/CLK _10695_/Q vdd gnd DFFPOSX1
XFILL_1__9998_ vdd gnd FILL
XFILL_2__8791_ vdd gnd FILL
X_12434_ _12434_/A _12434_/B _12434_/Y vdd gnd AND2X2
XFILL_1__8949_ vdd gnd FILL
XFILL_0__10170_ vdd gnd FILL
X_12365_ _12365_/A _12365_/B _12365_/Y vdd gnd AND2X2
XFILL_1__11460_ vdd gnd FILL
X_11316_ _11316_/A _11316_/B _11316_/Y vdd gnd NOR2X1
X_14104_ _14104_/A _14104_/B _14104_/Y vdd gnd NAND2X1
XFILL_2__9412_ vdd gnd FILL
X_12296_ _12296_/A _12296_/Y vdd gnd INVX1
XFILL_1__10411_ vdd gnd FILL
XFILL_2__12750_ vdd gnd FILL
XFILL_1__11391_ vdd gnd FILL
X_14035_ _14035_/A _14035_/B _14035_/C _14035_/Y vdd gnd AOI21X1
X_11247_ _11247_/A _11247_/Y vdd gnd INVX1
XFILL_1__13130_ vdd gnd FILL
XFILL_2__9343_ vdd gnd FILL
XFILL_1__10342_ vdd gnd FILL
XFILL_2__12681_ vdd gnd FILL
XFILL_0__13860_ vdd gnd FILL
X_11178_ _11178_/A _11178_/B _11178_/Y vdd gnd OR2X2
XFILL_2__9274_ vdd gnd FILL
XFILL_0__12811_ vdd gnd FILL
XFILL_1__13061_ vdd gnd FILL
XFILL_1__10273_ vdd gnd FILL
X_10129_ _10129_/A _10129_/B _10129_/C _10129_/Y vdd gnd OAI21X1
XFILL_0__13791_ vdd gnd FILL
XFILL_1__12012_ vdd gnd FILL
XFILL_2__14351_ vdd gnd FILL
XFILL_2__11563_ vdd gnd FILL
XFILL_0__12742_ vdd gnd FILL
XFILL_0__7240_ vdd gnd FILL
XFILL_2__14282_ vdd gnd FILL
XFILL_2__11494_ vdd gnd FILL
XFILL_0__12673_ vdd gnd FILL
XFILL_0__7171_ vdd gnd FILL
XFILL_2__7107_ vdd gnd FILL
X_14868_ _14868_/A _14868_/B _14868_/Y vdd gnd NOR2X1
XFILL_0__14412_ vdd gnd FILL
XFILL256650x201750 vdd gnd FILL
XFILL_1__13963_ vdd gnd FILL
X_13819_ _13819_/A _13819_/B _13819_/Y vdd gnd NAND2X1
XFILL_1__12914_ vdd gnd FILL
X_14799_ _14799_/A _14799_/B _14799_/C _14799_/Y vdd gnd AOI21X1
XFILL_0__14343_ vdd gnd FILL
XFILL_1__13894_ vdd gnd FILL
XFILL_0__11555_ vdd gnd FILL
XFILL_2__12115_ vdd gnd FILL
XFILL_0__10506_ vdd gnd FILL
XFILL_1__12845_ vdd gnd FILL
XFILL_0__14274_ vdd gnd FILL
X_8420_ _8420_/A _8420_/Y vdd gnd INVX1
XFILL_0__11486_ vdd gnd FILL
XFILL_2__12046_ vdd gnd FILL
XFILL_0__13225_ vdd gnd FILL
XFILL_0__10437_ vdd gnd FILL
XFILL_1__12776_ vdd gnd FILL
X_8351_ _8351_/A _8351_/B _8351_/Y vdd gnd NAND2X1
XFILL_1__11727_ vdd gnd FILL
XFILL_0__13156_ vdd gnd FILL
XFILL_0__10368_ vdd gnd FILL
X_7302_ _7302_/A _7302_/B _7302_/C _7302_/Y vdd gnd AOI21X1
XFILL_0__9743_ vdd gnd FILL
X_8282_ _8282_/A _8282_/B _8282_/C _8282_/Y vdd gnd NAND3X1
XFILL_1__14446_ vdd gnd FILL
XFILL_0__12107_ vdd gnd FILL
XFILL_0__13087_ vdd gnd FILL
XFILL_0__10299_ vdd gnd FILL
XFILL_2__13997_ vdd gnd FILL
X_7233_ _7233_/A _7233_/B _7233_/C _7233_/Y vdd gnd OAI21X1
XFILL_0__9674_ vdd gnd FILL
XFILL_1__10609_ vdd gnd FILL
XFILL_2__12948_ vdd gnd FILL
XFILL_0__12038_ vdd gnd FILL
XFILL_1__14377_ vdd gnd FILL
XFILL_1__11589_ vdd gnd FILL
XFILL_0__8625_ vdd gnd FILL
X_7164_ _7164_/A _7164_/B _7164_/Y vdd gnd NAND2X1
XFILL_1__13328_ vdd gnd FILL
XFILL_2__12879_ vdd gnd FILL
XFILL_0__8556_ vdd gnd FILL
X_7095_ _7095_/A _7095_/B _7095_/Y vdd gnd NAND2X1
XFILL_1__13259_ vdd gnd FILL
XFILL_0__7507_ vdd gnd FILL
XFILL_0__13989_ vdd gnd FILL
XFILL_1__7280_ vdd gnd FILL
XFILL_0__8487_ vdd gnd FILL
XFILL_0__7438_ vdd gnd FILL
X_9805_ _9805_/D _9805_/CLK _9805_/Q vdd gnd DFFPOSX1
XFILL_0__7369_ vdd gnd FILL
XFILL256650x111750 vdd gnd FILL
X_7997_ _7997_/A _7997_/Y vdd gnd INVX2
XFILL_0__9108_ vdd gnd FILL
X_9736_ _9736_/A _9736_/B _9736_/Y vdd gnd NAND2X1
XFILL_0__9039_ vdd gnd FILL
XFILL_1__9921_ vdd gnd FILL
XBUFX2_insert109 BUFX2_insert109/A BUFX2_insert109/Y vdd gnd BUFX2
X_9667_ _9667_/A _9667_/B _9667_/C _9667_/Y vdd gnd NAND3X1
X_8618_ _8618_/A _8618_/Y vdd gnd INVX1
XFILL_1__9852_ vdd gnd FILL
X_9598_ _9598_/A _9598_/B _9598_/C _9598_/Y vdd gnd OAI21X1
X_10480_ _10480_/A _10480_/Y vdd gnd INVX1
XFILL_1__8803_ vdd gnd FILL
X_8549_ _8549_/A _8549_/B _8549_/C _8549_/Y vdd gnd OAI21X1
XFILL_1__8734_ vdd gnd FILL
X_12150_ _12150_/A _12150_/B _12150_/Y vdd gnd NAND2X1
XFILL_1__8665_ vdd gnd FILL
X_11101_ _11101_/A _11101_/B _11101_/Y vdd gnd NAND2X1
X_12081_ _12081_/A _12081_/B _12081_/Y vdd gnd NAND2X1
XFILL_1__7616_ vdd gnd FILL
XFILL_1__8596_ vdd gnd FILL
X_11032_ _11032_/A _11032_/B _11032_/C _11032_/Y vdd gnd OAI21X1
XFILL_1__7547_ vdd gnd FILL
XFILL257550x176550 vdd gnd FILL
XFILL_1__7478_ vdd gnd FILL
XFILL_2__8010_ vdd gnd FILL
XFILL_1__9217_ vdd gnd FILL
X_12983_ _12983_/A _12983_/B _12983_/C _12983_/Y vdd gnd OAI21X1
X_14722_ _14722_/A _14722_/B _14722_/C _14722_/Y vdd gnd OAI21X1
X_11934_ _11934_/A _11934_/B _11934_/C _11934_/Y vdd gnd AOI21X1
XFILL_1__9148_ vdd gnd FILL
X_14653_ _14653_/A _14653_/B _14653_/Y vdd gnd NOR2X1
XFILL_1__9079_ vdd gnd FILL
X_11865_ _11865_/A _11865_/B _11865_/C _11865_/Y vdd gnd OAI21X1
XFILL_1__10960_ vdd gnd FILL
X_13604_ _13604_/A _13604_/B _13604_/S _13604_/Y vdd gnd MUX2X1
X_10816_ _10816_/A _10816_/B _10816_/C _10816_/Y vdd gnd OAI21X1
X_14584_ _14584_/A _14584_/B _14584_/C _14584_/Y vdd gnd OAI21X1
X_11796_ _11796_/A _11796_/B _11796_/Y vdd gnd NAND2X1
XFILL_0__11340_ vdd gnd FILL
XFILL257250x90150 vdd gnd FILL
XFILL_1__10891_ vdd gnd FILL
X_13535_ _13535_/A _13535_/B _13535_/C _13535_/D _13535_/Y vdd gnd AOI22X1
X_10747_ _10747_/D _10747_/CLK _10747_/Q vdd gnd DFFPOSX1
XFILL_1__12630_ vdd gnd FILL
XFILL_0__11271_ vdd gnd FILL
X_10678_ _10678_/A _10678_/B _10678_/Y vdd gnd NAND2X1
X_13466_ _13466_/D _13466_/CLK _13466_/Q vdd gnd DFFPOSX1
XFILL_0__13010_ vdd gnd FILL
XFILL_2__13920_ vdd gnd FILL
XFILL_0__10222_ vdd gnd FILL
X_12417_ _12417_/A _12417_/B _12417_/C _12417_/Y vdd gnd NAND3X1
XFILL_1__14300_ vdd gnd FILL
XFILL_2__7725_ vdd gnd FILL
XFILL_1__11512_ vdd gnd FILL
X_13397_ _13397_/A _13397_/B _13397_/C _13397_/Y vdd gnd OAI21X1
XFILL_2__13851_ vdd gnd FILL
XFILL_0__10153_ vdd gnd FILL
XFILL_1__12492_ vdd gnd FILL
X_12348_ _12348_/A _12348_/B _12348_/C _12348_/Y vdd gnd OAI21X1
XFILL_1__14231_ vdd gnd FILL
XFILL_2__7656_ vdd gnd FILL
XFILL_1__11443_ vdd gnd FILL
XFILL_0__10084_ vdd gnd FILL
XFILL_2__13782_ vdd gnd FILL
X_12279_ _12279_/A _12279_/B _12279_/C _12279_/Y vdd gnd OAI21X1
XFILL_0__13912_ vdd gnd FILL
XFILL_2__12733_ vdd gnd FILL
XFILL_1__11374_ vdd gnd FILL
XFILL_0__8410_ vdd gnd FILL
X_14018_ _14018_/A _14018_/B _14018_/C _14018_/Y vdd gnd OAI21X1
XFILL_0__9390_ vdd gnd FILL
XFILL_1__13113_ vdd gnd FILL
XFILL_2__9326_ vdd gnd FILL
XFILL_1__10325_ vdd gnd FILL
XFILL_2__12664_ vdd gnd FILL
XFILL_0__13843_ vdd gnd FILL
XFILL_1__14093_ vdd gnd FILL
XFILL_0__8341_ vdd gnd FILL
XFILL_2__9257_ vdd gnd FILL
XFILL_1__13044_ vdd gnd FILL
XFILL_1__10256_ vdd gnd FILL
XFILL_0__13774_ vdd gnd FILL
XFILL_0__10986_ vdd gnd FILL
X_7920_ _7920_/D _7920_/CLK _7920_/Q vdd gnd DFFPOSX1
XFILL_0__8272_ vdd gnd FILL
XFILL_2__11546_ vdd gnd FILL
XFILL_2__9188_ vdd gnd FILL
XFILL_0__12725_ vdd gnd FILL
XFILL_0__7223_ vdd gnd FILL
XFILL_1__10187_ vdd gnd FILL
X_7851_ _7851_/A _7851_/B _7851_/Y vdd gnd AND2X2
XFILL_2__11477_ vdd gnd FILL
XFILL_0__12656_ vdd gnd FILL
XFILL_0__7154_ vdd gnd FILL
X_7782_ _7782_/A _7782_/B _7782_/Y vdd gnd NAND2X1
XFILL_0__11607_ vdd gnd FILL
XFILL_1__13946_ vdd gnd FILL
X_9521_ _9521_/A _9521_/B _9521_/Y vdd gnd NOR2X1
XFILL_0__7085_ vdd gnd FILL
XFILL_0__14326_ vdd gnd FILL
XFILL_0__11538_ vdd gnd FILL
XFILL_1__13877_ vdd gnd FILL
X_9452_ _9452_/A _9452_/B _9452_/C _9452_/Y vdd gnd OAI21X1
XFILL257550x241350 vdd gnd FILL
XFILL_0__14257_ vdd gnd FILL
XFILL_1__12828_ vdd gnd FILL
X_8403_ _8403_/A _8403_/B _8403_/C _8403_/Y vdd gnd NAND3X1
XFILL_0__11469_ vdd gnd FILL
X_9383_ _9383_/A _9383_/B _9383_/C _9383_/Y vdd gnd OAI21X1
XFILL_2__12029_ vdd gnd FILL
XFILL_0__13208_ vdd gnd FILL
XFILL_1__12759_ vdd gnd FILL
X_8334_ _8334_/A _8334_/B _8334_/C _8334_/Y vdd gnd NAND3X1
XFILL_0__13139_ vdd gnd FILL
XFILL_0__9726_ vdd gnd FILL
X_8265_ _8265_/A _8265_/B _8265_/C _8265_/Y vdd gnd NAND3X1
XFILL_1__14429_ vdd gnd FILL
X_7216_ _7216_/A _7216_/B _7216_/Y vdd gnd NAND2X1
XFILL_0__9657_ vdd gnd FILL
XFILL_1__8450_ vdd gnd FILL
X_8196_ _8196_/A _8196_/B _8196_/Y vdd gnd NOR2X1
XFILL_1__7401_ vdd gnd FILL
XFILL_0__8608_ vdd gnd FILL
X_7147_ _7147_/A _7147_/B _7147_/S _7147_/Y vdd gnd MUX2X1
XFILL_1__8381_ vdd gnd FILL
XFILL_0__9588_ vdd gnd FILL
XFILL_1__7332_ vdd gnd FILL
XFILL_0__8539_ vdd gnd FILL
X_7078_ _7078_/A _7078_/B _7078_/Y vdd gnd NOR2X1
XFILL_1__7263_ vdd gnd FILL
XFILL257550x108150 vdd gnd FILL
XFILL_1__9002_ vdd gnd FILL
XFILL_1__7194_ vdd gnd FILL
X_11650_ _11650_/D _11650_/CLK _11650_/Q vdd gnd DFFPOSX1
X_9719_ _9719_/A _9719_/Y vdd gnd INVX1
X_10601_ _10601_/A _10601_/B _10601_/Y vdd gnd NAND2X1
XFILL_1__9904_ vdd gnd FILL
X_11581_ _11581_/A _11581_/B _11581_/C _11581_/Y vdd gnd OAI21X1
XFILL257550x151350 vdd gnd FILL
X_10532_ _10532_/A _10532_/B _10532_/Y vdd gnd NAND2X1
X_13320_ _13320_/A _13320_/B _13320_/Y vdd gnd NOR2X1
X_10463_ _10463_/A _10463_/B _10463_/Y vdd gnd NAND2X1
X_13251_ _13251_/A _13251_/B _13251_/Y vdd gnd NAND2X1
X_12202_ _12202_/A _12202_/B _12202_/Y vdd gnd NAND2X1
X_13182_ _13182_/A _13182_/B _13182_/Y vdd gnd NAND2X1
X_10394_ _10394_/A _10394_/Y vdd gnd INVX1
XFILL_2__7510_ vdd gnd FILL
XFILL_1__8717_ vdd gnd FILL
XFILL_1__9697_ vdd gnd FILL
X_12133_ _12133_/A _12133_/B _12133_/Y vdd gnd NOR2X1
XFILL_2__7441_ vdd gnd FILL
XFILL_1__8648_ vdd gnd FILL
X_12064_ _12064_/A _12064_/B _12064_/C _12064_/Y vdd gnd OAI21X1
XFILL_2__7372_ vdd gnd FILL
XFILL_1__8579_ vdd gnd FILL
X_11015_ _11015_/A _11015_/B _11015_/C _11015_/Y vdd gnd OAI21X1
XFILL_1__10110_ vdd gnd FILL
XFILL_0__10840_ vdd gnd FILL
XFILL_1__11090_ vdd gnd FILL
XFILL_1__10041_ vdd gnd FILL
XFILL_0__10771_ vdd gnd FILL
XBUFX2_insert9 BUFX2_insert9/A BUFX2_insert9/Y vdd gnd BUFX2
X_12966_ _12966_/A _12966_/B _12966_/C _12966_/Y vdd gnd NOR3X1
XFILL_0__12510_ vdd gnd FILL
X_14705_ _14705_/A _14705_/B _14705_/Y vdd gnd NAND2X1
X_11917_ _11917_/A _11917_/B _11917_/C _11917_/Y vdd gnd OAI21X1
X_12897_ _12897_/A _12897_/Y vdd gnd INVX1
XFILL_1__13800_ vdd gnd FILL
XFILL_1__14780_ vdd gnd FILL
XFILL_0__12441_ vdd gnd FILL
XFILL_1__11992_ vdd gnd FILL
X_14636_ _14636_/A _14636_/Y vdd gnd INVX1
XFILL_2__10213_ vdd gnd FILL
X_11848_ _11848_/A _11848_/Y vdd gnd INVX2
XFILL_1__13731_ vdd gnd FILL
XFILL_1__10943_ vdd gnd FILL
XFILL_0__12372_ vdd gnd FILL
X_14567_ _14567_/A _14567_/B _14567_/C _14567_/Y vdd gnd OAI21X1
XFILL_2__10144_ vdd gnd FILL
X_11779_ _11779_/A _11779_/B _11779_/Y vdd gnd NOR2X1
XFILL_0__14111_ vdd gnd FILL
XFILL_1__13662_ vdd gnd FILL
XFILL_0__11323_ vdd gnd FILL
XFILL_1__10874_ vdd gnd FILL
XFILL_0__7910_ vdd gnd FILL
X_13518_ _13518_/A _13518_/B _13518_/Y vdd gnd NAND2X1
X_14498_ _14498_/A _14498_/B _14498_/Y vdd gnd NAND2X1
XFILL_2__10075_ vdd gnd FILL
XFILL_0__14042_ vdd gnd FILL
XFILL_1__13593_ vdd gnd FILL
XFILL_0__11254_ vdd gnd FILL
X_13449_ _13449_/D _13449_/CLK _13449_/Q vdd gnd DFFPOSX1
XFILL_0__7841_ vdd gnd FILL
XFILL_0__10205_ vdd gnd FILL
XFILL_0__11185_ vdd gnd FILL
XFILL_0__7772_ vdd gnd FILL
XFILL_2__7708_ vdd gnd FILL
XFILL_0__10136_ vdd gnd FILL
XFILL_1__12475_ vdd gnd FILL
XFILL_0__9511_ vdd gnd FILL
X_8050_ _8050_/A _8050_/B _8050_/C _8050_/D _8050_/Y vdd gnd AOI22X1
XFILL_2__7639_ vdd gnd FILL
XFILL_1__11426_ vdd gnd FILL
XFILL_2__13765_ vdd gnd FILL
XFILL_2__10977_ vdd gnd FILL
XFILL_0__10067_ vdd gnd FILL
XFILL_0__9442_ vdd gnd FILL
XFILL_1_BUFX2_insert13 vdd gnd FILL
XFILL_1_BUFX2_insert24 vdd gnd FILL
XFILL_1__14145_ vdd gnd FILL
XFILL_1__11357_ vdd gnd FILL
XFILL_2__13696_ vdd gnd FILL
XFILL_0__9373_ vdd gnd FILL
XFILL_1__10308_ vdd gnd FILL
XFILL_1__14076_ vdd gnd FILL
XFILL_0__13826_ vdd gnd FILL
XFILL_1__11288_ vdd gnd FILL
XFILL_0__8324_ vdd gnd FILL
X_8952_ _8952_/A _8952_/B _8952_/Y vdd gnd NAND2X1
XFILL_1__13027_ vdd gnd FILL
XFILL_1__10239_ vdd gnd FILL
XFILL_0__13757_ vdd gnd FILL
XFILL_0__10969_ vdd gnd FILL
X_7903_ _7903_/A _7903_/B _7903_/C _7903_/Y vdd gnd OAI21X1
XFILL_0__8255_ vdd gnd FILL
X_8883_ _8883_/D _8883_/CLK _8883_/Q vdd gnd DFFPOSX1
XFILL_0__12708_ vdd gnd FILL
XFILL_0__7206_ vdd gnd FILL
XFILL_0__13688_ vdd gnd FILL
X_7834_ _7834_/A _7834_/B _7834_/Y vdd gnd NOR2X1
XFILL_0__8186_ vdd gnd FILL
XFILL_0__12639_ vdd gnd FILL
XFILL_0__7137_ vdd gnd FILL
XFILL_1_CLKBUF1_insert36 vdd gnd FILL
X_7765_ _7765_/A _7765_/B _7765_/C _7765_/Y vdd gnd OAI21X1
XFILL_1_CLKBUF1_insert47 vdd gnd FILL
XFILL_1_CLKBUF1_insert58 vdd gnd FILL
XFILL_1__13929_ vdd gnd FILL
XFILL_1_CLKBUF1_insert69 vdd gnd FILL
X_9504_ _9504_/A _9504_/B _9504_/C _9504_/Y vdd gnd AOI21X1
X_7696_ _7696_/A _7696_/B _7696_/C _7696_/Y vdd gnd AOI21X1
XFILL_0__14309_ vdd gnd FILL
X_9435_ _9435_/A _9435_/B _9435_/C _9435_/Y vdd gnd OAI21X1
XFILL_1__7881_ vdd gnd FILL
XFILL_1__9620_ vdd gnd FILL
X_9366_ _9366_/A _9366_/B _9366_/C _9366_/Y vdd gnd OAI21X1
X_8317_ _8317_/A _8317_/B _8317_/C _8317_/Y vdd gnd OAI21X1
XFILL_1__9551_ vdd gnd FILL
X_9297_ _9297_/A _9297_/B _9297_/Y vdd gnd AND2X2
XFILL_0__9709_ vdd gnd FILL
XFILL_1__8502_ vdd gnd FILL
X_8248_ _8248_/A _8248_/B _8248_/C _8248_/Y vdd gnd NAND3X1
XFILL_1__9482_ vdd gnd FILL
XFILL_1__8433_ vdd gnd FILL
X_8179_ _8179_/A _8179_/B _8179_/C _8179_/Y vdd gnd OAI21X1
XFILL_1__8364_ vdd gnd FILL
XFILL_1__7315_ vdd gnd FILL
XFILL_1__8295_ vdd gnd FILL
X_12820_ _12820_/A _12820_/Y vdd gnd INVX1
XFILL_1__7246_ vdd gnd FILL
X_12751_ _12751_/A _12751_/B _12751_/C _12751_/Y vdd gnd AOI21X1
XFILL_1__7177_ vdd gnd FILL
X_11702_ _11702_/A _11702_/B _11702_/C _11702_/D _11702_/Y vdd gnd AOI22X1
X_12682_ _12682_/A _12682_/B _12682_/Y vdd gnd NAND2X1
X_14421_ _14421_/A _14421_/Y vdd gnd INVX1
X_11633_ _11633_/D _11633_/CLK _11633_/Q vdd gnd DFFPOSX1
X_14352_ _14352_/A _14352_/Y vdd gnd INVX1
X_11564_ _11564_/A _11564_/Y vdd gnd INVX1
XFILL_2__9660_ vdd gnd FILL
X_13303_ _13303_/A _13303_/B _13303_/Y vdd gnd NAND2X1
X_10515_ _10515_/A _10515_/B _10515_/Y vdd gnd NAND2X1
X_14283_ _14283_/A _14283_/B _14283_/Y vdd gnd NAND2X1
X_11495_ _11495_/A _11495_/B _11495_/C _11495_/Y vdd gnd AOI21X1
XFILL_2__9591_ vdd gnd FILL
XFILL_1__10590_ vdd gnd FILL
X_10446_ _10446_/A _10446_/B _10446_/C _10446_/D _10446_/Y vdd gnd AOI22X1
X_13234_ _13234_/A _13234_/B _13234_/C _13234_/Y vdd gnd OAI21X1
XFILL_1__9749_ vdd gnd FILL
XFILL_2__10900_ vdd gnd FILL
X_13165_ _13165_/A _13165_/B _13165_/C _13165_/Y vdd gnd OAI21X1
X_10377_ _10377_/A _10377_/B _10377_/C _10377_/Y vdd gnd NAND3X1
XFILL_1__12260_ vdd gnd FILL
XFILL_2__10831_ vdd gnd FILL
X_12116_ _12116_/A _12116_/Y vdd gnd INVX1
XFILL_0__12990_ vdd gnd FILL
X_13096_ _13096_/A _13096_/B _13096_/C _13096_/Y vdd gnd NAND3X1
XFILL_1__11211_ vdd gnd FILL
XFILL_2__7424_ vdd gnd FILL
XFILL_0__11941_ vdd gnd FILL
XFILL_1__12191_ vdd gnd FILL
X_12047_ _12047_/A _12047_/B _12047_/Y vdd gnd NAND2X1
XFILL_2__12501_ vdd gnd FILL
XFILL_2__7355_ vdd gnd FILL
XFILL_1__11142_ vdd gnd FILL
XFILL_0__14660_ vdd gnd FILL
XFILL_0__11872_ vdd gnd FILL
XFILL_0__13611_ vdd gnd FILL
XFILL_2__12432_ vdd gnd FILL
XFILL_1__11073_ vdd gnd FILL
XFILL_2__7286_ vdd gnd FILL
XFILL_0__10823_ vdd gnd FILL
XFILL_0__14591_ vdd gnd FILL
XFILL_2_BUFX2_insert260 vdd gnd FILL
XFILL_1__10024_ vdd gnd FILL
XFILL_2__12363_ vdd gnd FILL
X_13998_ _13998_/A _13998_/B _13998_/Y vdd gnd NAND2X1
XFILL_0__13542_ vdd gnd FILL
XFILL_0__8040_ vdd gnd FILL
XFILL_2_BUFX2_insert282 vdd gnd FILL
X_12949_ _12949_/A _12949_/B _12949_/Y vdd gnd AND2X2
XFILL_1__14832_ vdd gnd FILL
XFILL_2__12294_ vdd gnd FILL
XFILL_0__10685_ vdd gnd FILL
XFILL_0__12424_ vdd gnd FILL
XFILL_1__14763_ vdd gnd FILL
XFILL_1__11975_ vdd gnd FILL
X_14619_ _14619_/A _14619_/B _14619_/Y vdd gnd NOR2X1
X_7550_ _7550_/A _7550_/B _7550_/C _7550_/D _7550_/Y vdd gnd AOI22X1
XFILL_0__9991_ vdd gnd FILL
XFILL_1__10926_ vdd gnd FILL
XFILL_1__13714_ vdd gnd FILL
XFILL_0__12355_ vdd gnd FILL
XFILL_1__14694_ vdd gnd FILL
XFILL_0__8942_ vdd gnd FILL
X_7481_ _7481_/A _7481_/B _7481_/Y vdd gnd NAND2X1
XFILL_2__10127_ vdd gnd FILL
XBUFX2_insert270 BUFX2_insert270/A BUFX2_insert270/Y vdd gnd BUFX2
XFILL_0__11306_ vdd gnd FILL
XFILL_1__13645_ vdd gnd FILL
XBUFX2_insert281 BUFX2_insert281/A BUFX2_insert281/Y vdd gnd BUFX2
XFILL_1__10857_ vdd gnd FILL
X_9220_ _9220_/A _9220_/B _9220_/Y vdd gnd AND2X2
XFILL_0__12286_ vdd gnd FILL
XBUFX2_insert292 BUFX2_insert292/A BUFX2_insert292/Y vdd gnd BUFX2
XFILL_2__10058_ vdd gnd FILL
XFILL_0__14025_ vdd gnd FILL
XFILL_0__11237_ vdd gnd FILL
XFILL_1__13576_ vdd gnd FILL
XFILL_1__10788_ vdd gnd FILL
X_9151_ _9151_/A _9151_/B _9151_/Y vdd gnd NAND2X1
XFILL_0__7824_ vdd gnd FILL
XFILL_1__12527_ vdd gnd FILL
XFILL_0__11168_ vdd gnd FILL
X_8102_ _8102_/A _8102_/B _8102_/S _8102_/Y vdd gnd MUX2X1
X_9082_ _9082_/A _9082_/Y vdd gnd INVX1
XFILL_0__7755_ vdd gnd FILL
XFILL_0__10119_ vdd gnd FILL
XFILL_1__12458_ vdd gnd FILL
X_8033_ _8033_/A _8033_/B _8033_/Y vdd gnd NAND2X1
XFILL_0__11099_ vdd gnd FILL
XFILL_0__7686_ vdd gnd FILL
XFILL_1__11409_ vdd gnd FILL
XFILL_1__12389_ vdd gnd FILL
XFILL_0__9425_ vdd gnd FILL
XFILL_1__14128_ vdd gnd FILL
XFILL_0__14858_ vdd gnd FILL
XFILL_0__9356_ vdd gnd FILL
X_9984_ _9984_/A _9984_/B _9984_/Y vdd gnd NAND2X1
XFILL_1__14059_ vdd gnd FILL
XFILL_0__13809_ vdd gnd FILL
XFILL_1__7100_ vdd gnd FILL
XFILL_0__14789_ vdd gnd FILL
XFILL_0__8307_ vdd gnd FILL
XFILL_1__8080_ vdd gnd FILL
XFILL_0__9287_ vdd gnd FILL
X_8935_ _8935_/A _8935_/Y vdd gnd INVX1
XFILL_0__8238_ vdd gnd FILL
X_8866_ _8866_/D _8866_/CLK _8866_/Q vdd gnd DFFPOSX1
X_7817_ _7817_/A _7817_/B _7817_/Y vdd gnd NAND2X1
XFILL_0__8169_ vdd gnd FILL
X_8797_ _8797_/A _8797_/B _8797_/C _8797_/Y vdd gnd OAI21X1
X_7748_ _7748_/A _7748_/B _7748_/C _7748_/Y vdd gnd OAI21X1
XFILL_1__8982_ vdd gnd FILL
X_7679_ _7679_/A _7679_/B _7679_/Y vdd gnd NOR2X1
X_9418_ _9418_/A _9418_/B _9418_/C _9418_/Y vdd gnd OAI21X1
XFILL_1__7864_ vdd gnd FILL
X_10300_ _10300_/A _10300_/B _10300_/C _10300_/D _10300_/Y vdd gnd AOI22X1
XFILL_1__9603_ vdd gnd FILL
X_11280_ _11280_/A _11280_/B _11280_/Y vdd gnd NAND2X1
X_9349_ _9349_/A _9349_/Y vdd gnd INVX1
XFILL_1__7795_ vdd gnd FILL
X_10231_ _10231_/A _10231_/B _10231_/Y vdd gnd NAND2X1
XFILL_1__9534_ vdd gnd FILL
X_10162_ _10162_/A _10162_/B _10162_/Y vdd gnd AND2X2
XFILL_1__9465_ vdd gnd FILL
X_10093_ _10093_/A _10093_/Y vdd gnd INVX1
XFILL_1__8416_ vdd gnd FILL
XFILL_1__9396_ vdd gnd FILL
X_13921_ _13921_/A _13921_/B _13921_/C _13921_/Y vdd gnd OAI21X1
XFILL_1__8347_ vdd gnd FILL
X_13852_ _13852_/A _13852_/B _13852_/Y vdd gnd NAND2X1
XFILL_1__8278_ vdd gnd FILL
X_12803_ _12803_/A _12803_/Y vdd gnd INVX2
XFILL_1_BUFX2_insert201 vdd gnd FILL
XFILL_1__7229_ vdd gnd FILL
XFILL_1_BUFX2_insert212 vdd gnd FILL
X_13783_ _13783_/A _13783_/B _13783_/C _13783_/Y vdd gnd OAI21X1
X_10995_ _10995_/A _10995_/Y vdd gnd INVX1
XFILL_1_BUFX2_insert223 vdd gnd FILL
XFILL_1_BUFX2_insert234 vdd gnd FILL
XFILL_1_BUFX2_insert245 vdd gnd FILL
X_12734_ _12734_/A _12734_/Y vdd gnd INVX1
XFILL_1_BUFX2_insert256 vdd gnd FILL
XFILL_1_BUFX2_insert267 vdd gnd FILL
XFILL_1_BUFX2_insert278 vdd gnd FILL
XFILL_0__10470_ vdd gnd FILL
XCLKBUF1_insert38 CLKBUF1_insert38/A CLKBUF1_insert38/Y vdd gnd CLKBUF1
XFILL_1_BUFX2_insert289 vdd gnd FILL
XCLKBUF1_insert49 CLKBUF1_insert49/A CLKBUF1_insert49/Y vdd gnd CLKBUF1
X_12665_ _12665_/A _12665_/B _12665_/C _12665_/D _12665_/Y vdd gnd AOI22X1
XFILL_1__11760_ vdd gnd FILL
X_14404_ _14404_/A _14404_/B _14404_/Y vdd gnd NAND2X1
X_11616_ _11616_/D _11616_/CLK _11616_/Q vdd gnd DFFPOSX1
X_12596_ _12596_/D _12596_/CLK _12596_/Q vdd gnd DFFPOSX1
XFILL_0__12140_ vdd gnd FILL
X_14335_ _14335_/A _14335_/Y vdd gnd INVX1
X_11547_ _11547_/A _11547_/B _11547_/Y vdd gnd AND2X2
XFILL_2__9643_ vdd gnd FILL
XFILL_1__10642_ vdd gnd FILL
XFILL_0__12071_ vdd gnd FILL
XFILL_2__12981_ vdd gnd FILL
X_14266_ _14266_/A _14266_/B _14266_/Y vdd gnd NOR2X1
XFILL_2__14720_ vdd gnd FILL
X_11478_ _11478_/A _11478_/B _11478_/Y vdd gnd NAND2X1
XFILL_0__11022_ vdd gnd FILL
XFILL_2__9574_ vdd gnd FILL
XFILL_1__13361_ vdd gnd FILL
XFILL_1__10573_ vdd gnd FILL
X_13217_ _13217_/A _13217_/B _13217_/C _13217_/Y vdd gnd AOI21X1
X_10429_ _10429_/A _10429_/B _10429_/Y vdd gnd NOR2X1
XFILL_1__12312_ vdd gnd FILL
X_14197_ _14197_/D _14197_/CLK _14197_/Q vdd gnd DFFPOSX1
XFILL_2__14651_ vdd gnd FILL
XFILL_1__13292_ vdd gnd FILL
X_13148_ _13148_/A _13148_/B _13148_/Y vdd gnd NAND2X1
XFILL_0__7540_ vdd gnd FILL
XFILL_1__12243_ vdd gnd FILL
XFILL_0__12973_ vdd gnd FILL
X_13079_ _13079_/A _13079_/B _13079_/C _13079_/Y vdd gnd NAND3X1
XFILL_0__7471_ vdd gnd FILL
XFILL_0__14712_ vdd gnd FILL
XFILL_0__11924_ vdd gnd FILL
XFILL_1__12174_ vdd gnd FILL
XFILL_0__9210_ vdd gnd FILL
XFILL_1__11125_ vdd gnd FILL
XFILL_0__14643_ vdd gnd FILL
XFILL_0__11855_ vdd gnd FILL
XFILL_0__9141_ vdd gnd FILL
XFILL_2__12415_ vdd gnd FILL
XFILL_1__11056_ vdd gnd FILL
XFILL_0__10806_ vdd gnd FILL
XFILL_0__14574_ vdd gnd FILL
XFILL_0__11786_ vdd gnd FILL
XFILL_0__9072_ vdd gnd FILL
X_8720_ _8720_/A _8720_/Y vdd gnd INVX1
XFILL_1__10007_ vdd gnd FILL
XFILL_2__12346_ vdd gnd FILL
XFILL_0__13525_ vdd gnd FILL
XFILL_0__8023_ vdd gnd FILL
X_8651_ _8651_/A _8651_/B _8651_/C _8651_/Y vdd gnd OAI21X1
XFILL_1__14815_ vdd gnd FILL
XFILL_2__12277_ vdd gnd FILL
X_7602_ _7602_/A _7602_/B _7602_/Y vdd gnd NOR2X1
XFILL_0__10668_ vdd gnd FILL
X_8582_ _8582_/A _8582_/B _8582_/C _8582_/Y vdd gnd NAND3X1
XFILL_2__14016_ vdd gnd FILL
XFILL_0__12407_ vdd gnd FILL
XFILL_1__14746_ vdd gnd FILL
XFILL_1__11958_ vdd gnd FILL
XFILL_0__13387_ vdd gnd FILL
X_7533_ _7533_/A _7533_/B _7533_/C _7533_/Y vdd gnd OAI21X1
XFILL_0__10599_ vdd gnd FILL
XFILL_0__9974_ vdd gnd FILL
XFILL_0__12338_ vdd gnd FILL
XFILL_1__10909_ vdd gnd FILL
XFILL_1__14677_ vdd gnd FILL
XFILL_0__8925_ vdd gnd FILL
XFILL_1__11889_ vdd gnd FILL
X_7464_ _7464_/A _7464_/B _7464_/Y vdd gnd NAND2X1
XFILL_1__13628_ vdd gnd FILL
XFILL_0__12269_ vdd gnd FILL
X_9203_ _9203_/A _9203_/Y vdd gnd INVX1
XFILL_0__14008_ vdd gnd FILL
X_7395_ _7395_/A _7395_/B _7395_/C _7395_/Y vdd gnd OAI21X1
XFILL_2__14918_ vdd gnd FILL
XFILL_1__13559_ vdd gnd FILL
X_9134_ _9134_/A _9134_/B _9134_/C _9134_/Y vdd gnd OAI21X1
XFILL_0__7807_ vdd gnd FILL
XFILL_1__7580_ vdd gnd FILL
XFILL_0__8787_ vdd gnd FILL
X_9065_ _9065_/A _9065_/Y vdd gnd INVX1
XFILL_0__7738_ vdd gnd FILL
X_8016_ _8016_/A _8016_/B _8016_/C _8016_/Y vdd gnd OAI21X1
XFILL_1__9250_ vdd gnd FILL
XFILL_0__7669_ vdd gnd FILL
XFILL_0__9408_ vdd gnd FILL
XFILL_1__8201_ vdd gnd FILL
XFILL_1__9181_ vdd gnd FILL
XFILL_0__9339_ vdd gnd FILL
XFILL_1__8132_ vdd gnd FILL
X_9967_ _9967_/A _9967_/B _9967_/C _9967_/Y vdd gnd OAI21X1
X_8918_ _8918_/D _8918_/CLK _8918_/Q vdd gnd DFFPOSX1
XFILL_1__8063_ vdd gnd FILL
X_9898_ _9898_/A _9898_/B _9898_/C _9898_/D _9898_/Y vdd gnd AOI22X1
X_10780_ _10780_/A _10780_/B _10780_/Y vdd gnd NOR2X1
X_8849_ _8849_/D _8849_/CLK _8849_/Q vdd gnd DFFPOSX1
XFILL_0_BUFX2_insert208 vdd gnd FILL
XFILL_0_BUFX2_insert219 vdd gnd FILL
X_12450_ _12450_/A _12450_/B _12450_/C _12450_/Y vdd gnd OAI21X1
XFILL_1__8965_ vdd gnd FILL
X_11401_ _11401_/A _11401_/B _11401_/Y vdd gnd NAND2X1
X_12381_ _12381_/A _12381_/B _12381_/C _12381_/D _12381_/Y vdd gnd OAI22X1
X_14120_ _14120_/A _14120_/B _14120_/C _14120_/Y vdd gnd OAI21X1
X_11332_ _11332_/A _11332_/B _11332_/Y vdd gnd OR2X2
XFILL_1__7847_ vdd gnd FILL
X_14051_ _14051_/A _14051_/B _14051_/C _14051_/Y vdd gnd OAI21X1
XFILL257250x187350 vdd gnd FILL
X_11263_ _11263_/A _11263_/B _11263_/Y vdd gnd NAND2X1
XFILL_1__7778_ vdd gnd FILL
X_13002_ _13002_/A _13002_/B _13002_/Y vdd gnd NAND2X1
X_10214_ _10214_/A _10214_/B _10214_/C _10214_/Y vdd gnd NAND3X1
XFILL_1__9517_ vdd gnd FILL
XFILL_2__8310_ vdd gnd FILL
X_11194_ _11194_/A _11194_/B _11194_/C _11194_/Y vdd gnd AOI21X1
X_10145_ _10145_/A _10145_/B _10145_/Y vdd gnd AND2X2
XFILL_1__9448_ vdd gnd FILL
XFILL_2__8241_ vdd gnd FILL
X_10076_ _10076_/A _10076_/B _10076_/C _10076_/Y vdd gnd OAI21X1
XFILL_2__10530_ vdd gnd FILL
XFILL_1__9379_ vdd gnd FILL
XFILL_2__8172_ vdd gnd FILL
X_13904_ _13904_/A _13904_/B _13904_/Y vdd gnd NAND2X1
X_14884_ _14884_/D _14884_/CLK _14884_/Q vdd gnd DFFPOSX1
XFILL_2__10461_ vdd gnd FILL
X_13835_ _13835_/A _13835_/Y vdd gnd INVX1
XFILL_1__12930_ vdd gnd FILL
XFILL_2__10392_ vdd gnd FILL
XFILL_0__11571_ vdd gnd FILL
X_13766_ _13766_/A _13766_/B _13766_/C _13766_/Y vdd gnd OAI21X1
X_10978_ _10978_/A _10978_/B _10978_/Y vdd gnd NAND2X1
XFILL_0__13310_ vdd gnd FILL
XFILL_0__10522_ vdd gnd FILL
XFILL256950x28950 vdd gnd FILL
XFILL_0__14290_ vdd gnd FILL
XFILL_1__12861_ vdd gnd FILL
X_12717_ _12717_/A _12717_/B _12717_/Y vdd gnd NAND2X1
XFILL_1__14600_ vdd gnd FILL
XFILL_2__12062_ vdd gnd FILL
X_13697_ _13697_/A _13697_/Y vdd gnd INVX1
XFILL_1__11812_ vdd gnd FILL
XFILL_0__13241_ vdd gnd FILL
XFILL_0__10453_ vdd gnd FILL
XFILL_1__12792_ vdd gnd FILL
X_12648_ _12648_/A _12648_/B _12648_/C _12648_/Y vdd gnd OAI21X1
XFILL_0__13172_ vdd gnd FILL
XFILL_1__11743_ vdd gnd FILL
XFILL_0__10384_ vdd gnd FILL
X_12579_ _12579_/D _12579_/CLK _12579_/Q vdd gnd DFFPOSX1
XFILL_0__12123_ vdd gnd FILL
XFILL_2__7887_ vdd gnd FILL
XFILL_1__14462_ vdd gnd FILL
X_14318_ _14318_/A _14318_/Y vdd gnd INVX1
XFILL_0__8710_ vdd gnd FILL
XFILL_0__9690_ vdd gnd FILL
XFILL_1__10625_ vdd gnd FILL
XFILL_1__13413_ vdd gnd FILL
XFILL_0__12054_ vdd gnd FILL
XFILL_1__14393_ vdd gnd FILL
X_14249_ _14249_/A _14249_/Y vdd gnd INVX1
XFILL_0__8641_ vdd gnd FILL
X_7180_ _7180_/A _7180_/B _7180_/Y vdd gnd NAND2X1
XFILL_2__14703_ vdd gnd FILL
XFILL_0__11005_ vdd gnd FILL
XFILL_2__11915_ vdd gnd FILL
XFILL_1__10556_ vdd gnd FILL
XFILL_1__13344_ vdd gnd FILL
XFILL_2__12895_ vdd gnd FILL
XFILL_0__8572_ vdd gnd FILL
XFILL_2__8508_ vdd gnd FILL
XFILL_2__14634_ vdd gnd FILL
XFILL_2__11846_ vdd gnd FILL
XFILL_1__13275_ vdd gnd FILL
XFILL_1__10487_ vdd gnd FILL
XFILL_0__7523_ vdd gnd FILL
XFILL_2__8439_ vdd gnd FILL
XFILL_1__12226_ vdd gnd FILL
XFILL_2__14565_ vdd gnd FILL
XFILL_0__12956_ vdd gnd FILL
XFILL_0__7454_ vdd gnd FILL
XFILL_1_BUFX2_insert9 vdd gnd FILL
XFILL_1__12157_ vdd gnd FILL
XFILL_0__11907_ vdd gnd FILL
XFILL_0__12887_ vdd gnd FILL
X_9821_ _9821_/D _9821_/CLK _9821_/Q vdd gnd DFFPOSX1
XFILL_0__7385_ vdd gnd FILL
XFILL_1__11108_ vdd gnd FILL
XFILL_0__14626_ vdd gnd FILL
XFILL_1__12088_ vdd gnd FILL
XFILL_0__11838_ vdd gnd FILL
XFILL_0__9124_ vdd gnd FILL
X_9752_ _9752_/A _9752_/B _9752_/Y vdd gnd NAND2X1
XFILL_1__11039_ vdd gnd FILL
XFILL257250x252150 vdd gnd FILL
XFILL_0__14557_ vdd gnd FILL
XFILL_0__11769_ vdd gnd FILL
XFILL_0__9055_ vdd gnd FILL
X_8703_ _8703_/A _8703_/B _8703_/Y vdd gnd NAND2X1
X_9683_ _9683_/A _9683_/B _9683_/Y vdd gnd NAND2X1
XFILL_2__12329_ vdd gnd FILL
XFILL_0__13508_ vdd gnd FILL
XFILL_0__8006_ vdd gnd FILL
XFILL_0__14488_ vdd gnd FILL
X_8634_ _8634_/A _8634_/B _8634_/C _8634_/Y vdd gnd OAI21X1
X_8565_ _8565_/A _8565_/B _8565_/Y vdd gnd NOR2X1
XFILL_1__14729_ vdd gnd FILL
X_7516_ _7516_/A _7516_/B _7516_/Y vdd gnd NAND2X1
XFILL_0__9957_ vdd gnd FILL
XFILL_1__8750_ vdd gnd FILL
X_8496_ _8496_/A _8496_/Y vdd gnd INVX1
XFILL_1__7701_ vdd gnd FILL
X_7447_ _7447_/A _7447_/B _7447_/S _7447_/Y vdd gnd MUX2X1
XFILL_0__9888_ vdd gnd FILL
XFILL_1__8681_ vdd gnd FILL
XFILL_1__7632_ vdd gnd FILL
XFILL_0__8839_ vdd gnd FILL
X_7378_ _7378_/A _7378_/Y vdd gnd INVX1
X_9117_ _9117_/A _9117_/B _9117_/Y vdd gnd NOR2X1
XFILL_1__7563_ vdd gnd FILL
XFILL_1__9302_ vdd gnd FILL
X_9048_ _9048_/A _9048_/B _9048_/C _9048_/Y vdd gnd OAI21X1
XFILL256650x150 vdd gnd FILL
XFILL_1__7494_ vdd gnd FILL
XFILL_1__9233_ vdd gnd FILL
X_11950_ _11950_/A _11950_/Y vdd gnd INVX1
XFILL_1__9164_ vdd gnd FILL
X_10901_ _10901_/A _10901_/B _10901_/Y vdd gnd NAND2X1
XFILL_1__8115_ vdd gnd FILL
X_11881_ _11881_/A _11881_/B _11881_/C _11881_/Y vdd gnd OAI21X1
XFILL_1__9095_ vdd gnd FILL
X_13620_ _13620_/A _13620_/B _13620_/C _13620_/Y vdd gnd OAI21X1
X_10832_ _10832_/A _10832_/B _10832_/C _10832_/Y vdd gnd OAI21X1
XFILL_1__8046_ vdd gnd FILL
X_13551_ _13551_/A _13551_/Y vdd gnd INVX1
X_10763_ _10763_/D _10763_/CLK _10763_/Q vdd gnd DFFPOSX1
X_12502_ _12502_/A _12502_/B _12502_/C _12502_/Y vdd gnd OAI21X1
XFILL_2__7810_ vdd gnd FILL
X_13482_ _13482_/D _13482_/CLK _13482_/Q vdd gnd DFFPOSX1
X_10694_ _10694_/D _10694_/CLK _10694_/Q vdd gnd DFFPOSX1
XFILL_1__9997_ vdd gnd FILL
X_12433_ _12433_/A _12433_/B _12433_/Y vdd gnd NAND2X1
XFILL_1__8948_ vdd gnd FILL
XFILL_2__7741_ vdd gnd FILL
X_12364_ _12364_/A _12364_/B _12364_/C _12364_/Y vdd gnd AOI21X1
XFILL_2__7672_ vdd gnd FILL
X_14103_ _14103_/A _14103_/B _14103_/C _14103_/Y vdd gnd OAI21X1
X_11315_ _11315_/A _11315_/B _11315_/C _11315_/Y vdd gnd OAI21X1
XFILL_1__10410_ vdd gnd FILL
X_12295_ _12295_/A _12295_/B _12295_/Y vdd gnd NAND2X1
XFILL_1__11390_ vdd gnd FILL
X_14034_ _14034_/A _14034_/B _14034_/Y vdd gnd NOR2X1
X_11246_ _11246_/A _11246_/B _11246_/C _11246_/D _11246_/Y vdd gnd AOI22X1
XFILL_2__11700_ vdd gnd FILL
XFILL_1__10341_ vdd gnd FILL
X_11177_ _11177_/A _11177_/B _11177_/Y vdd gnd NAND2X1
XFILL_1__13060_ vdd gnd FILL
XFILL_1__10272_ vdd gnd FILL
XFILL_0__12810_ vdd gnd FILL
XFILL_0__13790_ vdd gnd FILL
X_10128_ _10128_/A _10128_/B _10128_/Y vdd gnd OR2X2
XFILL_1__12011_ vdd gnd FILL
XFILL_2__8224_ vdd gnd FILL
XFILL_0__12741_ vdd gnd FILL
X_10059_ _10059_/A _10059_/B _10059_/C _10059_/Y vdd gnd NAND3X1
XFILL_2__13301_ vdd gnd FILL
XFILL_2__10513_ vdd gnd FILL
XFILL_2__8155_ vdd gnd FILL
XFILL_0__12672_ vdd gnd FILL
XFILL_0__7170_ vdd gnd FILL
X_14867_ _14867_/A _14867_/B _14867_/C _14867_/Y vdd gnd OAI21X1
XFILL_2__10444_ vdd gnd FILL
XFILL_0__14411_ vdd gnd FILL
XFILL_2__8086_ vdd gnd FILL
XFILL_1__13962_ vdd gnd FILL
X_13818_ _13818_/A _13818_/B _13818_/Y vdd gnd AND2X2
X_14798_ _14798_/A _14798_/B _14798_/Y vdd gnd NAND2X1
XFILL_1__12913_ vdd gnd FILL
XFILL_2__10375_ vdd gnd FILL
XFILL_0__14342_ vdd gnd FILL
XFILL_0__11554_ vdd gnd FILL
XFILL_1__13893_ vdd gnd FILL
X_13749_ _13749_/A _13749_/Y vdd gnd INVX1
XFILL_0__10505_ vdd gnd FILL
XFILL_0__14273_ vdd gnd FILL
XFILL_1__12844_ vdd gnd FILL
XFILL_0__11485_ vdd gnd FILL
XFILL_0__13224_ vdd gnd FILL
XFILL_2__8988_ vdd gnd FILL
XFILL_0__10436_ vdd gnd FILL
XFILL_1__12775_ vdd gnd FILL
X_8350_ _8350_/A _8350_/B _8350_/Y vdd gnd NAND2X1
XFILL_0__13155_ vdd gnd FILL
XFILL_1__11726_ vdd gnd FILL
XFILL_0__10367_ vdd gnd FILL
X_7301_ _7301_/A _7301_/B _7301_/C _7301_/Y vdd gnd NAND3X1
XFILL_0__9742_ vdd gnd FILL
X_8281_ _8281_/A _8281_/B _8281_/C _8281_/Y vdd gnd OAI21X1
XFILL_0__12106_ vdd gnd FILL
XFILL_1__14445_ vdd gnd FILL
XFILL_0__13086_ vdd gnd FILL
X_7232_ _7232_/A _7232_/Y vdd gnd INVX2
XFILL_0__10298_ vdd gnd FILL
XFILL_0__9673_ vdd gnd FILL
XFILL_1__10608_ vdd gnd FILL
XFILL_0__12037_ vdd gnd FILL
XFILL_1__14376_ vdd gnd FILL
XFILL_1__11588_ vdd gnd FILL
XFILL_0__8624_ vdd gnd FILL
X_7163_ _7163_/A _7163_/Y vdd gnd INVX2
XFILL_1__10539_ vdd gnd FILL
XFILL_1__13327_ vdd gnd FILL
XFILL_0__8555_ vdd gnd FILL
XFILL_2__14617_ vdd gnd FILL
X_7094_ _7094_/A _7094_/B _7094_/C _7094_/D _7094_/Y vdd gnd AOI22X1
XFILL_2__11829_ vdd gnd FILL
XFILL_1__13258_ vdd gnd FILL
XFILL_0__7506_ vdd gnd FILL
XFILL_0__13988_ vdd gnd FILL
XFILL_0__8486_ vdd gnd FILL
XFILL_1__12209_ vdd gnd FILL
XFILL_1__13189_ vdd gnd FILL
XFILL_0__12939_ vdd gnd FILL
XFILL_0__7437_ vdd gnd FILL
X_9804_ _9804_/D _9804_/CLK _9804_/Q vdd gnd DFFPOSX1
XFILL_0__7368_ vdd gnd FILL
XFILL_0__14609_ vdd gnd FILL
X_7996_ _7996_/A _7996_/Y vdd gnd INVX1
XFILL_0__9107_ vdd gnd FILL
X_9735_ _9735_/A _9735_/B _9735_/C _9735_/Y vdd gnd OAI21X1
XFILL_0__7299_ vdd gnd FILL
XFILL_0__9038_ vdd gnd FILL
XFILL_1__9920_ vdd gnd FILL
X_9666_ _9666_/A _9666_/B _9666_/C _9666_/Y vdd gnd OAI21X1
XFILL_1__9851_ vdd gnd FILL
X_8617_ _8617_/A _8617_/B _8617_/Y vdd gnd NAND2X1
X_9597_ _9597_/A _9597_/Y vdd gnd INVX1
XFILL_1__8802_ vdd gnd FILL
X_8548_ _8548_/A _8548_/Y vdd gnd INVX1
XFILL_1__8733_ vdd gnd FILL
X_8479_ _8479_/A _8479_/B _8479_/C _8479_/Y vdd gnd AOI21X1
XFILL_1__8664_ vdd gnd FILL
X_11100_ _11100_/A _11100_/B _11100_/Y vdd gnd AND2X2
XFILL_1__7615_ vdd gnd FILL
X_12080_ _12080_/A _12080_/B _12080_/C _12080_/Y vdd gnd OAI21X1
XFILL_1__8595_ vdd gnd FILL
X_11031_ _11031_/A _11031_/Y vdd gnd INVX1
XFILL_1__7546_ vdd gnd FILL
XFILL_1__7477_ vdd gnd FILL
XFILL_1__9216_ vdd gnd FILL
X_12982_ _12982_/A _12982_/B _12982_/Y vdd gnd NAND2X1
X_14721_ _14721_/A _14721_/B _14721_/Y vdd gnd NAND2X1
X_11933_ _11933_/A _11933_/B _11933_/Y vdd gnd NAND2X1
XFILL_1__9147_ vdd gnd FILL
X_14652_ _14652_/A _14652_/B _14652_/Y vdd gnd NAND2X1
X_11864_ _11864_/A _11864_/B _11864_/C _11864_/D _11864_/Y vdd gnd AOI22X1
XFILL_1__9078_ vdd gnd FILL
X_13603_ _13603_/A _13603_/B _13603_/S _13603_/Y vdd gnd MUX2X1
X_10815_ _10815_/A _10815_/B _10815_/C _10815_/Y vdd gnd OAI21X1
X_14583_ _14583_/A _14583_/B _14583_/Y vdd gnd NAND2X1
XFILL_1__8029_ vdd gnd FILL
XFILL_2__10160_ vdd gnd FILL
X_11795_ _11795_/A _11795_/Y vdd gnd INVX1
XFILL_1__10890_ vdd gnd FILL
X_13534_ _13534_/A _13534_/B _13534_/C _13534_/Y vdd gnd OAI21X1
X_10746_ _10746_/D _10746_/CLK _10746_/Q vdd gnd DFFPOSX1
XFILL_2__10091_ vdd gnd FILL
XFILL_0__11270_ vdd gnd FILL
X_13465_ _13465_/D _13465_/CLK _13465_/Q vdd gnd DFFPOSX1
X_10677_ _10677_/A _10677_/B _10677_/C _10677_/Y vdd gnd OAI21X1
XFILL_0__10221_ vdd gnd FILL
X_12416_ _12416_/A _12416_/Y vdd gnd INVX1
X_13396_ _13396_/A _13396_/B _13396_/C _13396_/Y vdd gnd OAI21X1
XFILL_1__11511_ vdd gnd FILL
XFILL_0__10152_ vdd gnd FILL
XFILL_1__12491_ vdd gnd FILL
X_12347_ _12347_/A _12347_/B _12347_/C _12347_/Y vdd gnd OAI21X1
XFILL_1__14230_ vdd gnd FILL
XFILL_1__11442_ vdd gnd FILL
XFILL_2__10993_ vdd gnd FILL
XFILL_0__10083_ vdd gnd FILL
X_12278_ _12278_/A _12278_/B _12278_/C _12278_/Y vdd gnd NAND3X1
XFILL_0__13911_ vdd gnd FILL
XFILL_2__7586_ vdd gnd FILL
XFILL_1__11373_ vdd gnd FILL
X_14017_ _14017_/A _14017_/Y vdd gnd INVX1
X_11229_ _11229_/A _11229_/B _11229_/C _11229_/Y vdd gnd OAI21X1
XFILL_1__13112_ vdd gnd FILL
XFILL_1__10324_ vdd gnd FILL
XFILL_1__14092_ vdd gnd FILL
XFILL_0__13842_ vdd gnd FILL
XFILL_0__8340_ vdd gnd FILL
XFILL_2__14402_ vdd gnd FILL
XFILL_1__13043_ vdd gnd FILL
XFILL_1__10255_ vdd gnd FILL
XFILL_0__10985_ vdd gnd FILL
XFILL_0__13773_ vdd gnd FILL
XFILL_2__8207_ vdd gnd FILL
XFILL_0__8271_ vdd gnd FILL
XFILL_1__10186_ vdd gnd FILL
XFILL_0__12724_ vdd gnd FILL
XFILL_0__7222_ vdd gnd FILL
X_14919_ _14919_/A _14919_/Y vdd gnd BUFX2
X_7850_ _7850_/A _7850_/B _7850_/C _7850_/Y vdd gnd OAI21X1
XFILL_2__8138_ vdd gnd FILL
XFILL_0__12655_ vdd gnd FILL
XFILL_0__7153_ vdd gnd FILL
XFILL_2__13215_ vdd gnd FILL
XFILL_2__10427_ vdd gnd FILL
X_7781_ _7781_/A _7781_/Y vdd gnd INVX1
XFILL_2__8069_ vdd gnd FILL
XFILL_0__11606_ vdd gnd FILL
XFILL_1__13945_ vdd gnd FILL
X_9520_ _9520_/A _9520_/B _9520_/Y vdd gnd NOR2X1
XFILL_0__7084_ vdd gnd FILL
XFILL_2__13146_ vdd gnd FILL
XFILL_2__10358_ vdd gnd FILL
XFILL_0__14325_ vdd gnd FILL
XFILL_0__11537_ vdd gnd FILL
XFILL_1__13876_ vdd gnd FILL
X_9451_ _9451_/A _9451_/Y vdd gnd INVX1
XFILL_2__13077_ vdd gnd FILL
XFILL_0__14256_ vdd gnd FILL
XFILL_1__12827_ vdd gnd FILL
XFILL_2__10289_ vdd gnd FILL
XFILL_0__11468_ vdd gnd FILL
X_8402_ _8402_/A _8402_/Y vdd gnd INVX1
X_9382_ _9382_/A _9382_/B _9382_/Y vdd gnd NAND2X1
XFILL_0__13207_ vdd gnd FILL
XFILL_0__10419_ vdd gnd FILL
XFILL_0_BUFX2_insert380 vdd gnd FILL
XFILL_1__12758_ vdd gnd FILL
XFILL_0__11399_ vdd gnd FILL
X_8333_ _8333_/A _8333_/B _8333_/C _8333_/Y vdd gnd AOI21X1
XFILL_0__13138_ vdd gnd FILL
XFILL_1__11709_ vdd gnd FILL
XFILL_0__9725_ vdd gnd FILL
XFILL_1__12689_ vdd gnd FILL
X_8264_ _8264_/A _8264_/B _8264_/Y vdd gnd NAND2X1
XFILL_1__14428_ vdd gnd FILL
XFILL_0__13069_ vdd gnd FILL
X_7215_ _7215_/A _7215_/B _7215_/C _7215_/Y vdd gnd AOI21X1
XFILL_0__9656_ vdd gnd FILL
X_8195_ _8195_/A _8195_/B _8195_/C _8195_/Y vdd gnd NAND3X1
XFILL_1__14359_ vdd gnd FILL
XFILL_1__7400_ vdd gnd FILL
XFILL_0__8607_ vdd gnd FILL
X_7146_ _7146_/A _7146_/B _7146_/C _7146_/Y vdd gnd OAI21X1
XFILL_0__9587_ vdd gnd FILL
XFILL_1__8380_ vdd gnd FILL
XFILL_1__7331_ vdd gnd FILL
XFILL_0__8538_ vdd gnd FILL
X_7077_ _7077_/A _7077_/Y vdd gnd INVX4
XFILL_1__7262_ vdd gnd FILL
XFILL_0__8469_ vdd gnd FILL
XFILL_1__9001_ vdd gnd FILL
XFILL_1__7193_ vdd gnd FILL
X_7979_ _7979_/D _7979_/CLK _7979_/Q vdd gnd DFFPOSX1
X_9718_ _9718_/A _9718_/B _9718_/C _9718_/Y vdd gnd OAI21X1
X_10600_ _10600_/A _10600_/B _10600_/C _10600_/Y vdd gnd OAI21X1
XFILL_1__9903_ vdd gnd FILL
X_11580_ _11580_/A _11580_/B _11580_/C _11580_/Y vdd gnd OAI21X1
X_9649_ _9649_/A _9649_/B _9649_/C _9649_/Y vdd gnd OAI21X1
X_10531_ _10531_/A _10531_/B _10531_/Y vdd gnd NAND2X1
X_13250_ _13250_/A _13250_/B _13250_/Y vdd gnd NOR2X1
X_10462_ _10462_/A _10462_/B _10462_/Y vdd gnd NAND2X1
X_12201_ _12201_/A _12201_/B _12201_/Y vdd gnd NAND2X1
X_13181_ _13181_/A _13181_/B _13181_/C _13181_/Y vdd gnd OAI21X1
XFILL_1__8716_ vdd gnd FILL
X_10393_ _10393_/A _10393_/B _10393_/C _10393_/Y vdd gnd AOI21X1
XFILL_1__9696_ vdd gnd FILL
X_12132_ _12132_/A _12132_/B _12132_/S _12132_/Y vdd gnd MUX2X1
XFILL_1__8647_ vdd gnd FILL
X_12063_ _12063_/A _12063_/B _12063_/Y vdd gnd NAND2X1
XFILL_1__8578_ vdd gnd FILL
X_11014_ _11014_/A _11014_/B _11014_/C _11014_/Y vdd gnd AOI21X1
XFILL_2__9110_ vdd gnd FILL
XFILL_1__7529_ vdd gnd FILL
XFILL_1__10040_ vdd gnd FILL
XFILL_0__10770_ vdd gnd FILL
X_12965_ _12965_/A _12965_/Y vdd gnd INVX1
X_14704_ _14704_/A _14704_/B _14704_/Y vdd gnd NAND2X1
X_11916_ _11916_/A _11916_/B _11916_/C _11916_/Y vdd gnd OAI21X1
X_12896_ _12896_/A _12896_/B _12896_/Y vdd gnd NOR2X1
XFILL_0__12440_ vdd gnd FILL
X_14635_ _14635_/A _14635_/B _14635_/C _14635_/Y vdd gnd NAND3X1
XFILL_1__11991_ vdd gnd FILL
X_11847_ _11847_/A _11847_/B _11847_/C _11847_/Y vdd gnd AOI21X1
XFILL_2__13000_ vdd gnd FILL
XFILL_2__9943_ vdd gnd FILL
XFILL_1__13730_ vdd gnd FILL
XFILL_1__10942_ vdd gnd FILL
XFILL_0__12371_ vdd gnd FILL
X_14566_ _14566_/A _14566_/B _14566_/Y vdd gnd NAND2X1
X_11778_ _11778_/A _11778_/B _11778_/Y vdd gnd NAND2X1
XFILL_0__14110_ vdd gnd FILL
XFILL_2__9874_ vdd gnd FILL
XFILL_0__11322_ vdd gnd FILL
XFILL_1__13661_ vdd gnd FILL
X_13517_ _13517_/A _13517_/B _13517_/C _13517_/D _13517_/Y vdd gnd AOI22X1
XFILL_1__10873_ vdd gnd FILL
X_10729_ _10729_/D _10729_/CLK _10729_/Q vdd gnd DFFPOSX1
XFILL_2__8825_ vdd gnd FILL
X_14497_ _14497_/A _14497_/B _14497_/C _14497_/Y vdd gnd OAI21X1
XFILL_0__14041_ vdd gnd FILL
XFILL_0__11253_ vdd gnd FILL
XFILL256050x21750 vdd gnd FILL
XFILL_1__13592_ vdd gnd FILL
X_13448_ _13448_/D _13448_/CLK _13448_/Q vdd gnd DFFPOSX1
XFILL_0__7840_ vdd gnd FILL
XFILL_0__10204_ vdd gnd FILL
XFILL_2__8756_ vdd gnd FILL
XFILL_0__11184_ vdd gnd FILL
XFILL_0__7771_ vdd gnd FILL
X_13379_ _13379_/A _13379_/B _13379_/C _13379_/Y vdd gnd OAI21X1
XFILL_0__10135_ vdd gnd FILL
XFILL_0__9510_ vdd gnd FILL
XFILL_1__12474_ vdd gnd FILL
XFILL256050x223350 vdd gnd FILL
XFILL_1__11425_ vdd gnd FILL
XFILL_0__10066_ vdd gnd FILL
XFILL_0__9441_ vdd gnd FILL
XFILL_1_BUFX2_insert14 vdd gnd FILL
XFILL_1__14144_ vdd gnd FILL
XFILL_1__11356_ vdd gnd FILL
XFILL_1_BUFX2_insert25 vdd gnd FILL
XFILL_0__9372_ vdd gnd FILL
XFILL_1__10307_ vdd gnd FILL
XFILL_1__11287_ vdd gnd FILL
XFILL_0__13825_ vdd gnd FILL
XFILL_1__14075_ vdd gnd FILL
XFILL_0__8323_ vdd gnd FILL
X_8951_ _8951_/A _8951_/B _8951_/C _8951_/D _8951_/Y vdd gnd AOI22X1
XFILL_1__10238_ vdd gnd FILL
XFILL_1__13026_ vdd gnd FILL
XFILL_0__13756_ vdd gnd FILL
XFILL_0__10968_ vdd gnd FILL
X_7902_ _7902_/A _7902_/B _7902_/Y vdd gnd NAND2X1
XFILL_0__8254_ vdd gnd FILL
XFILL_2__14316_ vdd gnd FILL
X_8882_ _8882_/D _8882_/CLK _8882_/Q vdd gnd DFFPOSX1
XFILL_1__10169_ vdd gnd FILL
XFILL_0__12707_ vdd gnd FILL
XFILL_0__7205_ vdd gnd FILL
XFILL_0__10899_ vdd gnd FILL
XFILL_0__13687_ vdd gnd FILL
X_7833_ _7833_/A _7833_/B _7833_/Y vdd gnd NAND2X1
XFILL_0__8185_ vdd gnd FILL
XFILL_2__14247_ vdd gnd FILL
XFILL_0__12638_ vdd gnd FILL
XFILL_0__7136_ vdd gnd FILL
XFILL_1_CLKBUF1_insert37 vdd gnd FILL
X_7764_ _7764_/A _7764_/B _7764_/Y vdd gnd NAND2X1
XFILL_1_CLKBUF1_insert48 vdd gnd FILL
XFILL_1__13928_ vdd gnd FILL
XFILL_1_CLKBUF1_insert59 vdd gnd FILL
X_9503_ _9503_/A _9503_/Y vdd gnd INVX1
XFILL_2__13129_ vdd gnd FILL
X_7695_ _7695_/A _7695_/B _7695_/Y vdd gnd NOR2X1
XFILL_0__14308_ vdd gnd FILL
XFILL_1__13859_ vdd gnd FILL
X_9434_ _9434_/A _9434_/B _9434_/Y vdd gnd NOR2X1
XFILL_1__7880_ vdd gnd FILL
XFILL_0__14239_ vdd gnd FILL
X_9365_ _9365_/A _9365_/B _9365_/Y vdd gnd OR2X2
XFILL_1__9550_ vdd gnd FILL
X_8316_ _8316_/A _8316_/B _8316_/C _8316_/Y vdd gnd OAI21X1
X_9296_ _9296_/A _9296_/B _9296_/Y vdd gnd NAND2X1
XFILL_1__8501_ vdd gnd FILL
XFILL_0__9708_ vdd gnd FILL
XFILL_1__9481_ vdd gnd FILL
X_8247_ _8247_/A _8247_/B _8247_/Y vdd gnd AND2X2
XFILL_0__9639_ vdd gnd FILL
XFILL_1__8432_ vdd gnd FILL
X_8178_ _8178_/A _8178_/B _8178_/C _8178_/Y vdd gnd AOI21X1
X_7129_ _7129_/A _7129_/B _7129_/C _7129_/Y vdd gnd OAI21X1
XFILL_1__8363_ vdd gnd FILL
XFILL_1__7314_ vdd gnd FILL
XFILL_1__8294_ vdd gnd FILL
XFILL_1__7245_ vdd gnd FILL
X_12750_ _12750_/A _12750_/B _12750_/C _12750_/D _12750_/Y vdd gnd OAI22X1
XFILL_1__7176_ vdd gnd FILL
X_11701_ _11701_/A _11701_/B _11701_/Y vdd gnd AND2X2
X_12681_ _12681_/A _12681_/Y vdd gnd INVX1
X_14420_ _14420_/A _14420_/B _14420_/Y vdd gnd NAND2X1
X_11632_ _11632_/D _11632_/CLK _11632_/Q vdd gnd DFFPOSX1
X_14351_ _14351_/A _14351_/Y vdd gnd INVX1
X_11563_ _11563_/A _11563_/B _11563_/C _11563_/Y vdd gnd OAI21X1
X_13302_ _13302_/A _13302_/Y vdd gnd INVX1
X_10514_ _10514_/A _10514_/B _10514_/Y vdd gnd NAND2X1
X_14282_ _14282_/A _14282_/B _14282_/C _14282_/Y vdd gnd OAI21X1
XFILL_2__8610_ vdd gnd FILL
X_11494_ _11494_/A _11494_/Y vdd gnd INVX1
X_13233_ _13233_/A _13233_/B _13233_/Y vdd gnd OR2X2
X_10445_ _10445_/A _10445_/B _10445_/Y vdd gnd NOR2X1
XFILL_2__8541_ vdd gnd FILL
XFILL_1__9748_ vdd gnd FILL
X_13164_ _13164_/A _13164_/B _13164_/C _13164_/Y vdd gnd NAND3X1
X_10376_ _10376_/A _10376_/B _10376_/C _10376_/Y vdd gnd OAI21X1
XFILL_1__9679_ vdd gnd FILL
XFILL_2__8472_ vdd gnd FILL
X_12115_ _12115_/A _12115_/B _12115_/C _12115_/Y vdd gnd AOI21X1
X_13095_ _13095_/A _13095_/Y vdd gnd INVX1
XFILL_1__11210_ vdd gnd FILL
XFILL_1__12190_ vdd gnd FILL
XFILL_0__11940_ vdd gnd FILL
X_12046_ _12046_/A _12046_/B _12046_/Y vdd gnd NAND2X1
XFILL_1__11141_ vdd gnd FILL
XFILL_0__11871_ vdd gnd FILL
XFILL_1__11072_ vdd gnd FILL
XFILL_0__13610_ vdd gnd FILL
XFILL_0__10822_ vdd gnd FILL
XFILL_0__14590_ vdd gnd FILL
XFILL_2__9024_ vdd gnd FILL
XFILL_1__10023_ vdd gnd FILL
X_13997_ _13997_/A _13997_/B _13997_/C _13997_/Y vdd gnd NAND3X1
XFILL_2_BUFX2_insert272 vdd gnd FILL
XFILL_0__13541_ vdd gnd FILL
X_12948_ _12948_/A _12948_/B _12948_/C _12948_/Y vdd gnd AOI21X1
XFILL_2__14101_ vdd gnd FILL
XFILL_2_BUFX2_insert294 vdd gnd FILL
XFILL_2__11313_ vdd gnd FILL
XFILL_1__14831_ vdd gnd FILL
XFILL_0__10684_ vdd gnd FILL
XFILL_2__14032_ vdd gnd FILL
X_12879_ _12879_/A _12879_/B _12879_/Y vdd gnd NAND2X1
XFILL_2__11244_ vdd gnd FILL
XFILL_1__14762_ vdd gnd FILL
XFILL_0__12423_ vdd gnd FILL
XFILL_1__11974_ vdd gnd FILL
X_14618_ _14618_/A _14618_/B _14618_/Y vdd gnd AND2X2
XFILL_0__9990_ vdd gnd FILL
XFILL_2__9926_ vdd gnd FILL
XFILL_1__13713_ vdd gnd FILL
XFILL_0__12354_ vdd gnd FILL
XFILL_1__10925_ vdd gnd FILL
XFILL_2__11175_ vdd gnd FILL
XFILL_1__14693_ vdd gnd FILL
XFILL_0__8941_ vdd gnd FILL
X_14549_ _14549_/D _14549_/CLK _14549_/Q vdd gnd DFFPOSX1
X_7480_ _7480_/A _7480_/B _7480_/Y vdd gnd AND2X2
XBUFX2_insert260 BUFX2_insert260/A BUFX2_insert260/Y vdd gnd BUFX2
XFILL_0__11305_ vdd gnd FILL
XFILL_2__9857_ vdd gnd FILL
XFILL_1__13644_ vdd gnd FILL
XBUFX2_insert271 BUFX2_insert271/A BUFX2_insert271/Y vdd gnd BUFX2
XFILL_0__12285_ vdd gnd FILL
XFILL_1__10856_ vdd gnd FILL
XBUFX2_insert282 BUFX2_insert282/A BUFX2_insert282/Y vdd gnd BUFX2
XBUFX2_insert293 BUFX2_insert293/A BUFX2_insert293/Y vdd gnd BUFX2
XFILL_2__8808_ vdd gnd FILL
XFILL_0__14024_ vdd gnd FILL
XFILL_0__11236_ vdd gnd FILL
XFILL_1__13575_ vdd gnd FILL
XFILL_0__7823_ vdd gnd FILL
XFILL_1__10787_ vdd gnd FILL
X_9150_ _9150_/A _9150_/B _9150_/C _9150_/Y vdd gnd AOI21X1
XFILL_2__14865_ vdd gnd FILL
XFILL_2__8739_ vdd gnd FILL
XFILL_1__12526_ vdd gnd FILL
XFILL_0__11167_ vdd gnd FILL
X_8101_ _8101_/A _8101_/B _8101_/C _8101_/Y vdd gnd OAI21X1
XFILL_0__7754_ vdd gnd FILL
X_9081_ _9081_/A _9081_/B _9081_/C _9081_/Y vdd gnd OAI21X1
XFILL_0__10118_ vdd gnd FILL
XFILL_2__14796_ vdd gnd FILL
XFILL_1__12457_ vdd gnd FILL
XFILL_0__11098_ vdd gnd FILL
X_8032_ _8032_/A _8032_/Y vdd gnd INVX1
XFILL_0__7685_ vdd gnd FILL
XFILL_1__11408_ vdd gnd FILL
XFILL_0__10049_ vdd gnd FILL
XFILL_0__9424_ vdd gnd FILL
XFILL_1__12388_ vdd gnd FILL
XFILL_1__14127_ vdd gnd FILL
XFILL_1__11339_ vdd gnd FILL
XFILL_0__14857_ vdd gnd FILL
XFILL_0__9355_ vdd gnd FILL
X_9983_ _9983_/A _9983_/B _9983_/S _9983_/Y vdd gnd MUX2X1
XFILL_2__12629_ vdd gnd FILL
XFILL_1__14058_ vdd gnd FILL
XFILL_0__13808_ vdd gnd FILL
XFILL_0__8306_ vdd gnd FILL
XFILL_0__14788_ vdd gnd FILL
XFILL_0__9286_ vdd gnd FILL
X_8934_ _8934_/A _8934_/B _8934_/C _8934_/Y vdd gnd OAI21X1
XFILL_1__13009_ vdd gnd FILL
XFILL_0__13739_ vdd gnd FILL
XFILL_0__8237_ vdd gnd FILL
X_8865_ _8865_/D _8865_/CLK _8865_/Q vdd gnd DFFPOSX1
X_7816_ _7816_/A _7816_/B _7816_/C _7816_/D _7816_/Y vdd gnd OAI22X1
XFILL_0__8168_ vdd gnd FILL
X_8796_ _8796_/A _8796_/B _8796_/C _8796_/Y vdd gnd OAI21X1
XFILL_0__7119_ vdd gnd FILL
XFILL_1__8981_ vdd gnd FILL
X_7747_ _7747_/A _7747_/B _7747_/C _7747_/Y vdd gnd OAI21X1
XFILL_0__8099_ vdd gnd FILL
X_7678_ _7678_/A _7678_/B _7678_/Y vdd gnd NAND2X1
X_9417_ _9417_/A _9417_/B _9417_/Y vdd gnd AND2X2
XFILL_1__7863_ vdd gnd FILL
XFILL_1__9602_ vdd gnd FILL
X_9348_ _9348_/A _9348_/B _9348_/C _9348_/Y vdd gnd NAND3X1
XFILL_1__7794_ vdd gnd FILL
X_10230_ _10230_/A _10230_/B _10230_/Y vdd gnd NOR2X1
XFILL_1__9533_ vdd gnd FILL
X_9279_ _9279_/A _9279_/B _9279_/C _9279_/Y vdd gnd OAI21X1
X_10161_ _10161_/A _10161_/B _10161_/Y vdd gnd AND2X2
XFILL_1__9464_ vdd gnd FILL
XFILL_1__8415_ vdd gnd FILL
X_10092_ _10092_/A _10092_/B _10092_/C _10092_/D _10092_/Y vdd gnd AOI22X1
XFILL_1__9395_ vdd gnd FILL
X_13920_ _13920_/A _13920_/B _13920_/C _13920_/Y vdd gnd OAI21X1
XFILL_1__8346_ vdd gnd FILL
X_13851_ _13851_/A _13851_/B _13851_/C _13851_/Y vdd gnd OAI21X1
XFILL_1__8277_ vdd gnd FILL
X_12802_ _12802_/A _12802_/B _12802_/C _12802_/Y vdd gnd OAI21X1
XFILL_1__7228_ vdd gnd FILL
X_13782_ _13782_/A _13782_/B _13782_/C _13782_/Y vdd gnd AOI21X1
X_10994_ _10994_/A _10994_/B _10994_/C _10994_/Y vdd gnd OAI21X1
XFILL_1_BUFX2_insert202 vdd gnd FILL
XFILL_1_BUFX2_insert213 vdd gnd FILL
XFILL_1_BUFX2_insert224 vdd gnd FILL
XFILL_1_BUFX2_insert235 vdd gnd FILL
X_12733_ _12733_/A _12733_/B _12733_/C _12733_/Y vdd gnd AOI21X1
XFILL_1__7159_ vdd gnd FILL
XFILL_1_BUFX2_insert246 vdd gnd FILL
XFILL_1_BUFX2_insert257 vdd gnd FILL
XFILL_1_BUFX2_insert268 vdd gnd FILL
XFILL_1_BUFX2_insert279 vdd gnd FILL
X_12664_ _12664_/A _12664_/B _12664_/C _12664_/Y vdd gnd OAI21X1
XCLKBUF1_insert39 CLKBUF1_insert39/A CLKBUF1_insert39/Y vdd gnd CLKBUF1
X_14403_ _14403_/A _14403_/B _14403_/Y vdd gnd NAND2X1
X_11615_ _11615_/D _11615_/CLK _11615_/Q vdd gnd DFFPOSX1
X_12595_ _12595_/D _12595_/CLK _12595_/Q vdd gnd DFFPOSX1
X_14334_ _14334_/A _14334_/B _14334_/Y vdd gnd NAND2X1
X_11546_ _11546_/A _11546_/B _11546_/C _11546_/Y vdd gnd OAI21X1
XFILL_1__10641_ vdd gnd FILL
XFILL_0__12070_ vdd gnd FILL
X_14265_ _14265_/A _14265_/B _14265_/Y vdd gnd OR2X2
X_11477_ _11477_/A _11477_/Y vdd gnd INVX1
XFILL_0__11021_ vdd gnd FILL
XFILL_2__11931_ vdd gnd FILL
XFILL_1__13360_ vdd gnd FILL
X_13216_ _13216_/A _13216_/B _13216_/Y vdd gnd NOR2X1
XFILL_1__10572_ vdd gnd FILL
X_10428_ _10428_/A _10428_/B _10428_/C _10428_/Y vdd gnd AOI21X1
XFILL_2__8524_ vdd gnd FILL
X_14196_ _14196_/D _14196_/CLK _14196_/Q vdd gnd DFFPOSX1
XFILL_1__12311_ vdd gnd FILL
XFILL_2__11862_ vdd gnd FILL
XFILL_1__13291_ vdd gnd FILL
X_13147_ _13147_/A _13147_/B _13147_/C _13147_/Y vdd gnd NAND3X1
XFILL_2__13601_ vdd gnd FILL
X_10359_ _10359_/A _10359_/B _10359_/C _10359_/Y vdd gnd OAI21X1
XFILL_2__8455_ vdd gnd FILL
XFILL_2__14581_ vdd gnd FILL
XFILL_1__12242_ vdd gnd FILL
XFILL_2__11793_ vdd gnd FILL
XFILL_0__12972_ vdd gnd FILL
X_13078_ _13078_/A _13078_/B _13078_/C _13078_/Y vdd gnd OAI21X1
XFILL_0__7470_ vdd gnd FILL
XFILL_2__13532_ vdd gnd FILL
XFILL_0__14711_ vdd gnd FILL
XFILL_2__8386_ vdd gnd FILL
XFILL_0__11923_ vdd gnd FILL
XFILL_1__12173_ vdd gnd FILL
X_12029_ _12029_/A _12029_/B _12029_/C _12029_/Y vdd gnd AOI21X1
XFILL_1__11124_ vdd gnd FILL
XFILL_0__14642_ vdd gnd FILL
XFILL_2__10675_ vdd gnd FILL
XFILL_0__9140_ vdd gnd FILL
XFILL_0__11854_ vdd gnd FILL
XFILL_1__11055_ vdd gnd FILL
XFILL_2__13394_ vdd gnd FILL
XFILL_0__10805_ vdd gnd FILL
XFILL_0__14573_ vdd gnd FILL
XFILL_0__9071_ vdd gnd FILL
XFILL_2__9007_ vdd gnd FILL
XFILL_0__11785_ vdd gnd FILL
XFILL_1__10006_ vdd gnd FILL
XFILL_0__13524_ vdd gnd FILL
XFILL_0__8022_ vdd gnd FILL
X_8650_ _8650_/A _8650_/B _8650_/C _8650_/Y vdd gnd OAI21X1
XFILL_1__14814_ vdd gnd FILL
XFILL_0__10667_ vdd gnd FILL
X_7601_ _7601_/A _7601_/B _7601_/Y vdd gnd NAND2X1
X_8581_ _8581_/A _8581_/B _8581_/Y vdd gnd NOR2X1
XFILL_2__11227_ vdd gnd FILL
XFILL_1__14745_ vdd gnd FILL
XFILL_0__12406_ vdd gnd FILL
XFILL_1__11957_ vdd gnd FILL
XFILL_0__10598_ vdd gnd FILL
XFILL_0__13386_ vdd gnd FILL
X_7532_ _7532_/A _7532_/B _7532_/Y vdd gnd NAND2X1
XFILL_2__9909_ vdd gnd FILL
XFILL_0__9973_ vdd gnd FILL
XFILL_1__10908_ vdd gnd FILL
XFILL_2__11158_ vdd gnd FILL
XFILL_1__14676_ vdd gnd FILL
XFILL_0__12337_ vdd gnd FILL
XFILL_1__11888_ vdd gnd FILL
XFILL_0__8924_ vdd gnd FILL
X_7463_ _7463_/A _7463_/B _7463_/S _7463_/Y vdd gnd MUX2X1
XFILL_1__13627_ vdd gnd FILL
XFILL_0__12268_ vdd gnd FILL
XFILL_1__10839_ vdd gnd FILL
XFILL_2__11089_ vdd gnd FILL
X_9202_ _9202_/A _9202_/B _9202_/C _9202_/Y vdd gnd AOI21X1
XFILL_0__14007_ vdd gnd FILL
X_7394_ _7394_/A _7394_/Y vdd gnd INVX1
XFILL_0__11219_ vdd gnd FILL
XFILL_1__13558_ vdd gnd FILL
XFILL_0__7806_ vdd gnd FILL
XFILL_0__12199_ vdd gnd FILL
X_9133_ _9133_/A _9133_/B _9133_/Y vdd gnd NAND2X1
XFILL_0__8786_ vdd gnd FILL
XFILL_1__12509_ vdd gnd FILL
XFILL_2__14848_ vdd gnd FILL
XFILL_0__7737_ vdd gnd FILL
X_9064_ _9064_/A _9064_/B _9064_/Y vdd gnd NAND2X1
XFILL_2__14779_ vdd gnd FILL
X_8015_ _8015_/A _8015_/B _8015_/Y vdd gnd NAND2X1
XFILL_0__7668_ vdd gnd FILL
XFILL_0__14909_ vdd gnd FILL
XFILL_0__9407_ vdd gnd FILL
XFILL_1__8200_ vdd gnd FILL
XFILL_1__9180_ vdd gnd FILL
XFILL_0__7599_ vdd gnd FILL
XFILL_0__9338_ vdd gnd FILL
XFILL_1__8131_ vdd gnd FILL
X_9966_ _9966_/A _9966_/B _9966_/S _9966_/Y vdd gnd MUX2X1
XFILL_0__9269_ vdd gnd FILL
X_8917_ _8917_/D _8917_/CLK _8917_/Q vdd gnd DFFPOSX1
XFILL_1__8062_ vdd gnd FILL
X_9897_ _9897_/A _9897_/B _9897_/C _9897_/Y vdd gnd OAI21X1
X_8848_ _8848_/D _8848_/CLK _8848_/Q vdd gnd DFFPOSX1
XFILL_0_BUFX2_insert209 vdd gnd FILL
X_8779_ _8779_/A _8779_/B _8779_/C _8779_/Y vdd gnd OAI21X1
XFILL_1__8964_ vdd gnd FILL
X_11400_ _11400_/A _11400_/B _11400_/Y vdd gnd NOR2X1
X_12380_ _12380_/A _12380_/B _12380_/Y vdd gnd NAND2X1
XFILL_1__7915_ vdd gnd FILL
XFILL256950x176550 vdd gnd FILL
X_11331_ _11331_/A _11331_/Y vdd gnd INVX1
XFILL_1__7846_ vdd gnd FILL
X_14050_ _14050_/A _14050_/B _14050_/Y vdd gnd OR2X2
X_11262_ _11262_/A _11262_/B _11262_/C _11262_/Y vdd gnd NAND3X1
XFILL_1__7777_ vdd gnd FILL
X_13001_ _13001_/A _13001_/B _13001_/Y vdd gnd NAND2X1
X_10213_ _10213_/A _10213_/B _10213_/C _10213_/D _10213_/Y vdd gnd AOI22X1
XFILL_1__9516_ vdd gnd FILL
X_11193_ _11193_/A _11193_/B _11193_/C _11193_/Y vdd gnd NAND3X1
X_10144_ _10144_/A _10144_/B _10144_/Y vdd gnd AND2X2
XFILL_1__9447_ vdd gnd FILL
X_10075_ _10075_/A _10075_/B _10075_/Y vdd gnd NAND2X1
XFILL_1__9378_ vdd gnd FILL
X_13903_ _13903_/A _13903_/B _13903_/C _13903_/Y vdd gnd OAI21X1
XFILL_2__7122_ vdd gnd FILL
XFILL_1__8329_ vdd gnd FILL
X_14883_ _14883_/D _14883_/CLK _14883_/Q vdd gnd DFFPOSX1
XFILL257250x75750 vdd gnd FILL
X_13834_ _13834_/A _13834_/B _13834_/Y vdd gnd NAND2X1
XFILL_0__11570_ vdd gnd FILL
X_13765_ _13765_/A _13765_/Y vdd gnd INVX1
X_10977_ _10977_/A _10977_/B _10977_/C _10977_/Y vdd gnd NAND3X1
XFILL_0__10521_ vdd gnd FILL
XFILL_1__12860_ vdd gnd FILL
X_12716_ _12716_/A _12716_/Y vdd gnd INVX1
X_13696_ _13696_/A _13696_/B _13696_/Y vdd gnd NAND2X1
XFILL_1__11811_ vdd gnd FILL
XFILL_0__10452_ vdd gnd FILL
XFILL_0__13240_ vdd gnd FILL
XFILL_1__12791_ vdd gnd FILL
X_12647_ _12647_/A _12647_/B _12647_/C _12647_/Y vdd gnd OAI21X1
XFILL_2__11012_ vdd gnd FILL
XFILL_0__13171_ vdd gnd FILL
XFILL_1__11742_ vdd gnd FILL
XFILL_0__10383_ vdd gnd FILL
X_12578_ _12578_/D _12578_/CLK _12578_/Q vdd gnd DFFPOSX1
XFILL_0__12122_ vdd gnd FILL
XFILL_1__14461_ vdd gnd FILL
X_14317_ _14317_/A _14317_/B _14317_/C _14317_/Y vdd gnd OAI21X1
X_11529_ _11529_/A _11529_/B _11529_/Y vdd gnd NAND2X1
XFILL_1__13412_ vdd gnd FILL
XFILL_1__10624_ vdd gnd FILL
XFILL_0__12053_ vdd gnd FILL
XFILL_1__14392_ vdd gnd FILL
X_14248_ _14248_/A _14248_/B _14248_/C _14248_/Y vdd gnd OAI21X1
XFILL_0__8640_ vdd gnd FILL
XFILL_0__11004_ vdd gnd FILL
XFILL_1__13343_ vdd gnd FILL
XFILL_1__10555_ vdd gnd FILL
XFILL_0__8571_ vdd gnd FILL
X_14179_ _14179_/D _14179_/CLK _14179_/Q vdd gnd DFFPOSX1
XFILL_1__13274_ vdd gnd FILL
XFILL_0__7522_ vdd gnd FILL
XFILL_1__10486_ vdd gnd FILL
XFILL_1__12225_ vdd gnd FILL
XFILL_2__11776_ vdd gnd FILL
XFILL_0__12955_ vdd gnd FILL
XFILL_0__7453_ vdd gnd FILL
XFILL_2__13515_ vdd gnd FILL
XFILL_2__8369_ vdd gnd FILL
XFILL_0__11906_ vdd gnd FILL
XFILL_1__12156_ vdd gnd FILL
X_9820_ _9820_/D _9820_/CLK _9820_/Q vdd gnd DFFPOSX1
XFILL_0__12886_ vdd gnd FILL
XFILL_0__7384_ vdd gnd FILL
XFILL_1__11107_ vdd gnd FILL
XFILL256950x241350 vdd gnd FILL
XFILL_0__14625_ vdd gnd FILL
XFILL_2__10658_ vdd gnd FILL
XFILL_0__9123_ vdd gnd FILL
XFILL_0__11837_ vdd gnd FILL
XFILL_1__12087_ vdd gnd FILL
XFILL257550x226950 vdd gnd FILL
X_9751_ _9751_/A _9751_/B _9751_/C _9751_/Y vdd gnd OAI21X1
XFILL_1__11038_ vdd gnd FILL
XFILL_2__13377_ vdd gnd FILL
XFILL_0__14556_ vdd gnd FILL
XFILL_2__10589_ vdd gnd FILL
XFILL_0__9054_ vdd gnd FILL
X_8702_ _8702_/A _8702_/B _8702_/Y vdd gnd NAND2X1
XFILL_0__11768_ vdd gnd FILL
X_9682_ _9682_/A _9682_/B _9682_/Y vdd gnd NOR2X1
XFILL_0__13507_ vdd gnd FILL
XFILL_0__8005_ vdd gnd FILL
XFILL_0__14487_ vdd gnd FILL
X_8633_ _8633_/A _8633_/B _8633_/C _8633_/Y vdd gnd OAI21X1
XFILL_0__11699_ vdd gnd FILL
XFILL_1__12989_ vdd gnd FILL
X_8564_ _8564_/A _8564_/B _8564_/Y vdd gnd NOR2X1
XFILL_1__14728_ vdd gnd FILL
XFILL_0__13369_ vdd gnd FILL
X_7515_ _7515_/A _7515_/B _7515_/Y vdd gnd NAND2X1
XFILL_0__9956_ vdd gnd FILL
X_8495_ _8495_/A _8495_/B _8495_/C _8495_/Y vdd gnd OAI21X1
XFILL_1__14659_ vdd gnd FILL
XFILL_1__7700_ vdd gnd FILL
X_7446_ _7446_/A _7446_/B _7446_/C _7446_/Y vdd gnd OAI21X1
XFILL_1__8680_ vdd gnd FILL
XFILL_0__9887_ vdd gnd FILL
XFILL_1__7631_ vdd gnd FILL
XFILL_0__8838_ vdd gnd FILL
X_7377_ _7377_/A _7377_/B _7377_/C _7377_/Y vdd gnd AOI21X1
XFILL256950x108150 vdd gnd FILL
X_9116_ _9116_/A _9116_/B _9116_/Y vdd gnd OR2X2
XFILL_1__7562_ vdd gnd FILL
XFILL_0__8769_ vdd gnd FILL
XFILL_1__9301_ vdd gnd FILL
X_9047_ _9047_/A _9047_/B _9047_/Y vdd gnd AND2X2
XFILL_1__7493_ vdd gnd FILL
XFILL_1__9232_ vdd gnd FILL
XFILL_1__9163_ vdd gnd FILL
XFILL257550x136950 vdd gnd FILL
X_10900_ _10900_/A _10900_/Y vdd gnd INVX1
XFILL_1__8114_ vdd gnd FILL
X_11880_ _11880_/A _11880_/B _11880_/Y vdd gnd NAND2X1
XFILL_1__9094_ vdd gnd FILL
X_9949_ _9949_/A _9949_/B _9949_/C _9949_/Y vdd gnd OAI21X1
X_10831_ _10831_/A _10831_/B _10831_/Y vdd gnd NAND2X1
XFILL_1__8045_ vdd gnd FILL
X_13550_ _13550_/A _13550_/B _13550_/C _13550_/Y vdd gnd OAI21X1
X_10762_ _10762_/D _10762_/CLK _10762_/Q vdd gnd DFFPOSX1
X_12501_ _12501_/A _12501_/B _12501_/C _12501_/Y vdd gnd OAI21X1
X_13481_ _13481_/D _13481_/CLK _13481_/Q vdd gnd DFFPOSX1
X_10693_ _10693_/D _10693_/CLK _10693_/Q vdd gnd DFFPOSX1
XFILL_1__9996_ vdd gnd FILL
X_12432_ _12432_/A _12432_/B _12432_/Y vdd gnd NAND2X1
XFILL_1__8947_ vdd gnd FILL
XFILL257250x50550 vdd gnd FILL
X_12363_ _12363_/A _12363_/B _12363_/Y vdd gnd NAND2X1
X_14102_ _14102_/A _14102_/B _14102_/Y vdd gnd NAND2X1
X_11314_ _11314_/A _11314_/B _11314_/C _11314_/D _11314_/Y vdd gnd AOI22X1
XFILL_2__9410_ vdd gnd FILL
X_12294_ _12294_/A _12294_/B _12294_/C _12294_/D _12294_/Y vdd gnd AOI22X1
XFILL_1__7829_ vdd gnd FILL
X_14033_ _14033_/A _14033_/B _14033_/C _14033_/Y vdd gnd OAI21X1
X_11245_ _11245_/A _11245_/B _11245_/Y vdd gnd NAND2X1
XFILL_2__9341_ vdd gnd FILL
XFILL_1__10340_ vdd gnd FILL
X_11176_ _11176_/A _11176_/B _11176_/Y vdd gnd AND2X2
XFILL_2__9272_ vdd gnd FILL
XFILL_1__10271_ vdd gnd FILL
X_10127_ _10127_/A _10127_/Y vdd gnd INVX1
XFILL_1__12010_ vdd gnd FILL
XFILL_2__11561_ vdd gnd FILL
XFILL_0__12740_ vdd gnd FILL
X_10058_ _10058_/A _10058_/B _10058_/C _10058_/Y vdd gnd OAI21X1
XFILL_2__14280_ vdd gnd FILL
XFILL_2__11492_ vdd gnd FILL
XFILL_0__12671_ vdd gnd FILL
XFILL_2__7105_ vdd gnd FILL
X_14866_ _14866_/A _14866_/B _14866_/Y vdd gnd NOR2X1
XFILL_2__13231_ vdd gnd FILL
XFILL_0__14410_ vdd gnd FILL
XFILL_1__13961_ vdd gnd FILL
X_13817_ _13817_/A _13817_/Y vdd gnd INVX1
XFILL_2__13162_ vdd gnd FILL
X_14797_ _14797_/A _14797_/B _14797_/Y vdd gnd NOR2X1
XFILL_1__12912_ vdd gnd FILL
XFILL_0__14341_ vdd gnd FILL
XFILL_1__13892_ vdd gnd FILL
XFILL_0__11553_ vdd gnd FILL
X_13748_ _13748_/A _13748_/B _13748_/C _13748_/Y vdd gnd NAND3X1
XFILL_0__10504_ vdd gnd FILL
XFILL_1__12843_ vdd gnd FILL
XFILL_2__13093_ vdd gnd FILL
XFILL_0__14272_ vdd gnd FILL
XFILL_0__11484_ vdd gnd FILL
X_13679_ _13679_/A _13679_/B _13679_/C _13679_/Y vdd gnd OAI21X1
XFILL_0__13223_ vdd gnd FILL
XFILL_0__10435_ vdd gnd FILL
XFILL_1__12774_ vdd gnd FILL
XFILL_1__11725_ vdd gnd FILL
XFILL_0__13154_ vdd gnd FILL
XFILL_0__10366_ vdd gnd FILL
X_7300_ _7300_/A _7300_/Y vdd gnd INVX1
XFILL_0__9741_ vdd gnd FILL
X_8280_ _8280_/A _8280_/B _8280_/Y vdd gnd OR2X2
XFILL_1__14444_ vdd gnd FILL
XFILL_0__12105_ vdd gnd FILL
XFILL257550x201750 vdd gnd FILL
XFILL_0__13085_ vdd gnd FILL
XFILL_0__10297_ vdd gnd FILL
X_7231_ _7231_/A _7231_/Y vdd gnd INVX1
XFILL_0__9672_ vdd gnd FILL
XFILL_2__9608_ vdd gnd FILL
XFILL_1__10607_ vdd gnd FILL
XFILL_2__12946_ vdd gnd FILL
XFILL_0__12036_ vdd gnd FILL
XFILL_1__14375_ vdd gnd FILL
XFILL_0__8623_ vdd gnd FILL
XFILL_1__11587_ vdd gnd FILL
X_7162_ _7162_/A _7162_/B _7162_/S _7162_/Y vdd gnd MUX2X1
XFILL_2__9539_ vdd gnd FILL
XFILL_1__13326_ vdd gnd FILL
XFILL_1__10538_ vdd gnd FILL
XFILL_0__8554_ vdd gnd FILL
X_7093_ _7093_/A _7093_/B _7093_/C _7093_/Y vdd gnd OAI21X1
XFILL_1__13257_ vdd gnd FILL
XFILL_0__7505_ vdd gnd FILL
XFILL_1__10469_ vdd gnd FILL
XFILL_0__13987_ vdd gnd FILL
XFILL_0__8485_ vdd gnd FILL
XFILL_1__12208_ vdd gnd FILL
XFILL_1__13188_ vdd gnd FILL
XFILL_0__12938_ vdd gnd FILL
XFILL_0__7436_ vdd gnd FILL
XFILL_2__14478_ vdd gnd FILL
XFILL_1__12139_ vdd gnd FILL
X_9803_ _9803_/D _9803_/CLK _9803_/Q vdd gnd DFFPOSX1
XFILL_0__12869_ vdd gnd FILL
XFILL_0__7367_ vdd gnd FILL
XFILL_0__14608_ vdd gnd FILL
X_7995_ _7995_/D _7995_/CLK _7995_/Q vdd gnd DFFPOSX1
XFILL_0__9106_ vdd gnd FILL
X_9734_ _9734_/A _9734_/B _9734_/Y vdd gnd NAND2X1
XFILL_0__7298_ vdd gnd FILL
XFILL_0__9037_ vdd gnd FILL
X_9665_ _9665_/A _9665_/B _9665_/Y vdd gnd NAND2X1
X_8616_ _8616_/A _8616_/B _8616_/C _8616_/Y vdd gnd OAI21X1
XFILL_1__9850_ vdd gnd FILL
X_9596_ _9596_/A _9596_/B _9596_/C _9596_/Y vdd gnd OAI21X1
XFILL_1__8801_ vdd gnd FILL
X_8547_ _8547_/A _8547_/B _8547_/C _8547_/Y vdd gnd NAND3X1
XFILL_0__9939_ vdd gnd FILL
XFILL_1__8732_ vdd gnd FILL
X_8478_ _8478_/A _8478_/B _8478_/Y vdd gnd NOR2X1
XFILL257550x111750 vdd gnd FILL
X_7429_ _7429_/A _7429_/B _7429_/C _7429_/Y vdd gnd NOR3X1
XFILL_1__8663_ vdd gnd FILL
XFILL_1__7614_ vdd gnd FILL
XFILL_1__8594_ vdd gnd FILL
X_11030_ _11030_/A _11030_/B _11030_/C _11030_/Y vdd gnd NAND3X1
XFILL_1__7545_ vdd gnd FILL
XFILL_1__7476_ vdd gnd FILL
XFILL_1__9215_ vdd gnd FILL
X_12981_ _12981_/A _12981_/B _12981_/C _12981_/Y vdd gnd OAI21X1
X_14720_ _14720_/A _14720_/B _14720_/Y vdd gnd OR2X2
XFILL_1__9146_ vdd gnd FILL
X_11932_ _11932_/A _11932_/B _11932_/C _11932_/Y vdd gnd NAND3X1
X_14651_ _14651_/A _14651_/B _14651_/Y vdd gnd NOR2X1
X_11863_ _11863_/A _11863_/B _11863_/Y vdd gnd NOR2X1
XFILL_1__9077_ vdd gnd FILL
X_10814_ _10814_/A _10814_/B _10814_/Y vdd gnd NAND2X1
X_13602_ _13602_/A _13602_/B _13602_/S _13602_/Y vdd gnd MUX2X1
XFILL_1__8028_ vdd gnd FILL
X_14582_ _14582_/A _14582_/B _14582_/C _14582_/Y vdd gnd OAI21X1
X_11794_ _11794_/A _11794_/B _11794_/C _11794_/Y vdd gnd OAI21X1
XFILL_2__9890_ vdd gnd FILL
X_10745_ _10745_/D _10745_/CLK _10745_/Q vdd gnd DFFPOSX1
X_13533_ _13533_/A _13533_/B _13533_/C _13533_/Y vdd gnd OAI21X1
X_13464_ _13464_/D _13464_/CLK _13464_/Q vdd gnd DFFPOSX1
X_10676_ _10676_/A _10676_/B _10676_/Y vdd gnd NAND2X1
XFILL_0__10220_ vdd gnd FILL
XFILL_1__9979_ vdd gnd FILL
XFILL_2__8772_ vdd gnd FILL
X_12415_ _12415_/A _12415_/B _12415_/Y vdd gnd NOR2X1
X_13395_ _13395_/A _13395_/B _13395_/C _13395_/Y vdd gnd OAI21X1
XFILL_1__11510_ vdd gnd FILL
XFILL_0__10151_ vdd gnd FILL
XFILL_1__12490_ vdd gnd FILL
X_12346_ _12346_/A _12346_/B _12346_/C _12346_/Y vdd gnd OAI21X1
XFILL_2__12800_ vdd gnd FILL
XFILL_1__11441_ vdd gnd FILL
XFILL_2__13780_ vdd gnd FILL
XFILL_0__10082_ vdd gnd FILL
X_12277_ _12277_/A _12277_/B _12277_/Y vdd gnd NOR2X1
XFILL_2__12731_ vdd gnd FILL
XFILL_0__13910_ vdd gnd FILL
XFILL_1__11372_ vdd gnd FILL
X_14016_ _14016_/A _14016_/B _14016_/Y vdd gnd NOR2X1
X_11228_ _11228_/A _11228_/B _11228_/Y vdd gnd NAND2X1
XFILL_2__9324_ vdd gnd FILL
XFILL_1__13111_ vdd gnd FILL
XFILL_2__12662_ vdd gnd FILL
XFILL_1__10323_ vdd gnd FILL
XFILL_1__14091_ vdd gnd FILL
XFILL_0__13841_ vdd gnd FILL
X_11159_ _11159_/A _11159_/B _11159_/S _11159_/Y vdd gnd MUX2X1
XFILL_1__13042_ vdd gnd FILL
XFILL_2__9255_ vdd gnd FILL
XFILL_1__10254_ vdd gnd FILL
XFILL_0__13772_ vdd gnd FILL
XFILL_0__10984_ vdd gnd FILL
XFILL_0__8270_ vdd gnd FILL
XFILL_2__14332_ vdd gnd FILL
XFILL_2__9186_ vdd gnd FILL
XFILL_2__11544_ vdd gnd FILL
XFILL_0__12723_ vdd gnd FILL
XFILL_0__7221_ vdd gnd FILL
XFILL_1__10185_ vdd gnd FILL
X_14918_ _14918_/A _14918_/Y vdd gnd BUFX2
XFILL_2__14263_ vdd gnd FILL
XFILL_2__11475_ vdd gnd FILL
XFILL_0__12654_ vdd gnd FILL
XFILL_0__7152_ vdd gnd FILL
X_14849_ _14849_/A _14849_/B _14849_/Y vdd gnd NOR2X1
X_7780_ _7780_/A _7780_/B _7780_/C _7780_/Y vdd gnd OAI21X1
XFILL_0__11605_ vdd gnd FILL
XFILL_1__13944_ vdd gnd FILL
XFILL_0__7083_ vdd gnd FILL
XFILL_0__14324_ vdd gnd FILL
XFILL_1__13875_ vdd gnd FILL
XFILL_0__11536_ vdd gnd FILL
X_9450_ _9450_/A _9450_/B _9450_/Y vdd gnd NOR2X1
XFILL_1__12826_ vdd gnd FILL
XFILL_0__14255_ vdd gnd FILL
X_8401_ _8401_/A _8401_/B _8401_/C _8401_/Y vdd gnd AOI21X1
XFILL_0__11467_ vdd gnd FILL
X_9381_ _9381_/A _9381_/B _9381_/C _9381_/Y vdd gnd OAI21X1
XFILL_2__12027_ vdd gnd FILL
XFILL_0__13206_ vdd gnd FILL
XFILL_0__10418_ vdd gnd FILL
XFILL_0_BUFX2_insert370 vdd gnd FILL
XFILL_1__12757_ vdd gnd FILL
X_8332_ _8332_/A _8332_/B _8332_/C _8332_/Y vdd gnd AOI21X1
XFILL_0__11398_ vdd gnd FILL
XFILL_0_BUFX2_insert381 vdd gnd FILL
XFILL_1__11708_ vdd gnd FILL
XFILL_0__13137_ vdd gnd FILL
XFILL_0__10349_ vdd gnd FILL
XFILL_1__12688_ vdd gnd FILL
XFILL_0__9724_ vdd gnd FILL
X_8263_ _8263_/A _8263_/B _8263_/C _8263_/Y vdd gnd NAND3X1
XFILL_1__14427_ vdd gnd FILL
XFILL_2__13978_ vdd gnd FILL
XFILL_0__13068_ vdd gnd FILL
X_7214_ _7214_/A _7214_/B _7214_/C _7214_/Y vdd gnd AOI21X1
XFILL_0__9655_ vdd gnd FILL
X_8194_ _8194_/A _8194_/B _8194_/C _8194_/Y vdd gnd OAI21X1
XFILL_2__12929_ vdd gnd FILL
XFILL_1__14358_ vdd gnd FILL
XFILL_0__12019_ vdd gnd FILL
XFILL_0__8606_ vdd gnd FILL
X_7145_ _7145_/A _7145_/B _7145_/Y vdd gnd NAND2X1
XFILL_0__9586_ vdd gnd FILL
XFILL_1__13309_ vdd gnd FILL
XFILL_1__14289_ vdd gnd FILL
XFILL_1__7330_ vdd gnd FILL
XFILL_0__8537_ vdd gnd FILL
X_7076_ _7076_/A _7076_/B _7076_/Y vdd gnd NOR2X1
XFILL_1__7261_ vdd gnd FILL
XFILL_0__8468_ vdd gnd FILL
XFILL_1__9000_ vdd gnd FILL
XFILL_0__7419_ vdd gnd FILL
XFILL_1__7192_ vdd gnd FILL
XFILL_0__8399_ vdd gnd FILL
X_7978_ _7978_/D _7978_/CLK _7978_/Q vdd gnd DFFPOSX1
X_9717_ _9717_/A _9717_/B _9717_/C _9717_/Y vdd gnd OAI21X1
XFILL_1__9902_ vdd gnd FILL
X_9648_ _9648_/A _9648_/B _9648_/Y vdd gnd NOR2X1
X_10530_ _10530_/A _10530_/B _10530_/Y vdd gnd NOR2X1
X_9579_ _9579_/A _9579_/Y vdd gnd INVX1
X_10461_ _10461_/A _10461_/B _10461_/Y vdd gnd NAND2X1
X_12200_ _12200_/A _12200_/B _12200_/C _12200_/Y vdd gnd OAI21X1
X_13180_ _13180_/A _13180_/Y vdd gnd INVX1
X_10392_ _10392_/A _10392_/B _10392_/Y vdd gnd NOR2X1
XFILL_1__8715_ vdd gnd FILL
XFILL_1__9695_ vdd gnd FILL
X_12131_ _12131_/A _12131_/B _12131_/C _12131_/Y vdd gnd OAI21X1
XFILL_1__8646_ vdd gnd FILL
XFILL_2_CLKBUF1_insert101 vdd gnd FILL
X_12062_ _12062_/A _12062_/B _12062_/C _12062_/Y vdd gnd NAND3X1
XFILL_2__7370_ vdd gnd FILL
XFILL_1__8577_ vdd gnd FILL
X_11013_ _11013_/A _11013_/B _11013_/Y vdd gnd NAND2X1
XFILL_1__7528_ vdd gnd FILL
XFILL_2__9040_ vdd gnd FILL
XFILL_1__7459_ vdd gnd FILL
X_12964_ _12964_/A _12964_/B _12964_/Y vdd gnd NAND2X1
X_14703_ _14703_/A _14703_/Y vdd gnd INVX1
X_11915_ _11915_/A _11915_/B _11915_/Y vdd gnd AND2X2
XFILL_1__9129_ vdd gnd FILL
XFILL_2__11260_ vdd gnd FILL
X_12895_ _12895_/A _12895_/B _12895_/C _12895_/Y vdd gnd NAND3X1
XFILL_1__11990_ vdd gnd FILL
X_14634_ _14634_/A _14634_/B _14634_/C _14634_/Y vdd gnd AOI21X1
X_11846_ _11846_/A _11846_/B _11846_/C _11846_/Y vdd gnd OAI21X1
XFILL_1__10941_ vdd gnd FILL
XFILL_2__11191_ vdd gnd FILL
XFILL_0__12370_ vdd gnd FILL
X_14565_ _14565_/A _14565_/B _14565_/C _14565_/Y vdd gnd OAI21X1
X_11777_ _11777_/A _11777_/Y vdd gnd INVX8
XFILL_1__13660_ vdd gnd FILL
XFILL_0__11321_ vdd gnd FILL
XFILL_1__10872_ vdd gnd FILL
X_10728_ _10728_/D _10728_/CLK _10728_/Q vdd gnd DFFPOSX1
X_13516_ _13516_/A _13516_/B _13516_/C _13516_/Y vdd gnd OAI21X1
X_14496_ _14496_/A _14496_/B _14496_/Y vdd gnd NAND2X1
XFILL_0__14040_ vdd gnd FILL
XFILL_0__11252_ vdd gnd FILL
XFILL_1__13591_ vdd gnd FILL
X_13447_ _13447_/D _13447_/CLK _13447_/Q vdd gnd DFFPOSX1
X_10659_ _10659_/A _10659_/B _10659_/C _10659_/Y vdd gnd OAI21X1
XFILL_2__13901_ vdd gnd FILL
XFILL_0__10203_ vdd gnd FILL
XFILL_0__11183_ vdd gnd FILL
XFILL_0__7770_ vdd gnd FILL
X_13378_ _13378_/A _13378_/B _13378_/Y vdd gnd NAND2X1
XFILL_2__7706_ vdd gnd FILL
XFILL_0__10134_ vdd gnd FILL
XFILL_2__13832_ vdd gnd FILL
XFILL_2__8686_ vdd gnd FILL
XFILL_1__12473_ vdd gnd FILL
X_12329_ _12329_/A _12329_/B _12329_/C _12329_/Y vdd gnd OAI21X1
XFILL_2__7637_ vdd gnd FILL
XFILL_1__11424_ vdd gnd FILL
XFILL_0__10065_ vdd gnd FILL
XFILL_2__13763_ vdd gnd FILL
XFILL_0__9440_ vdd gnd FILL
XFILL_2__12714_ vdd gnd FILL
XFILL_1__14143_ vdd gnd FILL
XFILL_1_BUFX2_insert15 vdd gnd FILL
XFILL_1__11355_ vdd gnd FILL
XFILL_2__13694_ vdd gnd FILL
XFILL_0__9371_ vdd gnd FILL
XFILL_1_BUFX2_insert26 vdd gnd FILL
XFILL_2__9307_ vdd gnd FILL
XFILL_1__10306_ vdd gnd FILL
XFILL_2__12645_ vdd gnd FILL
XFILL_0__13824_ vdd gnd FILL
XFILL_1__14074_ vdd gnd FILL
XFILL_0__8322_ vdd gnd FILL
XFILL_1__11286_ vdd gnd FILL
X_8950_ _8950_/A _8950_/B _8950_/C _8950_/Y vdd gnd OAI21X1
XFILL_2__9238_ vdd gnd FILL
XFILL_1__13025_ vdd gnd FILL
XFILL_1__10237_ vdd gnd FILL
XFILL_0__13755_ vdd gnd FILL
XFILL_0__10967_ vdd gnd FILL
X_7901_ _7901_/A _7901_/B _7901_/C _7901_/Y vdd gnd OAI21X1
XFILL_0__8253_ vdd gnd FILL
X_8881_ _8881_/D _8881_/CLK _8881_/Q vdd gnd DFFPOSX1
XFILL_2__11527_ vdd gnd FILL
XFILL_2__9169_ vdd gnd FILL
XFILL_0__12706_ vdd gnd FILL
XFILL_1__10168_ vdd gnd FILL
XFILL_0__7204_ vdd gnd FILL
XFILL_0__13686_ vdd gnd FILL
X_7832_ _7832_/A _7832_/B _7832_/Y vdd gnd NAND2X1
XFILL_0__8184_ vdd gnd FILL
XFILL_0__10898_ vdd gnd FILL
XFILL_2__11458_ vdd gnd FILL
XFILL_0__12637_ vdd gnd FILL
XFILL_0__7135_ vdd gnd FILL
XFILL_1__10099_ vdd gnd FILL
X_7763_ _7763_/A _7763_/Y vdd gnd INVX1
XFILL_1_CLKBUF1_insert38 vdd gnd FILL
XFILL_1__13927_ vdd gnd FILL
XFILL_1_CLKBUF1_insert49 vdd gnd FILL
XFILL_2__11389_ vdd gnd FILL
X_9502_ _9502_/A _9502_/Y vdd gnd INVX1
X_7694_ _7694_/A _7694_/Y vdd gnd INVX1
XFILL_0__14307_ vdd gnd FILL
XFILL_0__11519_ vdd gnd FILL
XFILL_1__13858_ vdd gnd FILL
X_9433_ _9433_/A _9433_/B _9433_/C _9433_/Y vdd gnd AOI21X1
XFILL_0__12499_ vdd gnd FILL
XFILL_0__14238_ vdd gnd FILL
XFILL_1__12809_ vdd gnd FILL
XFILL_1__13789_ vdd gnd FILL
X_9364_ _9364_/A _9364_/B _9364_/Y vdd gnd NAND2X1
X_8315_ _8315_/A _8315_/B _8315_/C _8315_/Y vdd gnd OAI21X1
X_9295_ _9295_/A _9295_/B _9295_/S _9295_/Y vdd gnd MUX2X1
XFILL_0__9707_ vdd gnd FILL
XFILL_1__8500_ vdd gnd FILL
X_8246_ _8246_/A _8246_/B _8246_/C _8246_/Y vdd gnd AOI21X1
XFILL_1__9480_ vdd gnd FILL
XFILL_0__7899_ vdd gnd FILL
XFILL_0__9638_ vdd gnd FILL
XFILL_1__8431_ vdd gnd FILL
X_8177_ _8177_/A _8177_/B _8177_/Y vdd gnd NAND2X1
X_7128_ _7128_/A _7128_/B _7128_/C _7128_/D _7128_/Y vdd gnd AOI22X1
XFILL_1__8362_ vdd gnd FILL
XFILL_0__9569_ vdd gnd FILL
XFILL_1__7313_ vdd gnd FILL
XFILL_1__8293_ vdd gnd FILL
XFILL_1__7244_ vdd gnd FILL
XFILL_1__7175_ vdd gnd FILL
X_11700_ _11700_/A _11700_/Y vdd gnd INVX2
X_12680_ _12680_/A _12680_/B _12680_/C _12680_/Y vdd gnd OAI21X1
X_11631_ _11631_/D _11631_/CLK _11631_/Q vdd gnd DFFPOSX1
X_14350_ _14350_/A _14350_/B _14350_/C _14350_/Y vdd gnd NAND3X1
X_11562_ _11562_/A _11562_/B _11562_/Y vdd gnd NAND2X1
X_10513_ _10513_/A _10513_/B _10513_/Y vdd gnd OR2X2
X_13301_ _13301_/A _13301_/B _13301_/Y vdd gnd NAND2X1
X_14281_ _14281_/A _14281_/B _14281_/Y vdd gnd AND2X2
X_11493_ _11493_/A _11493_/B _11493_/C _11493_/Y vdd gnd NAND3X1
X_13232_ _13232_/A _13232_/B _13232_/Y vdd gnd OR2X2
X_10444_ _10444_/A _10444_/B _10444_/Y vdd gnd NOR2X1
XFILL_1__9747_ vdd gnd FILL
X_13163_ _13163_/A _13163_/Y vdd gnd INVX1
X_10375_ _10375_/A _10375_/Y vdd gnd INVX1
XFILL_1__9678_ vdd gnd FILL
X_12114_ _12114_/A _12114_/B _12114_/Y vdd gnd NAND2X1
X_13094_ _13094_/A _13094_/B _13094_/C _13094_/Y vdd gnd OAI21X1
XFILL_2__7422_ vdd gnd FILL
XFILL_1__8629_ vdd gnd FILL
X_12045_ _12045_/A _12045_/B _12045_/Y vdd gnd NAND2X1
XFILL_2__7353_ vdd gnd FILL
XFILL_1__11140_ vdd gnd FILL
XFILL_0__11870_ vdd gnd FILL
XFILL_2__7284_ vdd gnd FILL
XFILL_1__11071_ vdd gnd FILL
XFILL_0__10821_ vdd gnd FILL
XFILL_1__10022_ vdd gnd FILL
XFILL_2_BUFX2_insert251 vdd gnd FILL
X_13996_ _13996_/A _13996_/B _13996_/Y vdd gnd NAND2X1
XFILL_0__13540_ vdd gnd FILL
X_12947_ _12947_/A _12947_/B _12947_/C _12947_/Y vdd gnd NAND3X1
XFILL_2_BUFX2_insert284 vdd gnd FILL
XFILL_1__14830_ vdd gnd FILL
XFILL_0__10683_ vdd gnd FILL
X_12878_ _12878_/A _12878_/B _12878_/C _12878_/Y vdd gnd NAND3X1
XFILL_1__14761_ vdd gnd FILL
XFILL_0__12422_ vdd gnd FILL
XFILL_1__11973_ vdd gnd FILL
X_14617_ _14617_/A _14617_/B _14617_/C _14617_/Y vdd gnd OAI21X1
X_11829_ _11829_/A _11829_/B _11829_/S _11829_/Y vdd gnd MUX2X1
XFILL_1__13712_ vdd gnd FILL
XFILL_1__10924_ vdd gnd FILL
XFILL_1__14692_ vdd gnd FILL
XFILL_0__12353_ vdd gnd FILL
XFILL_0__8940_ vdd gnd FILL
X_14548_ _14548_/D _14548_/CLK _14548_/Q vdd gnd DFFPOSX1
XFILL_2__10125_ vdd gnd FILL
XBUFX2_insert250 BUFX2_insert250/A BUFX2_insert250/Y vdd gnd BUFX2
XFILL_1__13643_ vdd gnd FILL
XFILL_0__11304_ vdd gnd FILL
XBUFX2_insert261 BUFX2_insert261/A BUFX2_insert261/Y vdd gnd BUFX2
XFILL_1__10855_ vdd gnd FILL
XBUFX2_insert272 BUFX2_insert272/A BUFX2_insert272/Y vdd gnd BUFX2
XFILL_0__12284_ vdd gnd FILL
XBUFX2_insert283 BUFX2_insert283/A BUFX2_insert283/Y vdd gnd BUFX2
X_14479_ _14479_/A _14479_/Y vdd gnd INVX1
XFILL_2__10056_ vdd gnd FILL
XBUFX2_insert294 BUFX2_insert294/A BUFX2_insert294/Y vdd gnd BUFX2
XFILL_0__14023_ vdd gnd FILL
XFILL_0__11235_ vdd gnd FILL
XFILL_1__13574_ vdd gnd FILL
XFILL_1__10786_ vdd gnd FILL
XFILL_0__7822_ vdd gnd FILL
XFILL_1__12525_ vdd gnd FILL
XFILL_0__11166_ vdd gnd FILL
X_8100_ _8100_/A _8100_/B _8100_/Y vdd gnd NAND2X1
X_9080_ _9080_/A _9080_/Y vdd gnd INVX2
XFILL_0__7753_ vdd gnd FILL
XFILL_2__13815_ vdd gnd FILL
XFILL_0__10117_ vdd gnd FILL
XFILL_1__12456_ vdd gnd FILL
X_8031_ _8031_/A _8031_/B _8031_/C _8031_/Y vdd gnd AOI21X1
XFILL_0__11097_ vdd gnd FILL
XFILL_0__7684_ vdd gnd FILL
XFILL_1__11407_ vdd gnd FILL
XFILL_2__13746_ vdd gnd FILL
XFILL_2__10958_ vdd gnd FILL
XFILL_0__10048_ vdd gnd FILL
XFILL_1__12387_ vdd gnd FILL
XFILL_0__9423_ vdd gnd FILL
XFILL256650x252150 vdd gnd FILL
XFILL257250x237750 vdd gnd FILL
XFILL_1__14126_ vdd gnd FILL
XFILL_1__11338_ vdd gnd FILL
XFILL_0__14856_ vdd gnd FILL
XFILL_2__10889_ vdd gnd FILL
XFILL_2__13677_ vdd gnd FILL
XFILL_0__9354_ vdd gnd FILL
X_9982_ _9982_/A _9982_/B _9982_/S _9982_/Y vdd gnd MUX2X1
XFILL_0__13807_ vdd gnd FILL
XFILL_1__14057_ vdd gnd FILL
XFILL_1__11269_ vdd gnd FILL
XFILL_0__14787_ vdd gnd FILL
XFILL_0__8305_ vdd gnd FILL
XFILL_0__9285_ vdd gnd FILL
X_8933_ _8933_/A _8933_/B _8933_/C _8933_/D _8933_/Y vdd gnd AOI22X1
XFILL_0__11999_ vdd gnd FILL
XFILL_1__13008_ vdd gnd FILL
XFILL_0__13738_ vdd gnd FILL
XFILL_0__8236_ vdd gnd FILL
X_8864_ _8864_/D _8864_/CLK _8864_/Q vdd gnd DFFPOSX1
XFILL_0__13669_ vdd gnd FILL
X_7815_ _7815_/A _7815_/B _7815_/C _7815_/Y vdd gnd OAI21X1
XFILL_0__8167_ vdd gnd FILL
X_8795_ _8795_/A _8795_/Y vdd gnd INVX1
XFILL_0__7118_ vdd gnd FILL
X_7746_ _7746_/A _7746_/B _7746_/C _7746_/Y vdd gnd OAI21X1
XFILL_0__8098_ vdd gnd FILL
XFILL_1__8980_ vdd gnd FILL
X_7677_ _7677_/A _7677_/B _7677_/C _7677_/Y vdd gnd AOI21X1
X_9416_ _9416_/A _9416_/B _9416_/Y vdd gnd NOR2X1
XFILL_1__7862_ vdd gnd FILL
XFILL_1__9601_ vdd gnd FILL
X_9347_ _9347_/A _9347_/B _9347_/C _9347_/Y vdd gnd OAI21X1
XFILL_1__7793_ vdd gnd FILL
XFILL_1__9532_ vdd gnd FILL
X_9278_ _9278_/A _9278_/B _9278_/C _9278_/Y vdd gnd AOI21X1
X_10160_ _10160_/A _10160_/B _10160_/C _10160_/Y vdd gnd NAND3X1
X_8229_ _8229_/A _8229_/B _8229_/C _8229_/Y vdd gnd NAND3X1
XFILL_1__9463_ vdd gnd FILL
X_10091_ _10091_/A _10091_/B _10091_/C _10091_/Y vdd gnd OAI21X1
XFILL_1__8414_ vdd gnd FILL
XFILL257250x147750 vdd gnd FILL
XFILL_1__9394_ vdd gnd FILL
XFILL_1__8345_ vdd gnd FILL
X_13850_ _13850_/A _13850_/B _13850_/Y vdd gnd NAND2X1
XFILL_1__8276_ vdd gnd FILL
X_12801_ _12801_/A _12801_/B _12801_/Y vdd gnd NAND2X1
X_10993_ _10993_/A _10993_/B _10993_/C _10993_/Y vdd gnd OAI21X1
XFILL_1__7227_ vdd gnd FILL
X_13781_ _13781_/A _13781_/Y vdd gnd INVX1
XFILL_1_BUFX2_insert203 vdd gnd FILL
XFILL_1_BUFX2_insert214 vdd gnd FILL
XFILL_1_BUFX2_insert225 vdd gnd FILL
X_12732_ _12732_/A _12732_/B _12732_/C _12732_/Y vdd gnd OAI21X1
XFILL_1__7158_ vdd gnd FILL
XFILL_1_BUFX2_insert236 vdd gnd FILL
XFILL257250x190950 vdd gnd FILL
XFILL_1_BUFX2_insert247 vdd gnd FILL
XFILL_1_BUFX2_insert258 vdd gnd FILL
XFILL_1_BUFX2_insert269 vdd gnd FILL
XCLKBUF1_insert29 CLKBUF1_insert29/A CLKBUF1_insert29/Y vdd gnd CLKBUF1
X_12663_ _12663_/A _12663_/B _12663_/C _12663_/D _12663_/Y vdd gnd AOI22X1
XFILL_1__7089_ vdd gnd FILL
X_14402_ _14402_/A _14402_/B _14402_/Y vdd gnd NAND2X1
X_11614_ _11614_/D _11614_/CLK _11614_/Q vdd gnd DFFPOSX1
XFILL_2__9710_ vdd gnd FILL
X_12594_ _12594_/D _12594_/CLK _12594_/Q vdd gnd DFFPOSX1
XFILL_0_CLKBUF1_insert384 vdd gnd FILL
X_14333_ _14333_/A _14333_/B _14333_/C _14333_/Y vdd gnd OAI21X1
X_11545_ _11545_/A _11545_/B _11545_/Y vdd gnd NAND2X1
XFILL_2__9641_ vdd gnd FILL
XFILL_1__10640_ vdd gnd FILL
X_14264_ _14264_/A _14264_/B _14264_/C _14264_/Y vdd gnd OAI21X1
X_11476_ _11476_/A _11476_/B _11476_/C _11476_/Y vdd gnd OAI21X1
XFILL_0__11020_ vdd gnd FILL
XFILL_2__9572_ vdd gnd FILL
XFILL_1__10571_ vdd gnd FILL
X_13215_ _13215_/A _13215_/B _13215_/Y vdd gnd NAND2X1
X_10427_ _10427_/A _10427_/Y vdd gnd INVX1
XFILL_1__12310_ vdd gnd FILL
X_14195_ _14195_/D _14195_/CLK _14195_/Q vdd gnd DFFPOSX1
XFILL_1__13290_ vdd gnd FILL
X_13146_ _13146_/A _13146_/B _13146_/C _13146_/Y vdd gnd NAND3X1
X_10358_ _10358_/A _10358_/B _10358_/Y vdd gnd NOR2X1
XFILL_1__12241_ vdd gnd FILL
XFILL_2__10812_ vdd gnd FILL
XFILL_0__12971_ vdd gnd FILL
X_13077_ _13077_/A _13077_/B _13077_/Y vdd gnd NOR2X1
X_10289_ _10289_/A _10289_/B _10289_/Y vdd gnd OR2X2
XFILL_2__7405_ vdd gnd FILL
XFILL_0__14710_ vdd gnd FILL
XFILL_0__11922_ vdd gnd FILL
XFILL_1__12172_ vdd gnd FILL
X_12028_ _12028_/A _12028_/B _12028_/C _12028_/Y vdd gnd AOI21X1
XFILL_2__7336_ vdd gnd FILL
XFILL_1__11123_ vdd gnd FILL
XFILL_0__14641_ vdd gnd FILL
XFILL_0__11853_ vdd gnd FILL
XFILL_2__12413_ vdd gnd FILL
XFILL_1__11054_ vdd gnd FILL
XFILL_0__10804_ vdd gnd FILL
XFILL_2__7267_ vdd gnd FILL
XFILL_0__14572_ vdd gnd FILL
XFILL_0__9070_ vdd gnd FILL
XFILL_0__11784_ vdd gnd FILL
X_13979_ _13979_/A _13979_/Y vdd gnd INVX1
XFILL_1__10005_ vdd gnd FILL
XFILL_2__12344_ vdd gnd FILL
XFILL_2__7198_ vdd gnd FILL
XFILL_0__13523_ vdd gnd FILL
XFILL_0__8021_ vdd gnd FILL
XFILL_1__14813_ vdd gnd FILL
XFILL_2__12275_ vdd gnd FILL
X_7600_ _7600_/A _7600_/Y vdd gnd INVX1
XFILL_0__10666_ vdd gnd FILL
X_8580_ _8580_/A _8580_/B _8580_/C _8580_/Y vdd gnd AOI21X1
XFILL_0__12405_ vdd gnd FILL
XFILL_1__14744_ vdd gnd FILL
XFILL_1__11956_ vdd gnd FILL
XFILL_0__13385_ vdd gnd FILL
X_7531_ _7531_/A _7531_/B _7531_/C _7531_/Y vdd gnd OAI21X1
XFILL_0__10597_ vdd gnd FILL
XFILL257250x212550 vdd gnd FILL
XFILL_0__9972_ vdd gnd FILL
XFILL_1__10907_ vdd gnd FILL
XFILL_0__12336_ vdd gnd FILL
XFILL_1__14675_ vdd gnd FILL
XFILL_1__11887_ vdd gnd FILL
XFILL_0__8923_ vdd gnd FILL
X_7462_ _7462_/A _7462_/B _7462_/C _7462_/Y vdd gnd OAI21X1
XFILL_2__10108_ vdd gnd FILL
XFILL_1__10838_ vdd gnd FILL
XFILL_1__13626_ vdd gnd FILL
X_9201_ _9201_/A _9201_/B _9201_/Y vdd gnd NOR2X1
XFILL_0__12267_ vdd gnd FILL
XFILL_0__14006_ vdd gnd FILL
X_7393_ _7393_/A _7393_/B _7393_/C _7393_/Y vdd gnd OAI21X1
XFILL_2__10039_ vdd gnd FILL
XFILL_2__14916_ vdd gnd FILL
XFILL_0__11218_ vdd gnd FILL
XFILL_1__13557_ vdd gnd FILL
XFILL_1__10769_ vdd gnd FILL
X_9132_ _9132_/A _9132_/B _9132_/C _9132_/Y vdd gnd AOI21X1
XFILL_0__7805_ vdd gnd FILL
XFILL_0__12198_ vdd gnd FILL
XFILL_0__8785_ vdd gnd FILL
XFILL_1__12508_ vdd gnd FILL
XFILL_0__11149_ vdd gnd FILL
X_9063_ _9063_/A _9063_/B _9063_/C _9063_/Y vdd gnd AOI21X1
XFILL_0__7736_ vdd gnd FILL
XFILL_1__12439_ vdd gnd FILL
X_8014_ _8014_/A _8014_/Y vdd gnd INVX1
XFILL_0__7667_ vdd gnd FILL
XFILL_0__14908_ vdd gnd FILL
XFILL_0__9406_ vdd gnd FILL
XFILL_0__7598_ vdd gnd FILL
XFILL_1__14109_ vdd gnd FILL
XFILL_0__14839_ vdd gnd FILL
XFILL_1__8130_ vdd gnd FILL
XFILL_0__9337_ vdd gnd FILL
X_9965_ _9965_/A _9965_/B _9965_/S _9965_/Y vdd gnd MUX2X1
XFILL_1__8061_ vdd gnd FILL
XFILL_0__9268_ vdd gnd FILL
X_8916_ _8916_/D _8916_/CLK _8916_/Q vdd gnd DFFPOSX1
X_9896_ _9896_/A _9896_/B _9896_/Y vdd gnd NOR2X1
XFILL_0__8219_ vdd gnd FILL
XFILL_0__9199_ vdd gnd FILL
X_8847_ _8847_/D _8847_/CLK _8847_/Q vdd gnd DFFPOSX1
X_8778_ _8778_/A _8778_/B _8778_/Y vdd gnd NAND2X1
X_7729_ _7729_/A _7729_/B _7729_/Y vdd gnd NOR2X1
XFILL257250x122550 vdd gnd FILL
XFILL_1__8963_ vdd gnd FILL
XFILL_1__7914_ vdd gnd FILL
X_11330_ _11330_/A _11330_/B _11330_/C _11330_/Y vdd gnd OAI21X1
XFILL_1__7845_ vdd gnd FILL
X_11261_ _11261_/A _11261_/Y vdd gnd INVX1
XFILL_1__7776_ vdd gnd FILL
X_10212_ _10212_/A _10212_/B _10212_/Y vdd gnd NOR2X1
X_13000_ _13000_/A _13000_/B _13000_/S _13000_/Y vdd gnd MUX2X1
XFILL_1__9515_ vdd gnd FILL
X_11192_ _11192_/A _11192_/Y vdd gnd INVX1
X_10143_ _10143_/A _10143_/B _10143_/Y vdd gnd NAND2X1
XFILL_1__9446_ vdd gnd FILL
X_10074_ _10074_/A _10074_/B _10074_/C _10074_/Y vdd gnd AOI21X1
XFILL_1__9377_ vdd gnd FILL
X_13902_ _13902_/A _13902_/B _13902_/Y vdd gnd NAND2X1
X_14882_ _14882_/D _14882_/CLK _14882_/Q vdd gnd DFFPOSX1
XFILL_1__8328_ vdd gnd FILL
X_13833_ _13833_/A _13833_/Y vdd gnd INVX1
XFILL_1__8259_ vdd gnd FILL
X_13764_ _13764_/A _13764_/B _13764_/C _13764_/Y vdd gnd OAI21X1
X_10976_ _10976_/A _10976_/Y vdd gnd INVX1
XFILL_0__10520_ vdd gnd FILL
X_12715_ _12715_/A _12715_/B _12715_/S _12715_/Y vdd gnd MUX2X1
X_13695_ _13695_/A _13695_/B _13695_/C _13695_/Y vdd gnd NAND3X1
XFILL_2__12060_ vdd gnd FILL
XFILL_1__11810_ vdd gnd FILL
XFILL_0__10451_ vdd gnd FILL
XFILL_1__12790_ vdd gnd FILL
X_12646_ _12646_/A _12646_/B _12646_/Y vdd gnd NAND2X1
XFILL_1__11741_ vdd gnd FILL
XFILL_0__13170_ vdd gnd FILL
XFILL_0__10382_ vdd gnd FILL
X_12577_ _12577_/D _12577_/CLK _12577_/Q vdd gnd DFFPOSX1
XFILL_1__14460_ vdd gnd FILL
XFILL_0__12121_ vdd gnd FILL
X_14316_ _14316_/A _14316_/B _14316_/Y vdd gnd NAND2X1
X_11528_ _11528_/A _11528_/B _11528_/Y vdd gnd NAND2X1
XFILL_2__9624_ vdd gnd FILL
XFILL_1__13411_ vdd gnd FILL
XFILL_1__10623_ vdd gnd FILL
XFILL_2__12962_ vdd gnd FILL
XFILL_0__12052_ vdd gnd FILL
XFILL_1__14391_ vdd gnd FILL
X_14247_ _14247_/A _14247_/B _14247_/Y vdd gnd NAND2X1
XFILL_2__14701_ vdd gnd FILL
X_11459_ _11459_/A _11459_/Y vdd gnd INVX1
XFILL_0__11003_ vdd gnd FILL
XFILL_2__9555_ vdd gnd FILL
XFILL_1__13342_ vdd gnd FILL
XFILL_1__10554_ vdd gnd FILL
XFILL_2__12893_ vdd gnd FILL
XFILL_0__8570_ vdd gnd FILL
X_14178_ _14178_/D _14178_/CLK _14178_/Q vdd gnd DFFPOSX1
XFILL_2__9486_ vdd gnd FILL
XFILL_1__13273_ vdd gnd FILL
XFILL_1__10485_ vdd gnd FILL
X_13129_ _13129_/A _13129_/B _13129_/C _13129_/Y vdd gnd NAND3X1
XFILL_0__7521_ vdd gnd FILL
XFILL_1__12224_ vdd gnd FILL
XFILL_0__12954_ vdd gnd FILL
XFILL_0__7452_ vdd gnd FILL
XFILL_0__11905_ vdd gnd FILL
XFILL_1__12155_ vdd gnd FILL
XFILL_2__14494_ vdd gnd FILL
XFILL_0__12885_ vdd gnd FILL
XFILL_0__7383_ vdd gnd FILL
XFILL_1__11106_ vdd gnd FILL
XFILL_0__14624_ vdd gnd FILL
XFILL_0__11836_ vdd gnd FILL
XFILL_1__12086_ vdd gnd FILL
XFILL_0__9122_ vdd gnd FILL
X_9750_ _9750_/A _9750_/B _9750_/Y vdd gnd NAND2X1
XFILL_1__11037_ vdd gnd FILL
XFILL_0__11767_ vdd gnd FILL
XFILL_0__9053_ vdd gnd FILL
X_8701_ _8701_/A _8701_/B _8701_/Y vdd gnd NOR2X1
X_9681_ _9681_/A _9681_/B _9681_/Y vdd gnd NAND2X1
XFILL_2__12327_ vdd gnd FILL
XFILL_0__13506_ vdd gnd FILL
XFILL_0__8004_ vdd gnd FILL
XFILL_0__14486_ vdd gnd FILL
X_8632_ _8632_/A _8632_/Y vdd gnd INVX1
XFILL_0__11698_ vdd gnd FILL
XFILL_2__12258_ vdd gnd FILL
XFILL_0__10649_ vdd gnd FILL
XFILL_1__12988_ vdd gnd FILL
X_8563_ _8563_/A _8563_/B _8563_/Y vdd gnd NAND2X1
XFILL_1__14727_ vdd gnd FILL
XFILL_2__12189_ vdd gnd FILL
XFILL_1__11939_ vdd gnd FILL
XFILL_0__13368_ vdd gnd FILL
X_7514_ _7514_/A _7514_/B _7514_/Y vdd gnd NAND2X1
XFILL_0__9955_ vdd gnd FILL
X_8494_ _8494_/A _8494_/B _8494_/C _8494_/Y vdd gnd OAI21X1
XFILL_0__12319_ vdd gnd FILL
XFILL_1__14658_ vdd gnd FILL
XFILL_0__13299_ vdd gnd FILL
X_7445_ _7445_/A _7445_/B _7445_/Y vdd gnd NAND2X1
XFILL_0__9886_ vdd gnd FILL
XFILL_1__13609_ vdd gnd FILL
XFILL_1__14589_ vdd gnd FILL
XFILL_1__7630_ vdd gnd FILL
XFILL_0__8837_ vdd gnd FILL
X_7376_ _7376_/A _7376_/Y vdd gnd INVX1
X_9115_ _9115_/A _9115_/B _9115_/C _9115_/Y vdd gnd OAI21X1
XFILL_1__7561_ vdd gnd FILL
XFILL_0__8768_ vdd gnd FILL
XFILL_1__9300_ vdd gnd FILL
X_9046_ _9046_/A _9046_/B _9046_/C _9046_/Y vdd gnd NAND3X1
XFILL_0__7719_ vdd gnd FILL
XFILL_1__7492_ vdd gnd FILL
XFILL_0__8699_ vdd gnd FILL
XFILL_1__9231_ vdd gnd FILL
XFILL_1__9162_ vdd gnd FILL
XFILL_1__8113_ vdd gnd FILL
XFILL_1__9093_ vdd gnd FILL
X_9948_ _9948_/A _9948_/B _9948_/Y vdd gnd NAND2X1
X_10830_ _10830_/A _10830_/Y vdd gnd INVX1
XFILL_1__8044_ vdd gnd FILL
X_9879_ _9879_/A _9879_/B _9879_/C _9879_/Y vdd gnd AOI21X1
X_10761_ _10761_/D _10761_/CLK _10761_/Q vdd gnd DFFPOSX1
X_12500_ _12500_/A _12500_/B _12500_/Y vdd gnd NAND2X1
X_10692_ _10692_/D _10692_/CLK _10692_/Q vdd gnd DFFPOSX1
X_13480_ _13480_/D _13480_/CLK _13480_/Q vdd gnd DFFPOSX1
XFILL_1__9995_ vdd gnd FILL
X_12431_ _12431_/A _12431_/B _12431_/Y vdd gnd OR2X2
XFILL_1__8946_ vdd gnd FILL
X_12362_ _12362_/A _12362_/B _12362_/Y vdd gnd NAND2X1
XFILL_2__7670_ vdd gnd FILL
X_14101_ _14101_/A _14101_/B _14101_/Y vdd gnd NOR2X1
X_11313_ _11313_/A _11313_/B _11313_/C _11313_/Y vdd gnd AOI21X1
X_12293_ _12293_/A _12293_/B _12293_/Y vdd gnd NOR2X1
XFILL_1__7828_ vdd gnd FILL
X_14032_ _14032_/A _14032_/B _14032_/C _14032_/D _14032_/Y vdd gnd AOI22X1
X_11244_ _11244_/A _11244_/B _11244_/Y vdd gnd NAND2X1
XFILL_1__7759_ vdd gnd FILL
X_11175_ _11175_/A _11175_/B _11175_/C _11175_/Y vdd gnd NAND3X1
XFILL_1__10270_ vdd gnd FILL
X_10126_ _10126_/A _10126_/B _10126_/C _10126_/Y vdd gnd AOI21X1
XFILL_1__9429_ vdd gnd FILL
XFILL_2__8222_ vdd gnd FILL
X_10057_ _10057_/A _10057_/B _10057_/Y vdd gnd NAND2X1
XFILL_2__10511_ vdd gnd FILL
XFILL_2__8153_ vdd gnd FILL
XFILL_0__12670_ vdd gnd FILL
X_14865_ _14865_/A _14865_/B _14865_/C _14865_/Y vdd gnd AOI21X1
XFILL_2__10442_ vdd gnd FILL
XFILL_2__8084_ vdd gnd FILL
XFILL_1__13960_ vdd gnd FILL
X_13816_ _13816_/A _13816_/B _13816_/Y vdd gnd NAND2X1
X_14796_ _14796_/A _14796_/B _14796_/Y vdd gnd NAND2X1
XFILL_0__14340_ vdd gnd FILL
XFILL_1__12911_ vdd gnd FILL
XFILL_0__11552_ vdd gnd FILL
XFILL_1__13891_ vdd gnd FILL
XFILL_2__12112_ vdd gnd FILL
X_13747_ _13747_/A _13747_/B _13747_/C _13747_/Y vdd gnd OAI21X1
X_10959_ _10959_/A _10959_/B _10959_/C _10959_/Y vdd gnd OAI21X1
XFILL_0__10503_ vdd gnd FILL
XFILL_0__14271_ vdd gnd FILL
XFILL_1__12842_ vdd gnd FILL
XFILL_0__11483_ vdd gnd FILL
XFILL_2__12043_ vdd gnd FILL
X_13678_ _13678_/A _13678_/B _13678_/Y vdd gnd NAND2X1
XFILL_0__13222_ vdd gnd FILL
XFILL_2__8986_ vdd gnd FILL
XFILL_0__10434_ vdd gnd FILL
XFILL_1__12773_ vdd gnd FILL
X_12629_ _12629_/A _12629_/B _12629_/C _12629_/Y vdd gnd OAI21X1
XFILL_1__11724_ vdd gnd FILL
XFILL_0__13153_ vdd gnd FILL
XFILL_0__10365_ vdd gnd FILL
XFILL_0__9740_ vdd gnd FILL
XFILL_0__12104_ vdd gnd FILL
XFILL_2__7868_ vdd gnd FILL
XFILL_1__14443_ vdd gnd FILL
XFILL_0__13084_ vdd gnd FILL
XFILL_2__13994_ vdd gnd FILL
XFILL_0__10296_ vdd gnd FILL
X_7230_ _7230_/A _7230_/B _7230_/C _7230_/Y vdd gnd OAI21X1
XFILL_0__9671_ vdd gnd FILL
XFILL_1__10606_ vdd gnd FILL
XFILL_0__12035_ vdd gnd FILL
XFILL_1__14374_ vdd gnd FILL
XFILL_2__7799_ vdd gnd FILL
XFILL_1__11586_ vdd gnd FILL
XFILL_0__8622_ vdd gnd FILL
X_7161_ _7161_/A _7161_/B _7161_/S _7161_/Y vdd gnd MUX2X1
XFILL_1__10537_ vdd gnd FILL
XFILL_1__13325_ vdd gnd FILL
XFILL_2__12876_ vdd gnd FILL
XFILL_0__8553_ vdd gnd FILL
XFILL_2__14615_ vdd gnd FILL
X_7092_ _7092_/A _7092_/B _7092_/C _7092_/Y vdd gnd OAI21X1
XFILL_2__9469_ vdd gnd FILL
XFILL_1__13256_ vdd gnd FILL
XFILL_1__10468_ vdd gnd FILL
XFILL_0__7504_ vdd gnd FILL
XFILL_0__13986_ vdd gnd FILL
XFILL_0__8484_ vdd gnd FILL
XFILL_1__12207_ vdd gnd FILL
XFILL_1__13187_ vdd gnd FILL
XFILL_0__12937_ vdd gnd FILL
XFILL_1__10399_ vdd gnd FILL
XFILL_0__7435_ vdd gnd FILL
XFILL_1__12138_ vdd gnd FILL
XFILL_0__12868_ vdd gnd FILL
X_9802_ _9802_/D _9802_/CLK _9802_/Q vdd gnd DFFPOSX1
XFILL_0__7366_ vdd gnd FILL
X_7994_ _7994_/D _7994_/CLK _7994_/Q vdd gnd DFFPOSX1
XFILL_0__14607_ vdd gnd FILL
XFILL_0__11819_ vdd gnd FILL
XFILL_1__12069_ vdd gnd FILL
XFILL_0__9105_ vdd gnd FILL
XFILL_0__12799_ vdd gnd FILL
XFILL_0__7297_ vdd gnd FILL
X_9733_ _9733_/A _9733_/B _9733_/C _9733_/Y vdd gnd OAI21X1
XFILL_0__9036_ vdd gnd FILL
X_9664_ _9664_/A _9664_/B _9664_/C _9664_/D _9664_/Y vdd gnd OAI22X1
XFILL_0__14469_ vdd gnd FILL
X_8615_ _8615_/A _8615_/B _8615_/Y vdd gnd NAND2X1
X_9595_ _9595_/A _9595_/B _9595_/C _9595_/Y vdd gnd OAI21X1
XFILL_1__8800_ vdd gnd FILL
X_8546_ _8546_/A _8546_/Y vdd gnd INVX1
XFILL_0__9938_ vdd gnd FILL
XFILL_1__8731_ vdd gnd FILL
X_8477_ _8477_/A _8477_/B _8477_/Y vdd gnd NAND2X1
X_7428_ _7428_/A _7428_/Y vdd gnd INVX1
XFILL_0__9869_ vdd gnd FILL
XFILL_1__8662_ vdd gnd FILL
XFILL_1__7613_ vdd gnd FILL
X_7359_ _7359_/A _7359_/B _7359_/Y vdd gnd NOR2X1
XFILL_1__8593_ vdd gnd FILL
XFILL_1__7544_ vdd gnd FILL
X_9029_ _9029_/A _9029_/B _9029_/C _9029_/Y vdd gnd OAI21X1
XFILL_1__7475_ vdd gnd FILL
XFILL_1__9214_ vdd gnd FILL
X_12980_ _12980_/A _12980_/B _12980_/Y vdd gnd NAND2X1
X_11931_ _11931_/A _11931_/B _11931_/Y vdd gnd NAND2X1
XFILL_1__9145_ vdd gnd FILL
X_14650_ _14650_/A _14650_/B _14650_/Y vdd gnd NOR2X1
X_11862_ _11862_/A _11862_/B _11862_/Y vdd gnd NOR2X1
XFILL_1__9076_ vdd gnd FILL
X_13601_ _13601_/A _13601_/B _13601_/C _13601_/Y vdd gnd NAND3X1
X_10813_ _10813_/A _10813_/Y vdd gnd INVX1
X_14581_ _14581_/A _14581_/B _14581_/Y vdd gnd NAND2X1
XFILL_1__8027_ vdd gnd FILL
X_11793_ _11793_/A _11793_/B _11793_/Y vdd gnd NAND2X1
X_13532_ _13532_/A _13532_/B _13532_/Y vdd gnd NAND2X1
X_10744_ _10744_/D _10744_/CLK _10744_/Q vdd gnd DFFPOSX1
X_13463_ _13463_/D _13463_/CLK _13463_/Q vdd gnd DFFPOSX1
X_10675_ _10675_/A _10675_/B _10675_/C _10675_/Y vdd gnd OAI21X1
XFILL_1__9978_ vdd gnd FILL
X_12414_ _12414_/A _12414_/B _12414_/Y vdd gnd NAND2X1
XFILL_1__8929_ vdd gnd FILL
XFILL_2__7722_ vdd gnd FILL
X_13394_ _13394_/A _13394_/B _13394_/C _13394_/Y vdd gnd OAI21X1
XFILL_0__10150_ vdd gnd FILL
X_12345_ _12345_/A _12345_/B _12345_/Y vdd gnd NOR2X1
XFILL_2__7653_ vdd gnd FILL
XFILL_1__11440_ vdd gnd FILL
XFILL_2__10991_ vdd gnd FILL
XFILL_0__10081_ vdd gnd FILL
X_12276_ _12276_/A _12276_/B _12276_/C _12276_/Y vdd gnd AOI21X1
XFILL_2__7584_ vdd gnd FILL
XFILL_1__11371_ vdd gnd FILL
X_14015_ _14015_/A _14015_/B _14015_/Y vdd gnd NAND2X1
X_11227_ _11227_/A _11227_/B _11227_/C _11227_/Y vdd gnd OAI21X1
XFILL_1__13110_ vdd gnd FILL
XFILL_1__10322_ vdd gnd FILL
XFILL_1__14090_ vdd gnd FILL
XFILL_0__13840_ vdd gnd FILL
X_11158_ _11158_/A _11158_/B _11158_/C _11158_/Y vdd gnd OAI21X1
XFILL_1__13041_ vdd gnd FILL
XFILL_1__10253_ vdd gnd FILL
XFILL_0__13771_ vdd gnd FILL
XFILL_0__10983_ vdd gnd FILL
X_10109_ _10109_/A _10109_/B _10109_/Y vdd gnd NAND2X1
XFILL_2__8205_ vdd gnd FILL
X_11089_ _11089_/A _11089_/B _11089_/C _11089_/Y vdd gnd OAI21X1
XFILL_0__12722_ vdd gnd FILL
XFILL_1__10184_ vdd gnd FILL
XFILL_0__7220_ vdd gnd FILL
X_14917_ _14917_/A _14917_/Y vdd gnd BUFX2
XFILL_2__8136_ vdd gnd FILL
XFILL_0__12653_ vdd gnd FILL
XFILL_0__7151_ vdd gnd FILL
X_14848_ _14848_/A _14848_/B _14848_/C _14848_/Y vdd gnd OAI21X1
XFILL_2__10425_ vdd gnd FILL
XFILL_2__8067_ vdd gnd FILL
XFILL_0__11604_ vdd gnd FILL
XFILL_1__13943_ vdd gnd FILL
XFILL_0__7082_ vdd gnd FILL
X_14779_ _14779_/A _14779_/B _14779_/C _14779_/Y vdd gnd AOI21X1
XFILL_2__10356_ vdd gnd FILL
XFILL_0__14323_ vdd gnd FILL
XFILL_0__11535_ vdd gnd FILL
XFILL_1__13874_ vdd gnd FILL
XFILL_2__10287_ vdd gnd FILL
XFILL_0__14254_ vdd gnd FILL
XFILL_1__12825_ vdd gnd FILL
XFILL_0__11466_ vdd gnd FILL
X_8400_ _8400_/A _8400_/B _8400_/C _8400_/Y vdd gnd OAI21X1
X_9380_ _9380_/A _9380_/B _9380_/Y vdd gnd NAND2X1
XFILL_0__13205_ vdd gnd FILL
XFILL_2__8969_ vdd gnd FILL
XFILL_0__10417_ vdd gnd FILL
XFILL_0_BUFX2_insert360 vdd gnd FILL
XFILL_1__12756_ vdd gnd FILL
XFILL_0_BUFX2_insert371 vdd gnd FILL
X_8331_ _8331_/A _8331_/B _8331_/Y vdd gnd NAND2X1
XFILL_0__11397_ vdd gnd FILL
XFILL_0_BUFX2_insert382 vdd gnd FILL
XFILL_0__13136_ vdd gnd FILL
XFILL_1__11707_ vdd gnd FILL
XFILL_0__10348_ vdd gnd FILL
XFILL_0__9723_ vdd gnd FILL
XFILL_1__12687_ vdd gnd FILL
X_8262_ _8262_/A _8262_/B _8262_/C _8262_/Y vdd gnd NAND3X1
XFILL_1__14426_ vdd gnd FILL
XFILL_0__13067_ vdd gnd FILL
X_7213_ _7213_/A _7213_/B _7213_/C _7213_/D _7213_/Y vdd gnd OAI22X1
XFILL_0__10279_ vdd gnd FILL
XFILL_0__9654_ vdd gnd FILL
X_8193_ _8193_/A _8193_/B _8193_/Y vdd gnd NOR2X1
XFILL_0__12018_ vdd gnd FILL
XFILL_1__14357_ vdd gnd FILL
XFILL_1__11569_ vdd gnd FILL
XFILL_0__8605_ vdd gnd FILL
X_7144_ _7144_/A _7144_/Y vdd gnd INVX1
XFILL_0__9585_ vdd gnd FILL
XFILL_1__13308_ vdd gnd FILL
XFILL_1__14288_ vdd gnd FILL
XFILL_0__8536_ vdd gnd FILL
X_7075_ _7075_/A _7075_/Y vdd gnd INVX2
XFILL_1__13239_ vdd gnd FILL
XFILL_0__13969_ vdd gnd FILL
XFILL_1__7260_ vdd gnd FILL
XFILL_0__8467_ vdd gnd FILL
XFILL_0__7418_ vdd gnd FILL
XFILL_1__7191_ vdd gnd FILL
XFILL_0__8398_ vdd gnd FILL
XFILL_0__7349_ vdd gnd FILL
X_7977_ _7977_/D _7977_/CLK _7977_/Q vdd gnd DFFPOSX1
X_9716_ _9716_/A _9716_/Y vdd gnd INVX1
XFILL_1__9901_ vdd gnd FILL
XFILL_0__9019_ vdd gnd FILL
X_9647_ _9647_/A _9647_/B _9647_/C _9647_/Y vdd gnd AOI21X1
X_9578_ _9578_/A _9578_/B _9578_/Y vdd gnd NAND2X1
X_10460_ _10460_/A _10460_/B _10460_/Y vdd gnd NOR2X1
XFILL_1__9763_ vdd gnd FILL
X_8529_ _8529_/A _8529_/B _8529_/C _8529_/Y vdd gnd NAND3X1
X_10391_ _10391_/A _10391_/B _10391_/C _10391_/Y vdd gnd OAI21X1
XFILL_1__8714_ vdd gnd FILL
XFILL_1__9694_ vdd gnd FILL
X_12130_ _12130_/A _12130_/B _12130_/Y vdd gnd NAND2X1
XFILL_1__8645_ vdd gnd FILL
X_12061_ _12061_/A _12061_/B _12061_/C _12061_/D _12061_/Y vdd gnd AOI22X1
XFILL_1__8576_ vdd gnd FILL
X_11012_ _11012_/A _11012_/B _11012_/C _11012_/Y vdd gnd OAI21X1
XFILL_1__7527_ vdd gnd FILL
XFILL_1__7458_ vdd gnd FILL
X_12963_ _12963_/A _12963_/B _12963_/Y vdd gnd NAND2X1
XFILL_1__7389_ vdd gnd FILL
X_14702_ _14702_/A _14702_/Y vdd gnd INVX1
X_11914_ _11914_/A _11914_/B _11914_/Y vdd gnd NAND2X1
XFILL_1__9128_ vdd gnd FILL
X_12894_ _12894_/A _12894_/B _12894_/C _12894_/Y vdd gnd OAI21X1
X_14633_ _14633_/A _14633_/B _14633_/Y vdd gnd NAND2X1
XFILL_2__10210_ vdd gnd FILL
X_11845_ _11845_/A _11845_/Y vdd gnd INVX1
XFILL_1__9059_ vdd gnd FILL
XFILL_1__10940_ vdd gnd FILL
X_14564_ _14564_/A _14564_/B _14564_/Y vdd gnd NAND2X1
XFILL_2__10141_ vdd gnd FILL
X_11776_ _11776_/A _11776_/B _11776_/C _11776_/Y vdd gnd OAI21X1
XFILL_0__11320_ vdd gnd FILL
XFILL_1__10871_ vdd gnd FILL
X_13515_ _13515_/A _13515_/B _13515_/C _13515_/Y vdd gnd OAI21X1
X_10727_ _10727_/D _10727_/CLK _10727_/Q vdd gnd DFFPOSX1
X_14495_ _14495_/A _14495_/B _14495_/C _14495_/Y vdd gnd OAI21X1
XFILL_2__10072_ vdd gnd FILL
XFILL_0__11251_ vdd gnd FILL
XFILL_1__13590_ vdd gnd FILL
X_13446_ _13446_/D _13446_/CLK _13446_/Q vdd gnd DFFPOSX1
X_10658_ _10658_/A _10658_/B _10658_/Y vdd gnd NAND2X1
XFILL_0__10202_ vdd gnd FILL
XFILL_0__11182_ vdd gnd FILL
X_13377_ _13377_/A _13377_/B _13377_/C _13377_/Y vdd gnd OAI21X1
X_10589_ _10589_/A _10589_/B _10589_/Y vdd gnd NAND2X1
XFILL_0__10133_ vdd gnd FILL
XFILL_1__12472_ vdd gnd FILL
X_12328_ _12328_/A _12328_/Y vdd gnd INVX1
XFILL_1__11423_ vdd gnd FILL
XFILL_0__10064_ vdd gnd FILL
XFILL_2__10974_ vdd gnd FILL
X_12259_ _12259_/A _12259_/B _12259_/Y vdd gnd NAND2X1
XFILL_2__7567_ vdd gnd FILL
XFILL_1__11354_ vdd gnd FILL
XFILL_1__14142_ vdd gnd FILL
XFILL_1_BUFX2_insert16 vdd gnd FILL
XFILL_0__9370_ vdd gnd FILL
XFILL_1_BUFX2_insert27 vdd gnd FILL
XFILL_1__10305_ vdd gnd FILL
XFILL_1__14073_ vdd gnd FILL
XFILL_2__7498_ vdd gnd FILL
XFILL_1__11285_ vdd gnd FILL
XFILL_0__13823_ vdd gnd FILL
XFILL_0__8321_ vdd gnd FILL
XFILL_1__13024_ vdd gnd FILL
XFILL_1__10236_ vdd gnd FILL
XFILL_0__10966_ vdd gnd FILL
XFILL_0__13754_ vdd gnd FILL
X_7900_ _7900_/A _7900_/B _7900_/Y vdd gnd NAND2X1
XFILL_0__8252_ vdd gnd FILL
XFILL256350x75750 vdd gnd FILL
X_8880_ _8880_/D _8880_/CLK _8880_/Q vdd gnd DFFPOSX1
XFILL_1__10167_ vdd gnd FILL
XFILL_0__12705_ vdd gnd FILL
XFILL_0__7203_ vdd gnd FILL
XFILL_0__13685_ vdd gnd FILL
XFILL_0__10897_ vdd gnd FILL
X_7831_ _7831_/A _7831_/B _7831_/C _7831_/Y vdd gnd OAI21X1
XFILL_0__8183_ vdd gnd FILL
XFILL_2__8119_ vdd gnd FILL
XFILL_0__12636_ vdd gnd FILL
XFILL_1__10098_ vdd gnd FILL
XFILL_0__7134_ vdd gnd FILL
XFILL_2__10408_ vdd gnd FILL
X_7762_ _7762_/A _7762_/B _7762_/Y vdd gnd NAND2X1
XFILL_1__13926_ vdd gnd FILL
XFILL_1_CLKBUF1_insert39 vdd gnd FILL
X_9501_ _9501_/A _9501_/B _9501_/C _9501_/Y vdd gnd OAI21X1
XFILL_2__13127_ vdd gnd FILL
X_7693_ _7693_/A _7693_/B _7693_/Y vdd gnd NAND2X1
XFILL_2__10339_ vdd gnd FILL
XFILL_0__14306_ vdd gnd FILL
XFILL_0__11518_ vdd gnd FILL
XFILL_1__13857_ vdd gnd FILL
XFILL_0__12498_ vdd gnd FILL
X_9432_ _9432_/A _9432_/B _9432_/Y vdd gnd NAND2X1
XFILL_0__14237_ vdd gnd FILL
XFILL_1__12808_ vdd gnd FILL
XFILL_2__13058_ vdd gnd FILL
XFILL_0__11449_ vdd gnd FILL
XFILL_1__13788_ vdd gnd FILL
X_9363_ _9363_/A _9363_/B _9363_/Y vdd gnd NAND2X1
XFILL_0_BUFX2_insert190 vdd gnd FILL
XFILL_1__12739_ vdd gnd FILL
X_8314_ _8314_/A _8314_/B _8314_/Y vdd gnd AND2X2
X_9294_ _9294_/A _9294_/B _9294_/C _9294_/Y vdd gnd OAI21X1
XFILL_0__13119_ vdd gnd FILL
XFILL_0__9706_ vdd gnd FILL
XFILL_0__14099_ vdd gnd FILL
X_8245_ _8245_/A _8245_/Y vdd gnd INVX1
XFILL_0__7898_ vdd gnd FILL
XFILL_1__14409_ vdd gnd FILL
XFILL_0__9637_ vdd gnd FILL
XFILL_1__8430_ vdd gnd FILL
X_8176_ _8176_/A _8176_/Y vdd gnd INVX1
X_7127_ _7127_/A _7127_/B _7127_/C _7127_/Y vdd gnd OAI21X1
XFILL_0__9568_ vdd gnd FILL
XFILL_1__8361_ vdd gnd FILL
XFILL_1__7312_ vdd gnd FILL
XFILL_0__8519_ vdd gnd FILL
XFILL_0__9499_ vdd gnd FILL
XFILL_1__8292_ vdd gnd FILL
XFILL_1__7243_ vdd gnd FILL
XFILL_1__7174_ vdd gnd FILL
X_11630_ _11630_/D _11630_/CLK _11630_/Q vdd gnd DFFPOSX1
X_11561_ _11561_/A _11561_/B _11561_/C _11561_/Y vdd gnd OAI21X1
X_13300_ _13300_/A _13300_/Y vdd gnd INVX1
X_10512_ _10512_/A _10512_/B _10512_/C _10512_/Y vdd gnd OAI21X1
X_14280_ _14280_/A _14280_/Y vdd gnd INVX1
X_11492_ _11492_/A _11492_/Y vdd gnd INVX1
X_13231_ _13231_/A _13231_/B _13231_/Y vdd gnd AND2X2
X_10443_ _10443_/A _10443_/B _10443_/Y vdd gnd AND2X2
XFILL_1__9746_ vdd gnd FILL
X_13162_ _13162_/A _13162_/B _13162_/C _13162_/Y vdd gnd OAI21X1
X_10374_ _10374_/A _10374_/B _10374_/Y vdd gnd NOR2X1
XFILL_1__9677_ vdd gnd FILL
XFILL_2__8470_ vdd gnd FILL
X_12113_ _12113_/A _12113_/B _12113_/Y vdd gnd NAND2X1
XFILL_1__8628_ vdd gnd FILL
X_13093_ _13093_/A _13093_/B _13093_/Y vdd gnd NAND2X1
X_12044_ _12044_/A _12044_/Y vdd gnd INVX1
XFILL_1__8559_ vdd gnd FILL
XFILL_1__11070_ vdd gnd FILL
XFILL_0__10820_ vdd gnd FILL
XFILL_1__10021_ vdd gnd FILL
X_13995_ _13995_/A _13995_/B _13995_/Y vdd gnd NAND2X1
XFILL_2__12360_ vdd gnd FILL
XFILL_2_BUFX2_insert241 vdd gnd FILL
XFILL_2_BUFX2_insert263 vdd gnd FILL
X_12946_ _12946_/A _12946_/B _12946_/C _12946_/Y vdd gnd AOI21X1
XFILL_2_BUFX2_insert296 vdd gnd FILL
XFILL_2__12291_ vdd gnd FILL
XFILL_0__10682_ vdd gnd FILL
XFILL_2__14030_ vdd gnd FILL
X_12877_ _12877_/A _12877_/B _12877_/Y vdd gnd NAND2X1
XFILL_0__12421_ vdd gnd FILL
XFILL_1__14760_ vdd gnd FILL
X_14616_ _14616_/A _14616_/B _14616_/C _14616_/Y vdd gnd AOI21X1
XFILL_1__11972_ vdd gnd FILL
X_11828_ _11828_/A _11828_/B _11828_/C _11828_/Y vdd gnd AOI21X1
XFILL_2__9924_ vdd gnd FILL
XFILL_1__13711_ vdd gnd FILL
XFILL_0__12352_ vdd gnd FILL
XFILL_1__10923_ vdd gnd FILL
XFILL_1__14691_ vdd gnd FILL
X_14547_ _14547_/D _14547_/CLK _14547_/Q vdd gnd DFFPOSX1
X_11759_ _11759_/A _11759_/B _11759_/C _11759_/Y vdd gnd OAI21X1
XBUFX2_insert240 BUFX2_insert240/A BUFX2_insert240/Y vdd gnd BUFX2
XFILL_0__11303_ vdd gnd FILL
XFILL_1__13642_ vdd gnd FILL
XBUFX2_insert251 BUFX2_insert251/A BUFX2_insert251/Y vdd gnd BUFX2
XFILL_0__12283_ vdd gnd FILL
XFILL_1__10854_ vdd gnd FILL
XBUFX2_insert262 BUFX2_insert262/A BUFX2_insert262/Y vdd gnd BUFX2
XBUFX2_insert273 BUFX2_insert273/A BUFX2_insert273/Y vdd gnd BUFX2
XFILL_2__8806_ vdd gnd FILL
X_14478_ _14478_/A _14478_/B _14478_/C _14478_/Y vdd gnd OAI21X1
XBUFX2_insert284 BUFX2_insert284/A BUFX2_insert284/Y vdd gnd BUFX2
XFILL_0__14022_ vdd gnd FILL
XBUFX2_insert295 BUFX2_insert295/A BUFX2_insert295/Y vdd gnd BUFX2
XFILL_0__11234_ vdd gnd FILL
XFILL_1__10785_ vdd gnd FILL
XFILL_1__13573_ vdd gnd FILL
XFILL_0__7821_ vdd gnd FILL
X_13429_ _13429_/D _13429_/CLK _13429_/Q vdd gnd DFFPOSX1
XFILL_2__14863_ vdd gnd FILL
XFILL_1__12524_ vdd gnd FILL
XFILL_0__11165_ vdd gnd FILL
XFILL_0__7752_ vdd gnd FILL
XFILL_0__10116_ vdd gnd FILL
XFILL_2__14794_ vdd gnd FILL
XFILL_1__12455_ vdd gnd FILL
X_8030_ _8030_/A _8030_/B _8030_/C _8030_/Y vdd gnd OAI21X1
XFILL_0__11096_ vdd gnd FILL
XFILL_0__7683_ vdd gnd FILL
XFILL_1__11406_ vdd gnd FILL
XFILL_0__10047_ vdd gnd FILL
XFILL_1__12386_ vdd gnd FILL
XFILL_0__9422_ vdd gnd FILL
XFILL_1__11337_ vdd gnd FILL
XFILL_1__14125_ vdd gnd FILL
XFILL_0__14855_ vdd gnd FILL
XFILL_0__9353_ vdd gnd FILL
X_9981_ _9981_/A _9981_/B _9981_/S _9981_/Y vdd gnd MUX2X1
XFILL_1__11268_ vdd gnd FILL
XFILL_0__13806_ vdd gnd FILL
XFILL_1__14056_ vdd gnd FILL
XFILL_0__8304_ vdd gnd FILL
XFILL_0__14786_ vdd gnd FILL
XFILL_0__11998_ vdd gnd FILL
XFILL_0__9284_ vdd gnd FILL
X_8932_ _8932_/A _8932_/B _8932_/Y vdd gnd NOR2X1
XFILL_1__10219_ vdd gnd FILL
XFILL_1__13007_ vdd gnd FILL
XFILL_1__11199_ vdd gnd FILL
XFILL_0__13737_ vdd gnd FILL
XFILL_0__10949_ vdd gnd FILL
XFILL_0__8235_ vdd gnd FILL
X_8863_ _8863_/D _8863_/CLK _8863_/Q vdd gnd DFFPOSX1
XFILL_2__12489_ vdd gnd FILL
XFILL_0__13668_ vdd gnd FILL
X_7814_ _7814_/A _7814_/B _7814_/Y vdd gnd AND2X2
XFILL_0__8166_ vdd gnd FILL
XFILL_2__14228_ vdd gnd FILL
X_8794_ _8794_/A _8794_/B _8794_/C _8794_/Y vdd gnd OAI21X1
XFILL_0__12619_ vdd gnd FILL
XFILL_0__13599_ vdd gnd FILL
XFILL_0__7117_ vdd gnd FILL
X_7745_ _7745_/A _7745_/B _7745_/Y vdd gnd AND2X2
XFILL_0__8097_ vdd gnd FILL
XFILL_1__13909_ vdd gnd FILL
X_7676_ _7676_/A _7676_/Y vdd gnd INVX1
X_9415_ _9415_/A _9415_/B _9415_/Y vdd gnd NAND2X1
XFILL_1__7861_ vdd gnd FILL
XFILL_1__9600_ vdd gnd FILL
X_9346_ _9346_/A _9346_/B _9346_/C _9346_/Y vdd gnd AOI21X1
XFILL_0__8999_ vdd gnd FILL
XFILL_1__7792_ vdd gnd FILL
XFILL_1__9531_ vdd gnd FILL
X_9277_ _9277_/A _9277_/B _9277_/C _9277_/Y vdd gnd NOR3X1
XFILL256950x136950 vdd gnd FILL
XFILL_1__9462_ vdd gnd FILL
X_8228_ _8228_/A _8228_/B _8228_/C _8228_/Y vdd gnd OAI21X1
X_10090_ _10090_/A _10090_/B _10090_/C _10090_/Y vdd gnd AOI21X1
XFILL_1__8413_ vdd gnd FILL
XFILL_1__9393_ vdd gnd FILL
X_8159_ _8159_/A _8159_/Y vdd gnd INVX1
XFILL_1__8344_ vdd gnd FILL
XFILL_1__8275_ vdd gnd FILL
X_12800_ _12800_/A _12800_/B _12800_/C _12800_/Y vdd gnd OAI21X1
XFILL_1__7226_ vdd gnd FILL
X_13780_ _13780_/A _13780_/B _13780_/Y vdd gnd AND2X2
X_10992_ _10992_/A _10992_/B _10992_/C _10992_/Y vdd gnd OAI21X1
XFILL_1_BUFX2_insert204 vdd gnd FILL
XFILL_1_BUFX2_insert215 vdd gnd FILL
X_12731_ _12731_/A _12731_/B _12731_/S _12731_/Y vdd gnd MUX2X1
XFILL_1_BUFX2_insert226 vdd gnd FILL
XFILL_1__7157_ vdd gnd FILL
XFILL_1_BUFX2_insert237 vdd gnd FILL
XFILL_1_BUFX2_insert248 vdd gnd FILL
XFILL_1_BUFX2_insert259 vdd gnd FILL
X_12662_ _12662_/A _12662_/B _12662_/C _12662_/Y vdd gnd OAI21X1
XFILL_1__7088_ vdd gnd FILL
X_14401_ _14401_/A _14401_/B _14401_/Y vdd gnd OR2X2
X_11613_ _11613_/D _11613_/CLK _11613_/Q vdd gnd DFFPOSX1
X_12593_ _12593_/D _12593_/CLK _12593_/Q vdd gnd DFFPOSX1
X_14332_ _14332_/A _14332_/B _14332_/C _14332_/Y vdd gnd NAND3X1
XFILL_0_CLKBUF1_insert385 vdd gnd FILL
X_11544_ _11544_/A _11544_/B _11544_/C _11544_/Y vdd gnd OAI21X1
X_14263_ _14263_/A _14263_/Y vdd gnd INVX1
X_11475_ _11475_/A _11475_/B _11475_/Y vdd gnd NAND2X1
XFILL_1__10570_ vdd gnd FILL
X_13214_ _13214_/A _13214_/B _13214_/C _13214_/Y vdd gnd AOI21X1
X_10426_ _10426_/A _10426_/Y vdd gnd INVX1
XFILL_1__9729_ vdd gnd FILL
XFILL_2__8522_ vdd gnd FILL
X_14194_ _14194_/D _14194_/CLK _14194_/Q vdd gnd DFFPOSX1
XFILL_2__11860_ vdd gnd FILL
X_13145_ _13145_/A _13145_/B _13145_/Y vdd gnd NAND2X1
X_10357_ _10357_/A _10357_/B _10357_/C _10357_/Y vdd gnd AOI21X1
XFILL_2__8453_ vdd gnd FILL
XFILL_1__12240_ vdd gnd FILL
XFILL_2__11791_ vdd gnd FILL
XFILL_0__12970_ vdd gnd FILL
X_13076_ _13076_/A _13076_/B _13076_/Y vdd gnd OR2X2
X_10288_ _10288_/A _10288_/B _10288_/Y vdd gnd NAND2X1
XFILL_2__13530_ vdd gnd FILL
XFILL_2__8384_ vdd gnd FILL
XFILL_1__12171_ vdd gnd FILL
XFILL_0__11921_ vdd gnd FILL
X_12027_ _12027_/A _12027_/B _12027_/Y vdd gnd NAND2X1
XFILL_1__11122_ vdd gnd FILL
XFILL_0__14640_ vdd gnd FILL
XFILL_2__10673_ vdd gnd FILL
XFILL_0__11852_ vdd gnd FILL
XFILL_1__11053_ vdd gnd FILL
XFILL_0__10803_ vdd gnd FILL
XFILL_0__14571_ vdd gnd FILL
XFILL_0__11783_ vdd gnd FILL
XFILL_2__9005_ vdd gnd FILL
X_13978_ _13978_/A _13978_/B _13978_/C _13978_/Y vdd gnd AOI21X1
XFILL_1__10004_ vdd gnd FILL
XFILL_0__13522_ vdd gnd FILL
XFILL_0__8020_ vdd gnd FILL
X_12929_ _12929_/A _12929_/B _12929_/C _12929_/Y vdd gnd OAI21X1
XFILL_1__14812_ vdd gnd FILL
XFILL_0__10665_ vdd gnd FILL
XFILL256950x201750 vdd gnd FILL
XFILL_2__14013_ vdd gnd FILL
XFILL_2__11225_ vdd gnd FILL
XFILL_1__14743_ vdd gnd FILL
XFILL_0__12404_ vdd gnd FILL
XFILL_1__11955_ vdd gnd FILL
XFILL_0__13384_ vdd gnd FILL
XFILL_0__10596_ vdd gnd FILL
X_7530_ _7530_/A _7530_/B _7530_/Y vdd gnd NAND2X1
XFILL_0__9971_ vdd gnd FILL
XFILL_2__9907_ vdd gnd FILL
XFILL_0__12335_ vdd gnd FILL
XFILL_1__10906_ vdd gnd FILL
XFILL_1__14674_ vdd gnd FILL
XFILL_0__8922_ vdd gnd FILL
XFILL_1__11886_ vdd gnd FILL
X_7461_ _7461_/A _7461_/B _7461_/Y vdd gnd NAND2X1
XFILL_1__13625_ vdd gnd FILL
XFILL_0__12266_ vdd gnd FILL
XFILL_1__10837_ vdd gnd FILL
X_9200_ _9200_/A _9200_/B _9200_/C _9200_/Y vdd gnd OAI21X1
X_7392_ _7392_/A _7392_/B _7392_/C _7392_/Y vdd gnd OAI21X1
XFILL_0__14005_ vdd gnd FILL
XFILL_0__11217_ vdd gnd FILL
XFILL_1__13556_ vdd gnd FILL
XFILL_0__7804_ vdd gnd FILL
XFILL_1__10768_ vdd gnd FILL
XFILL_0__12197_ vdd gnd FILL
X_9131_ _9131_/A _9131_/Y vdd gnd INVX1
XFILL_0__8784_ vdd gnd FILL
XFILL_2__14846_ vdd gnd FILL
XFILL_1__12507_ vdd gnd FILL
XFILL_0__11148_ vdd gnd FILL
X_9062_ _9062_/A _9062_/B _9062_/C _9062_/Y vdd gnd AOI21X1
XFILL_0__7735_ vdd gnd FILL
XFILL_2__14777_ vdd gnd FILL
XFILL_1__12438_ vdd gnd FILL
XFILL_0__11079_ vdd gnd FILL
XFILL_2__11989_ vdd gnd FILL
X_8013_ _8013_/A _8013_/B _8013_/C _8013_/Y vdd gnd AOI21X1
XFILL_0__7666_ vdd gnd FILL
XFILL_0__9405_ vdd gnd FILL
XFILL_1__12369_ vdd gnd FILL
XFILL_0__7597_ vdd gnd FILL
XFILL_1__14108_ vdd gnd FILL
XFILL_0__14838_ vdd gnd FILL
XFILL_0__9336_ vdd gnd FILL
X_9964_ _9964_/A _9964_/B _9964_/S _9964_/Y vdd gnd MUX2X1
XFILL_1__14039_ vdd gnd FILL
XFILL_0__14769_ vdd gnd FILL
XFILL_0__9267_ vdd gnd FILL
X_8915_ _8915_/D _8915_/CLK _8915_/Q vdd gnd DFFPOSX1
XFILL_1__8060_ vdd gnd FILL
X_9895_ _9895_/A _9895_/Y vdd gnd INVX1
XFILL_0__8218_ vdd gnd FILL
XFILL_0__9198_ vdd gnd FILL
X_8846_ _8846_/D _8846_/CLK _8846_/Q vdd gnd DFFPOSX1
XFILL256950x111750 vdd gnd FILL
XFILL_0__8149_ vdd gnd FILL
X_8777_ _8777_/A _8777_/B _8777_/C _8777_/Y vdd gnd OAI21X1
XFILL_1__8962_ vdd gnd FILL
X_7728_ _7728_/A _7728_/B _7728_/C _7728_/Y vdd gnd OAI21X1
XFILL_1__7913_ vdd gnd FILL
X_7659_ _7659_/A _7659_/B _7659_/C _7659_/Y vdd gnd OAI21X1
XFILL_1__7844_ vdd gnd FILL
X_11260_ _11260_/A _11260_/B _11260_/C _11260_/Y vdd gnd AOI21X1
X_9329_ _9329_/A _9329_/B _9329_/Y vdd gnd NAND2X1
XFILL_1__7775_ vdd gnd FILL
X_10211_ _10211_/A _10211_/B _10211_/Y vdd gnd NOR2X1
XFILL_1__9514_ vdd gnd FILL
X_11191_ _11191_/A _11191_/B _11191_/C _11191_/Y vdd gnd AOI21X1
XFILL257250x10950 vdd gnd FILL
X_10142_ _10142_/A _10142_/B _10142_/C _10142_/D _10142_/Y vdd gnd AOI22X1
XFILL_1__9445_ vdd gnd FILL
X_10073_ _10073_/A _10073_/B _10073_/C _10073_/Y vdd gnd NAND3X1
XFILL_1__9376_ vdd gnd FILL
X_13901_ _13901_/A _13901_/B _13901_/Y vdd gnd NAND2X1
X_14881_ _14881_/D _14881_/CLK _14881_/Q vdd gnd DFFPOSX1
XFILL_1__8327_ vdd gnd FILL
X_13832_ _13832_/A _13832_/B _13832_/Y vdd gnd NAND2X1
XFILL_1__8258_ vdd gnd FILL
XFILL_1__7209_ vdd gnd FILL
X_13763_ _13763_/A _13763_/B _13763_/C _13763_/Y vdd gnd OAI21X1
X_10975_ _10975_/A _10975_/B _10975_/C _10975_/Y vdd gnd OAI21X1
XFILL_1__8189_ vdd gnd FILL
X_12714_ _12714_/A _12714_/B _12714_/C _12714_/Y vdd gnd OAI21X1
X_13694_ _13694_/A _13694_/Y vdd gnd INVX1
XFILL_0__10450_ vdd gnd FILL
X_12645_ _12645_/A _12645_/Y vdd gnd INVX1
XFILL_2__11010_ vdd gnd FILL
XFILL_1__11740_ vdd gnd FILL
XFILL_0__10381_ vdd gnd FILL
X_12576_ _12576_/D _12576_/CLK _12576_/Q vdd gnd DFFPOSX1
XFILL_0__12120_ vdd gnd FILL
XFILL_2__7884_ vdd gnd FILL
X_14315_ _14315_/A _14315_/B _14315_/Y vdd gnd NAND2X1
X_11527_ _11527_/A _11527_/B _11527_/C _11527_/Y vdd gnd OAI21X1
XFILL_1__13410_ vdd gnd FILL
XFILL_1__10622_ vdd gnd FILL
XFILL_0__12051_ vdd gnd FILL
XFILL_1__14390_ vdd gnd FILL
X_14246_ _14246_/A _14246_/Y vdd gnd INVX1
X_11458_ _11458_/A _11458_/B _11458_/Y vdd gnd NAND2X1
XFILL_0__11002_ vdd gnd FILL
XFILL_2__11912_ vdd gnd FILL
XFILL_1__13341_ vdd gnd FILL
XFILL_1__10553_ vdd gnd FILL
X_10409_ _10409_/A _10409_/B _10409_/C _10409_/Y vdd gnd OAI21X1
XFILL_2__8505_ vdd gnd FILL
X_14177_ _14177_/D _14177_/CLK _14177_/Q vdd gnd DFFPOSX1
XFILL_2__14631_ vdd gnd FILL
X_11389_ _11389_/A _11389_/B _11389_/Y vdd gnd NAND2X1
XFILL_2__11843_ vdd gnd FILL
XFILL_1__10484_ vdd gnd FILL
XFILL_1__13272_ vdd gnd FILL
X_13128_ _13128_/A _13128_/B _13128_/Y vdd gnd AND2X2
XFILL_0__7520_ vdd gnd FILL
XFILL_2__8436_ vdd gnd FILL
XFILL_2__14562_ vdd gnd FILL
XFILL_1__12223_ vdd gnd FILL
XFILL_2__11774_ vdd gnd FILL
XFILL_0__12953_ vdd gnd FILL
XFILL_0__7451_ vdd gnd FILL
X_13059_ _13059_/A _13059_/Y vdd gnd INVX1
XFILL_2__13513_ vdd gnd FILL
XFILL_2__8367_ vdd gnd FILL
XFILL_0__11904_ vdd gnd FILL
XFILL_1__12154_ vdd gnd FILL
XFILL_0__12884_ vdd gnd FILL
XFILL_0__7382_ vdd gnd FILL
XFILL_1__11105_ vdd gnd FILL
XFILL_0__14623_ vdd gnd FILL
XFILL_2__10656_ vdd gnd FILL
XFILL_1__12085_ vdd gnd FILL
XFILL_2__8298_ vdd gnd FILL
XFILL_0__9121_ vdd gnd FILL
XFILL_0__11835_ vdd gnd FILL
XFILL_1__11036_ vdd gnd FILL
XFILL_2__10587_ vdd gnd FILL
XFILL_0__9052_ vdd gnd FILL
X_8700_ _8700_/A _8700_/Y vdd gnd INVX1
XFILL_0__11766_ vdd gnd FILL
X_9680_ _9680_/A _9680_/B _9680_/Y vdd gnd NAND2X1
XFILL_0__13505_ vdd gnd FILL
XFILL_0__8003_ vdd gnd FILL
XFILL_0__11697_ vdd gnd FILL
XFILL_0__14485_ vdd gnd FILL
X_8631_ _8631_/A _8631_/B _8631_/C _8631_/Y vdd gnd OAI21X1
XFILL_0__10648_ vdd gnd FILL
XFILL_1__12987_ vdd gnd FILL
XFILL_2__11208_ vdd gnd FILL
X_8562_ _8562_/A _8562_/B _8562_/C _8562_/D _8562_/Y vdd gnd OAI22X1
XFILL_1__14726_ vdd gnd FILL
XFILL_1__11938_ vdd gnd FILL
XFILL_0__10579_ vdd gnd FILL
XFILL_0__13367_ vdd gnd FILL
X_7513_ _7513_/A _7513_/B _7513_/Y vdd gnd NOR2X1
XFILL_0__9954_ vdd gnd FILL
XFILL_2__11139_ vdd gnd FILL
X_8493_ _8493_/A _8493_/B _8493_/Y vdd gnd AND2X2
XFILL_1__14657_ vdd gnd FILL
XFILL_0__12318_ vdd gnd FILL
XFILL_1__11869_ vdd gnd FILL
XFILL_0__13298_ vdd gnd FILL
X_7444_ _7444_/A _7444_/B _7444_/C _7444_/Y vdd gnd OAI21X1
XFILL_0__9885_ vdd gnd FILL
XFILL_1__13608_ vdd gnd FILL
XFILL_0__12249_ vdd gnd FILL
XFILL_1__14588_ vdd gnd FILL
XFILL_0__8836_ vdd gnd FILL
X_7375_ _7375_/A _7375_/B _7375_/C _7375_/Y vdd gnd OAI21X1
XFILL_1__13539_ vdd gnd FILL
X_9114_ _9114_/A _9114_/Y vdd gnd INVX2
XFILL_1__7560_ vdd gnd FILL
XFILL_0__8767_ vdd gnd FILL
XFILL_2_CLKBUF1_insert91 vdd gnd FILL
XFILL_2__14829_ vdd gnd FILL
XFILL_0__7718_ vdd gnd FILL
X_9045_ _9045_/A _9045_/Y vdd gnd INVX1
XFILL_1__7491_ vdd gnd FILL
XFILL_0__8698_ vdd gnd FILL
XFILL_1__9230_ vdd gnd FILL
XFILL_0__7649_ vdd gnd FILL
XFILL_1__9161_ vdd gnd FILL
XFILL_0__9319_ vdd gnd FILL
XFILL_1__8112_ vdd gnd FILL
X_9947_ _9947_/A _9947_/Y vdd gnd INVX1
XFILL_1__9092_ vdd gnd FILL
XFILL_1__8043_ vdd gnd FILL
X_9878_ _9878_/A _9878_/B _9878_/C _9878_/Y vdd gnd OAI21X1
X_10760_ _10760_/D _10760_/CLK _10760_/Q vdd gnd DFFPOSX1
X_8829_ _8829_/A _8829_/B _8829_/C _8829_/Y vdd gnd OAI21X1
X_10691_ _10691_/D _10691_/CLK _10691_/Q vdd gnd DFFPOSX1
XFILL_1__9994_ vdd gnd FILL
X_12430_ _12430_/A _12430_/B _12430_/C _12430_/Y vdd gnd AOI21X1
XFILL_1__8945_ vdd gnd FILL
X_12361_ _12361_/A _12361_/B _12361_/Y vdd gnd OR2X2
X_14100_ _14100_/A _14100_/B _14100_/Y vdd gnd NAND2X1
X_11312_ _11312_/A _11312_/Y vdd gnd INVX1
XFILL_1__7827_ vdd gnd FILL
X_12292_ _12292_/A _12292_/B _12292_/Y vdd gnd NOR2X1
X_14031_ _14031_/A _14031_/B _14031_/C _14031_/Y vdd gnd AOI21X1
X_11243_ _11243_/A _11243_/B _11243_/Y vdd gnd OR2X2
XFILL_1__7758_ vdd gnd FILL
X_11174_ _11174_/A _11174_/Y vdd gnd INVX1
XFILL_1__7689_ vdd gnd FILL
X_10125_ _10125_/A _10125_/B _10125_/Y vdd gnd NOR2X1
XFILL_1__9428_ vdd gnd FILL
X_10056_ _10056_/A _10056_/B _10056_/C _10056_/Y vdd gnd AOI21X1
XFILL_1__9359_ vdd gnd FILL
XFILL_2__7103_ vdd gnd FILL
X_14864_ _14864_/A _14864_/B _14864_/C _14864_/Y vdd gnd OAI21X1
X_13815_ _13815_/A _13815_/B _13815_/C _13815_/Y vdd gnd OAI21X1
X_14795_ _14795_/A _14795_/B _14795_/Y vdd gnd NOR2X1
XFILL_2__13160_ vdd gnd FILL
XFILL_1__12910_ vdd gnd FILL
XFILL_2__10372_ vdd gnd FILL
XFILL_0__11551_ vdd gnd FILL
XFILL_1__13890_ vdd gnd FILL
X_13746_ _13746_/A _13746_/Y vdd gnd INVX1
X_10958_ _10958_/A _10958_/B _10958_/Y vdd gnd NAND2X1
XFILL_0__10502_ vdd gnd FILL
XFILL_1__12841_ vdd gnd FILL
XFILL_2__13091_ vdd gnd FILL
XFILL_0__14270_ vdd gnd FILL
XFILL_0__11482_ vdd gnd FILL
X_13677_ _13677_/A _13677_/B _13677_/C _13677_/Y vdd gnd OAI21X1
X_10889_ _10889_/A _10889_/B _10889_/S _10889_/Y vdd gnd MUX2X1
XFILL_0__10433_ vdd gnd FILL
XFILL_0__13221_ vdd gnd FILL
XFILL_1__12772_ vdd gnd FILL
X_12628_ _12628_/A _12628_/B _12628_/Y vdd gnd NAND2X1
XFILL_0__13152_ vdd gnd FILL
XFILL_1__11723_ vdd gnd FILL
XFILL_0__10364_ vdd gnd FILL
X_12559_ _12559_/D _12559_/CLK _12559_/Q vdd gnd DFFPOSX1
XFILL_0__12103_ vdd gnd FILL
XFILL_1__14442_ vdd gnd FILL
XFILL_0__13083_ vdd gnd FILL
XFILL_0__10295_ vdd gnd FILL
XFILL_0__9670_ vdd gnd FILL
XFILL_1__10605_ vdd gnd FILL
XFILL_0__12034_ vdd gnd FILL
XFILL_1__14373_ vdd gnd FILL
X_14229_ _14229_/A _14229_/B _14229_/Y vdd gnd NAND2X1
XFILL_0__8621_ vdd gnd FILL
XFILL_1__11585_ vdd gnd FILL
X_7160_ _7160_/A _7160_/B _7160_/S _7160_/Y vdd gnd MUX2X1
XFILL_1__13324_ vdd gnd FILL
XFILL_1__10536_ vdd gnd FILL
XFILL_0__8552_ vdd gnd FILL
X_7091_ _7091_/A _7091_/B _7091_/Y vdd gnd NAND2X1
XFILL_2__11826_ vdd gnd FILL
XFILL_1__13255_ vdd gnd FILL
XFILL_0__7503_ vdd gnd FILL
XFILL_1__10467_ vdd gnd FILL
XFILL_0__13985_ vdd gnd FILL
XFILL_0__8483_ vdd gnd FILL
XFILL_1__12206_ vdd gnd FILL
XFILL_2__11757_ vdd gnd FILL
XFILL_1__13186_ vdd gnd FILL
XFILL_0__12936_ vdd gnd FILL
XFILL_1__10398_ vdd gnd FILL
XFILL_0__7434_ vdd gnd FILL
XFILL_1__12137_ vdd gnd FILL
X_9801_ _9801_/D _9801_/CLK _9801_/Q vdd gnd DFFPOSX1
XFILL_0__12867_ vdd gnd FILL
XFILL_0__7365_ vdd gnd FILL
XFILL_2__13427_ vdd gnd FILL
XFILL_2__10639_ vdd gnd FILL
XFILL_0__14606_ vdd gnd FILL
X_7993_ _7993_/D _7993_/CLK _7993_/Q vdd gnd DFFPOSX1
XFILL_0__9104_ vdd gnd FILL
XFILL_0__11818_ vdd gnd FILL
XFILL_1__12068_ vdd gnd FILL
X_9732_ _9732_/A _9732_/B _9732_/C _9732_/Y vdd gnd OAI21X1
XFILL_0__12798_ vdd gnd FILL
XFILL_0__7296_ vdd gnd FILL
XFILL_1__11019_ vdd gnd FILL
XFILL_2__13358_ vdd gnd FILL
XFILL_0__9035_ vdd gnd FILL
XFILL_0__11749_ vdd gnd FILL
X_9663_ _9663_/A _9663_/B _9663_/C _9663_/Y vdd gnd OAI21X1
XFILL_2__13289_ vdd gnd FILL
XFILL_0__14468_ vdd gnd FILL
X_8614_ _8614_/A _8614_/B _8614_/Y vdd gnd NAND2X1
X_9594_ _9594_/A _9594_/B _9594_/C _9594_/Y vdd gnd OAI21X1
XFILL_0__13419_ vdd gnd FILL
XFILL_0__14399_ vdd gnd FILL
X_8545_ _8545_/A _8545_/B _8545_/C _8545_/Y vdd gnd AOI21X1
XFILL_1__14709_ vdd gnd FILL
XFILL_1__8730_ vdd gnd FILL
XFILL_0__9937_ vdd gnd FILL
X_8476_ _8476_/A _8476_/B _8476_/C _8476_/Y vdd gnd OAI21X1
X_7427_ _7427_/A _7427_/B _7427_/Y vdd gnd NAND2X1
XFILL_1__8661_ vdd gnd FILL
XFILL_0__9868_ vdd gnd FILL
XFILL_1__7612_ vdd gnd FILL
XFILL_0__8819_ vdd gnd FILL
X_7358_ _7358_/A _7358_/B _7358_/C _7358_/Y vdd gnd NAND3X1
XFILL_1__8592_ vdd gnd FILL
XFILL_1__7543_ vdd gnd FILL
X_7289_ _7289_/A _7289_/Y vdd gnd INVX1
X_9028_ _9028_/A _9028_/B _9028_/Y vdd gnd NAND2X1
XFILL_1__7474_ vdd gnd FILL
XFILL_1__9213_ vdd gnd FILL
X_11930_ _11930_/A _11930_/B _11930_/C _11930_/Y vdd gnd NAND3X1
XFILL_1__9144_ vdd gnd FILL
X_11861_ _11861_/A _11861_/B _11861_/C _11861_/Y vdd gnd OAI21X1
XFILL_1__9075_ vdd gnd FILL
X_13600_ _13600_/A _13600_/B _13600_/S _13600_/Y vdd gnd MUX2X1
X_10812_ _10812_/A _10812_/B _10812_/C _10812_/Y vdd gnd AOI21X1
X_14580_ _14580_/A _14580_/Y vdd gnd INVX1
XFILL_1__8026_ vdd gnd FILL
X_11792_ _11792_/A _11792_/Y vdd gnd INVX1
XFILL257550x36150 vdd gnd FILL
X_13531_ _13531_/A _13531_/Y vdd gnd INVX1
X_10743_ _10743_/D _10743_/CLK _10743_/Q vdd gnd DFFPOSX1
X_13462_ _13462_/D _13462_/CLK _13462_/Q vdd gnd DFFPOSX1
X_10674_ _10674_/A _10674_/B _10674_/Y vdd gnd NAND2X1
XFILL_2__8770_ vdd gnd FILL
XFILL_1__9977_ vdd gnd FILL
X_12413_ _12413_/A _12413_/B _12413_/C _12413_/D _12413_/Y vdd gnd AOI22X1
X_13393_ _13393_/A _13393_/B _13393_/C _13393_/Y vdd gnd OAI21X1
XFILL_1__8928_ vdd gnd FILL
X_12344_ _12344_/A _12344_/Y vdd gnd INVX1
XFILL_0__10080_ vdd gnd FILL
X_12275_ _12275_/A _12275_/Y vdd gnd INVX1
XFILL_1__11370_ vdd gnd FILL
X_14014_ _14014_/A _14014_/Y vdd gnd INVX1
X_11226_ _11226_/A _11226_/B _11226_/Y vdd gnd NAND2X1
XFILL_2__9322_ vdd gnd FILL
XFILL_1__10321_ vdd gnd FILL
XFILL_2__12660_ vdd gnd FILL
X_11157_ _11157_/A _11157_/B _11157_/Y vdd gnd NAND2X1
XFILL_2__9253_ vdd gnd FILL
XFILL_2__11611_ vdd gnd FILL
XFILL_1__10252_ vdd gnd FILL
XFILL_1__13040_ vdd gnd FILL
X_10108_ _10108_/A _10108_/B _10108_/C _10108_/Y vdd gnd OAI21X1
XFILL_0__13770_ vdd gnd FILL
XFILL_0__10982_ vdd gnd FILL
X_11088_ _11088_/A _11088_/B _11088_/C _11088_/Y vdd gnd OAI21X1
XFILL_2__14330_ vdd gnd FILL
XFILL_2__11542_ vdd gnd FILL
XFILL_0__12721_ vdd gnd FILL
XFILL_1__10183_ vdd gnd FILL
X_10039_ _10039_/A _10039_/B _10039_/C _10039_/Y vdd gnd OAI21X1
X_14916_ _14916_/A _14916_/Y vdd gnd BUFX2
XFILL_2__14261_ vdd gnd FILL
XFILL_0__12652_ vdd gnd FILL
XFILL_0__7150_ vdd gnd FILL
XFILL_2__13212_ vdd gnd FILL
X_14847_ _14847_/A _14847_/B _14847_/Y vdd gnd NOR2X1
XFILL_0__11603_ vdd gnd FILL
XFILL_1__13942_ vdd gnd FILL
XFILL_0__7081_ vdd gnd FILL
XFILL_2__13143_ vdd gnd FILL
X_14778_ _14778_/A _14778_/B _14778_/Y vdd gnd NAND2X1
XFILL_0__14322_ vdd gnd FILL
XFILL_1__13873_ vdd gnd FILL
XFILL_0__11534_ vdd gnd FILL
X_13729_ _13729_/A _13729_/B _13729_/Y vdd gnd NOR2X1
XFILL_1__12824_ vdd gnd FILL
XFILL_2__13074_ vdd gnd FILL
XFILL_0__14253_ vdd gnd FILL
XFILL_0__11465_ vdd gnd FILL
XFILL_0__13204_ vdd gnd FILL
XFILL_0_BUFX2_insert350 vdd gnd FILL
XFILL_0__10416_ vdd gnd FILL
XFILL_1__12755_ vdd gnd FILL
XFILL_0_BUFX2_insert361 vdd gnd FILL
XFILL_0__11396_ vdd gnd FILL
X_8330_ _8330_/A _8330_/B _8330_/C _8330_/Y vdd gnd NAND3X1
XFILL_0_BUFX2_insert372 vdd gnd FILL
XFILL_1__11706_ vdd gnd FILL
XFILL_0_BUFX2_insert383 vdd gnd FILL
XFILL_0__13135_ vdd gnd FILL
XFILL_0__10347_ vdd gnd FILL
XFILL_1__12686_ vdd gnd FILL
XFILL_0__9722_ vdd gnd FILL
X_8261_ _8261_/A _8261_/B _8261_/Y vdd gnd NAND2X1
XFILL_1__14425_ vdd gnd FILL
XFILL_0__13066_ vdd gnd FILL
XFILL_0__10278_ vdd gnd FILL
X_7212_ _7212_/A _7212_/B _7212_/Y vdd gnd NAND2X1
XFILL_0__9653_ vdd gnd FILL
X_8192_ _8192_/A _8192_/B _8192_/Y vdd gnd OR2X2
XFILL_0__12017_ vdd gnd FILL
XFILL_1__14356_ vdd gnd FILL
XFILL_0__8604_ vdd gnd FILL
XFILL_1__11568_ vdd gnd FILL
X_7143_ _7143_/A _7143_/B _7143_/C _7143_/Y vdd gnd OAI21X1
XFILL_0__9584_ vdd gnd FILL
XFILL_1__13307_ vdd gnd FILL
XFILL_1__10519_ vdd gnd FILL
XFILL_1__14287_ vdd gnd FILL
XFILL_0__8535_ vdd gnd FILL
XFILL_1__11499_ vdd gnd FILL
X_7074_ _7074_/A _7074_/B _7074_/Y vdd gnd NOR2X1
XFILL_1__13238_ vdd gnd FILL
XFILL_0__13968_ vdd gnd FILL
XFILL_0__8466_ vdd gnd FILL
XFILL_1__13169_ vdd gnd FILL
XFILL_0__12919_ vdd gnd FILL
XFILL_0__7417_ vdd gnd FILL
XFILL_0__13899_ vdd gnd FILL
XFILL_1__7190_ vdd gnd FILL
XFILL_0__8397_ vdd gnd FILL
XFILL_2__14459_ vdd gnd FILL
XFILL_0__7348_ vdd gnd FILL
X_7976_ _7976_/D _7976_/CLK _7976_/Q vdd gnd DFFPOSX1
X_9715_ _9715_/A _9715_/B _9715_/C _9715_/Y vdd gnd OAI21X1
XFILL_0__7279_ vdd gnd FILL
XFILL_0__9018_ vdd gnd FILL
XFILL_1__9900_ vdd gnd FILL
X_9646_ _9646_/A _9646_/Y vdd gnd INVX1
X_9577_ _9577_/A _9577_/B _9577_/Y vdd gnd NOR2X1
X_8528_ _8528_/A _8528_/B _8528_/C _8528_/Y vdd gnd OAI21X1
XFILL_1__9762_ vdd gnd FILL
X_10390_ _10390_/A _10390_/B _10390_/C _10390_/D _10390_/Y vdd gnd AOI22X1
XFILL_1__8713_ vdd gnd FILL
XFILL_1__9693_ vdd gnd FILL
X_8459_ _8459_/A _8459_/B _8459_/C _8459_/Y vdd gnd OAI21X1
XFILL_1__8644_ vdd gnd FILL
X_12060_ _12060_/A _12060_/B _12060_/Y vdd gnd NOR2X1
XFILL_2_CLKBUF1_insert103 vdd gnd FILL
XFILL_1__8575_ vdd gnd FILL
X_11011_ _11011_/A _11011_/B _11011_/Y vdd gnd NOR2X1
XFILL_1__7526_ vdd gnd FILL
XFILL_1__7457_ vdd gnd FILL
X_12962_ _12962_/A _12962_/B _12962_/Y vdd gnd NAND2X1
XFILL_1__7388_ vdd gnd FILL
X_14701_ _14701_/A _14701_/B _14701_/Y vdd gnd NAND2X1
X_11913_ _11913_/A _11913_/Y vdd gnd INVX1
XFILL_1__9127_ vdd gnd FILL
X_12893_ _12893_/A _12893_/B _12893_/Y vdd gnd OR2X2
X_14632_ _14632_/A _14632_/B _14632_/C _14632_/Y vdd gnd OAI21X1
X_11844_ _11844_/A _11844_/B _11844_/Y vdd gnd NOR2X1
XFILL_1__9058_ vdd gnd FILL
XFILL_2__9940_ vdd gnd FILL
X_14563_ _14563_/A _14563_/B _14563_/C _14563_/Y vdd gnd OAI21X1
XFILL_1__8009_ vdd gnd FILL
X_11775_ _11775_/A _11775_/B _11775_/C _11775_/Y vdd gnd OAI21X1
XFILL_2__9871_ vdd gnd FILL
XFILL_1__10870_ vdd gnd FILL
X_10726_ _10726_/D _10726_/CLK _10726_/Q vdd gnd DFFPOSX1
X_13514_ _13514_/A _13514_/B _13514_/Y vdd gnd NAND2X1
X_14494_ _14494_/A _14494_/B _14494_/Y vdd gnd NAND2X1
XFILL_2__8822_ vdd gnd FILL
XFILL_0__11250_ vdd gnd FILL
X_13445_ _13445_/D _13445_/CLK _13445_/Q vdd gnd DFFPOSX1
X_10657_ _10657_/A _10657_/B _10657_/C _10657_/Y vdd gnd OAI21X1
XFILL_0__10201_ vdd gnd FILL
XFILL_2__8753_ vdd gnd FILL
XFILL_0__11181_ vdd gnd FILL
X_13376_ _13376_/A _13376_/B _13376_/Y vdd gnd NAND2X1
X_10588_ _10588_/A _10588_/B _10588_/C _10588_/D _10588_/Y vdd gnd OAI22X1
XFILL_2__13830_ vdd gnd FILL
XFILL_0__10132_ vdd gnd FILL
XFILL_2__8684_ vdd gnd FILL
XFILL_1__12471_ vdd gnd FILL
X_12327_ _12327_/A _12327_/B _12327_/C _12327_/Y vdd gnd OAI21X1
XFILL_1__11422_ vdd gnd FILL
XFILL_2__13761_ vdd gnd FILL
XFILL_0__10063_ vdd gnd FILL
X_12258_ _12258_/A _12258_/B _12258_/C _12258_/D _12258_/Y vdd gnd OAI22X1
XFILL_2__12712_ vdd gnd FILL
XFILL_1__14141_ vdd gnd FILL
XFILL_2__13692_ vdd gnd FILL
XFILL_1__11353_ vdd gnd FILL
X_11209_ _11209_/A _11209_/B _11209_/Y vdd gnd NOR2X1
XFILL_2__9305_ vdd gnd FILL
XFILL_1_BUFX2_insert17 vdd gnd FILL
X_12189_ _12189_/A _12189_/B _12189_/Y vdd gnd AND2X2
XFILL_2__12643_ vdd gnd FILL
XFILL_1__10304_ vdd gnd FILL
XFILL_1_BUFX2_insert28 vdd gnd FILL
XFILL_1__14072_ vdd gnd FILL
XFILL_0__13822_ vdd gnd FILL
XFILL_0__8320_ vdd gnd FILL
XFILL_1__11284_ vdd gnd FILL
XFILL_2__9236_ vdd gnd FILL
XFILL_1__13023_ vdd gnd FILL
XFILL_1__10235_ vdd gnd FILL
XFILL_0__13753_ vdd gnd FILL
XFILL_0__10965_ vdd gnd FILL
XFILL_0__8251_ vdd gnd FILL
XFILL_2__14313_ vdd gnd FILL
XFILL_2__9167_ vdd gnd FILL
XFILL_2__11525_ vdd gnd FILL
XFILL_0__12704_ vdd gnd FILL
XFILL_0__7202_ vdd gnd FILL
XFILL_1__10166_ vdd gnd FILL
XFILL_0__13684_ vdd gnd FILL
X_7830_ _7830_/A _7830_/B _7830_/C _7830_/Y vdd gnd OAI21X1
XFILL_0__8182_ vdd gnd FILL
XFILL_0__10896_ vdd gnd FILL
XFILL_2__14244_ vdd gnd FILL
XFILL_2__9098_ vdd gnd FILL
XFILL_2__11456_ vdd gnd FILL
XFILL_0__12635_ vdd gnd FILL
XFILL_1__10097_ vdd gnd FILL
XFILL_0__7133_ vdd gnd FILL
X_7761_ _7761_/A _7761_/B _7761_/C _7761_/D _7761_/Y vdd gnd OAI22X1
XFILL_1__13925_ vdd gnd FILL
XFILL_1_CLKBUF1_insert29 vdd gnd FILL
XFILL_2__11387_ vdd gnd FILL
X_9500_ _9500_/A _9500_/B _9500_/C _9500_/Y vdd gnd OAI21X1
X_7692_ _7692_/A _7692_/B _7692_/C _7692_/Y vdd gnd OAI21X1
XFILL_0__14305_ vdd gnd FILL
XFILL_1__13856_ vdd gnd FILL
XFILL_0__11517_ vdd gnd FILL
X_9431_ _9431_/A _9431_/B _9431_/C _9431_/Y vdd gnd NAND3X1
XFILL_0__12497_ vdd gnd FILL
XFILL_1__12807_ vdd gnd FILL
XFILL_0__14236_ vdd gnd FILL
XFILL_0__11448_ vdd gnd FILL
XFILL_1__13787_ vdd gnd FILL
XFILL_1__10999_ vdd gnd FILL
X_9362_ _9362_/A _9362_/B _9362_/Y vdd gnd NAND2X1
XFILL_2__12008_ vdd gnd FILL
XFILL_0_BUFX2_insert180 vdd gnd FILL
XFILL_1__12738_ vdd gnd FILL
XFILL_0_BUFX2_insert191 vdd gnd FILL
X_8313_ _8313_/A _8313_/B _8313_/Y vdd gnd AND2X2
XFILL_0__11379_ vdd gnd FILL
X_9293_ _9293_/A _9293_/B _9293_/Y vdd gnd NAND2X1
XFILL_0__13118_ vdd gnd FILL
XFILL_1__12669_ vdd gnd FILL
XFILL_0__9705_ vdd gnd FILL
XFILL_0__14098_ vdd gnd FILL
X_8244_ _8244_/A _8244_/B _8244_/C _8244_/D _8244_/Y vdd gnd AOI22X1
XFILL_0__7897_ vdd gnd FILL
XFILL_1__14408_ vdd gnd FILL
XFILL_0__13049_ vdd gnd FILL
XFILL_0__9636_ vdd gnd FILL
X_8175_ _8175_/A _8175_/B _8175_/C _8175_/Y vdd gnd AOI21X1
XFILL_1__14339_ vdd gnd FILL
X_7126_ _7126_/A _7126_/B _7126_/C _7126_/D _7126_/Y vdd gnd AOI22X1
XFILL_0__9567_ vdd gnd FILL
XFILL_1__8360_ vdd gnd FILL
XFILL_1__7311_ vdd gnd FILL
XFILL_0__8518_ vdd gnd FILL
XFILL_0__9498_ vdd gnd FILL
XFILL_1__8291_ vdd gnd FILL
XFILL_1__7242_ vdd gnd FILL
XFILL_0__8449_ vdd gnd FILL
XFILL_1__7173_ vdd gnd FILL
X_7959_ _7959_/D _7959_/CLK _7959_/Q vdd gnd DFFPOSX1
X_11560_ _11560_/A _11560_/B _11560_/Y vdd gnd NAND2X1
X_9629_ _9629_/A _9629_/Y vdd gnd INVX1
X_10511_ _10511_/A _10511_/B _10511_/C _10511_/Y vdd gnd OAI21X1
X_11491_ _11491_/A _11491_/B _11491_/Y vdd gnd NOR2X1
XBUFX2_insert20 BUFX2_insert20/A BUFX2_insert20/Y vdd gnd BUFX2
X_13230_ _13230_/A _13230_/B _13230_/C _13230_/Y vdd gnd OAI21X1
X_10442_ _10442_/A _10442_/B _10442_/Y vdd gnd NAND2X1
XFILL_1__9745_ vdd gnd FILL
X_13161_ _13161_/A _13161_/Y vdd gnd INVX1
X_10373_ _10373_/A _10373_/B _10373_/Y vdd gnd NAND2X1
XFILL_1__9676_ vdd gnd FILL
X_12112_ _12112_/A _12112_/B _12112_/Y vdd gnd NAND2X1
XFILL_2__7420_ vdd gnd FILL
X_13092_ _13092_/A _13092_/B _13092_/C _13092_/Y vdd gnd AOI21X1
XFILL_1__8627_ vdd gnd FILL
XFILL257550x187350 vdd gnd FILL
X_12043_ _12043_/A _12043_/B _12043_/Y vdd gnd NAND2X1
XFILL_2__7351_ vdd gnd FILL
XFILL_1__8558_ vdd gnd FILL
XFILL_1__7509_ vdd gnd FILL
XFILL_1__8489_ vdd gnd FILL
XFILL_2__9021_ vdd gnd FILL
XFILL_2_BUFX2_insert220 vdd gnd FILL
XFILL_1__10020_ vdd gnd FILL
X_13994_ _13994_/A _13994_/B _13994_/C _13994_/Y vdd gnd OAI21X1
XFILL_2_BUFX2_insert253 vdd gnd FILL
X_12945_ _12945_/A _12945_/B _12945_/C _12945_/Y vdd gnd AOI21X1
XFILL_2__11310_ vdd gnd FILL
XFILL_2_BUFX2_insert275 vdd gnd FILL
XFILL_0__10681_ vdd gnd FILL
XFILL_2__11241_ vdd gnd FILL
X_12876_ _12876_/A _12876_/B _12876_/C _12876_/Y vdd gnd NAND3X1
XFILL_0__12420_ vdd gnd FILL
XFILL_1__11971_ vdd gnd FILL
X_14615_ _14615_/A _14615_/B _14615_/C _14615_/Y vdd gnd OAI21X1
X_11827_ _11827_/A _11827_/B _11827_/Y vdd gnd NAND2X1
XFILL_1__13710_ vdd gnd FILL
XFILL_1__10922_ vdd gnd FILL
XFILL_2__11172_ vdd gnd FILL
XFILL_1__14690_ vdd gnd FILL
XFILL_0__12351_ vdd gnd FILL
X_14546_ _14546_/D _14546_/CLK _14546_/Q vdd gnd DFFPOSX1
X_11758_ _11758_/A _11758_/B _11758_/Y vdd gnd NAND2X1
XBUFX2_insert230 BUFX2_insert230/A BUFX2_insert230/Y vdd gnd BUFX2
XFILL_1__13641_ vdd gnd FILL
XFILL_2__9854_ vdd gnd FILL
XFILL_0__11302_ vdd gnd FILL
XFILL_1__10853_ vdd gnd FILL
XBUFX2_insert241 BUFX2_insert241/A BUFX2_insert241/Y vdd gnd BUFX2
X_10709_ _10709_/D _10709_/CLK _10709_/Q vdd gnd DFFPOSX1
XFILL_0__12282_ vdd gnd FILL
XBUFX2_insert252 BUFX2_insert252/A BUFX2_insert252/Y vdd gnd BUFX2
XBUFX2_insert263 BUFX2_insert263/A BUFX2_insert263/Y vdd gnd BUFX2
XBUFX2_insert274 BUFX2_insert274/A BUFX2_insert274/Y vdd gnd BUFX2
X_14477_ _14477_/A _14477_/B _14477_/Y vdd gnd NAND2X1
X_11689_ _11689_/D _11689_/CLK _11689_/Q vdd gnd DFFPOSX1
XFILL_0__14021_ vdd gnd FILL
XBUFX2_insert285 BUFX2_insert285/A BUFX2_insert285/Y vdd gnd BUFX2
XFILL_1__13572_ vdd gnd FILL
XFILL_0__11233_ vdd gnd FILL
XFILL_0__7820_ vdd gnd FILL
XBUFX2_insert296 BUFX2_insert296/A BUFX2_insert296/Y vdd gnd BUFX2
XFILL_1__10784_ vdd gnd FILL
X_13428_ _13428_/D _13428_/CLK _13428_/Q vdd gnd DFFPOSX1
XFILL_2__8736_ vdd gnd FILL
XFILL_1__12523_ vdd gnd FILL
XFILL_0__11164_ vdd gnd FILL
XFILL_0__7751_ vdd gnd FILL
X_13359_ _13359_/A _13359_/B _13359_/Y vdd gnd NAND2X1
XFILL_0__10115_ vdd gnd FILL
XFILL_2__13813_ vdd gnd FILL
XFILL_1__12454_ vdd gnd FILL
XFILL_2__8667_ vdd gnd FILL
XFILL_0__11095_ vdd gnd FILL
XFILL_0__7682_ vdd gnd FILL
XFILL_1__11405_ vdd gnd FILL
XFILL_0__10046_ vdd gnd FILL
XFILL_2__13744_ vdd gnd FILL
XFILL_0__9421_ vdd gnd FILL
XFILL_2__8598_ vdd gnd FILL
XFILL_1__12385_ vdd gnd FILL
XFILL_1__14124_ vdd gnd FILL
XFILL_1__11336_ vdd gnd FILL
XFILL_2__13675_ vdd gnd FILL
XFILL_0__14854_ vdd gnd FILL
XFILL_0__9352_ vdd gnd FILL
X_9980_ _9980_/A _9980_/B _9980_/C _9980_/Y vdd gnd AOI21X1
XFILL_2__12626_ vdd gnd FILL
XFILL_1__14055_ vdd gnd FILL
XFILL_0__13805_ vdd gnd FILL
XFILL_0__8303_ vdd gnd FILL
XFILL_1__11267_ vdd gnd FILL
XFILL_0__14785_ vdd gnd FILL
XFILL_0__9283_ vdd gnd FILL
X_8931_ _8931_/A _8931_/B _8931_/C _8931_/Y vdd gnd OAI21X1
XFILL_0__11997_ vdd gnd FILL
XFILL_2__9219_ vdd gnd FILL
XFILL_1__13006_ vdd gnd FILL
XFILL_1__10218_ vdd gnd FILL
XFILL_0__13736_ vdd gnd FILL
XFILL_0__8234_ vdd gnd FILL
XFILL_1__11198_ vdd gnd FILL
XFILL_0__10948_ vdd gnd FILL
X_8862_ _8862_/D _8862_/CLK _8862_/Q vdd gnd DFFPOSX1
XFILL_2__11508_ vdd gnd FILL
XFILL_1__10149_ vdd gnd FILL
XFILL_0__13667_ vdd gnd FILL
X_7813_ _7813_/A _7813_/B _7813_/Y vdd gnd NAND2X1
XFILL_0__8165_ vdd gnd FILL
XFILL_0__10879_ vdd gnd FILL
X_8793_ _8793_/A _8793_/B _8793_/C _8793_/Y vdd gnd OAI21X1
XFILL_2__11439_ vdd gnd FILL
XFILL_0__12618_ vdd gnd FILL
XFILL_0__7116_ vdd gnd FILL
XFILL_0__13598_ vdd gnd FILL
XFILL257550x252150 vdd gnd FILL
X_7744_ _7744_/A _7744_/B _7744_/C _7744_/Y vdd gnd AOI21X1
XFILL_0__8096_ vdd gnd FILL
XFILL_1__13908_ vdd gnd FILL
X_7675_ _7675_/A _7675_/B _7675_/Y vdd gnd NAND2X1
XFILL_1__13839_ vdd gnd FILL
X_9414_ _9414_/A _9414_/B _9414_/C _9414_/Y vdd gnd NAND3X1
XFILL_1__7860_ vdd gnd FILL
XFILL_0__14219_ vdd gnd FILL
X_9345_ _9345_/A _9345_/B _9345_/C _9345_/Y vdd gnd NAND3X1
XFILL_1__7791_ vdd gnd FILL
XFILL_0__8998_ vdd gnd FILL
XFILL_1__9530_ vdd gnd FILL
X_9276_ _9276_/A _9276_/Y vdd gnd INVX1
XFILL_1__9461_ vdd gnd FILL
X_8227_ _8227_/A _8227_/B _8227_/Y vdd gnd NAND2X1
XFILL_0__9619_ vdd gnd FILL
XFILL_1__8412_ vdd gnd FILL
XFILL_1__9392_ vdd gnd FILL
X_8158_ _8158_/A _8158_/Y vdd gnd INVX1
X_7109_ _7109_/A _7109_/B _7109_/Y vdd gnd NAND2X1
XFILL_1__8343_ vdd gnd FILL
X_8089_ _8089_/A _8089_/B _8089_/C _8089_/Y vdd gnd AOI21X1
XFILL_1__8274_ vdd gnd FILL
XFILL_1__7225_ vdd gnd FILL
X_10991_ _10991_/A _10991_/B _10991_/Y vdd gnd AND2X2
XFILL_1_BUFX2_insert205 vdd gnd FILL
X_12730_ _12730_/A _12730_/B _12730_/S _12730_/Y vdd gnd MUX2X1
XFILL_1__7156_ vdd gnd FILL
XFILL_1_BUFX2_insert216 vdd gnd FILL
XFILL_1_BUFX2_insert227 vdd gnd FILL
XFILL_1_BUFX2_insert238 vdd gnd FILL
X_12661_ _12661_/A _12661_/B _12661_/Y vdd gnd NOR2X1
XFILL_1_BUFX2_insert249 vdd gnd FILL
XFILL_1__7087_ vdd gnd FILL
X_14400_ _14400_/A _14400_/B _14400_/C _14400_/Y vdd gnd OAI21X1
X_11612_ _11612_/D _11612_/CLK _11612_/Q vdd gnd DFFPOSX1
X_12592_ _12592_/D _12592_/CLK _12592_/Q vdd gnd DFFPOSX1
X_14331_ _14331_/A _14331_/B _14331_/Y vdd gnd NAND2X1
X_11543_ _11543_/A _11543_/B _11543_/Y vdd gnd NAND2X1
XFILL_0_CLKBUF1_insert386 vdd gnd FILL
X_14262_ _14262_/A _14262_/B _14262_/C _14262_/Y vdd gnd OAI21X1
X_11474_ _11474_/A _11474_/B _11474_/Y vdd gnd NAND2X1
XFILL_2__9570_ vdd gnd FILL
X_13213_ _13213_/A _13213_/Y vdd gnd INVX1
X_10425_ _10425_/A _10425_/B _10425_/C _10425_/Y vdd gnd OAI21X1
X_14193_ _14193_/D _14193_/CLK _14193_/Q vdd gnd DFFPOSX1
XFILL_1__9728_ vdd gnd FILL
X_13144_ _13144_/A _13144_/B _13144_/C _13144_/Y vdd gnd OAI21X1
X_10356_ _10356_/A _10356_/B _10356_/Y vdd gnd NAND2X1
XFILL_2__10810_ vdd gnd FILL
XFILL_1__9659_ vdd gnd FILL
X_13075_ _13075_/A _13075_/B _13075_/C _13075_/Y vdd gnd OAI21X1
XFILL_2__7403_ vdd gnd FILL
X_10287_ _10287_/A _10287_/B _10287_/Y vdd gnd NAND2X1
XFILL_0__11920_ vdd gnd FILL
XFILL_1__12170_ vdd gnd FILL
X_12026_ _12026_/A _12026_/B _12026_/C _12026_/Y vdd gnd NAND3X1
XFILL_2__7334_ vdd gnd FILL
XFILL_1__11121_ vdd gnd FILL
XFILL_0__11851_ vdd gnd FILL
XFILL_2__7265_ vdd gnd FILL
XFILL_1__11052_ vdd gnd FILL
XFILL_0__10802_ vdd gnd FILL
XFILL_2__13391_ vdd gnd FILL
XFILL_0__14570_ vdd gnd FILL
XFILL_0__11782_ vdd gnd FILL
X_13977_ _13977_/A _13977_/B _13977_/Y vdd gnd NAND2X1
XFILL_1__10003_ vdd gnd FILL
XFILL_2__7196_ vdd gnd FILL
XFILL_0__13521_ vdd gnd FILL
X_12928_ _12928_/A _12928_/B _12928_/C _12928_/Y vdd gnd OAI21X1
XFILL_1__14811_ vdd gnd FILL
XFILL_0__10664_ vdd gnd FILL
X_12859_ _12859_/A _12859_/B _12859_/C _12859_/Y vdd gnd AOI21X1
XFILL_1__14742_ vdd gnd FILL
XFILL_0__12403_ vdd gnd FILL
XFILL_1__11954_ vdd gnd FILL
XFILL_0__13383_ vdd gnd FILL
XFILL_0__10595_ vdd gnd FILL
XFILL_0__9970_ vdd gnd FILL
XFILL_1__10905_ vdd gnd FILL
XFILL_2__11155_ vdd gnd FILL
XFILL_1__14673_ vdd gnd FILL
XFILL_0__12334_ vdd gnd FILL
XFILL_1__11885_ vdd gnd FILL
XFILL_0__8921_ vdd gnd FILL
X_14529_ _14529_/D _14529_/CLK _14529_/Q vdd gnd DFFPOSX1
X_7460_ _7460_/A _7460_/B _7460_/C _7460_/Y vdd gnd OAI21X1
XFILL_2__10106_ vdd gnd FILL
XFILL_1__13624_ vdd gnd FILL
XFILL_2__11086_ vdd gnd FILL
XFILL_1__10836_ vdd gnd FILL
XFILL_0__12265_ vdd gnd FILL
X_7391_ _7391_/A _7391_/B _7391_/C _7391_/Y vdd gnd OAI21X1
XFILL_2__14914_ vdd gnd FILL
XFILL_0__14004_ vdd gnd FILL
XFILL_0__11216_ vdd gnd FILL
XFILL_1__13555_ vdd gnd FILL
X_9130_ _9130_/A _9130_/B _9130_/Y vdd gnd NAND2X1
XFILL_0__7803_ vdd gnd FILL
XFILL_0__12196_ vdd gnd FILL
XFILL_0__8783_ vdd gnd FILL
XFILL_1__12506_ vdd gnd FILL
XFILL_0__11147_ vdd gnd FILL
X_9061_ _9061_/A _9061_/B _9061_/C _9061_/D _9061_/Y vdd gnd OAI22X1
XFILL_0__7734_ vdd gnd FILL
XFILL_1__12437_ vdd gnd FILL
XFILL_0__11078_ vdd gnd FILL
X_8012_ _8012_/A _8012_/B _8012_/C _8012_/Y vdd gnd OAI21X1
XFILL_0__7665_ vdd gnd FILL
XFILL_2__13727_ vdd gnd FILL
XFILL_0__10029_ vdd gnd FILL
XFILL_1__12368_ vdd gnd FILL
XFILL_2__10939_ vdd gnd FILL
XFILL_0__9404_ vdd gnd FILL
XFILL_0__7596_ vdd gnd FILL
XFILL_1__14107_ vdd gnd FILL
XFILL_1__11319_ vdd gnd FILL
XFILL_2__13658_ vdd gnd FILL
XFILL_0__14837_ vdd gnd FILL
XFILL_1__12299_ vdd gnd FILL
XFILL_0__9335_ vdd gnd FILL
X_9963_ _9963_/A _9963_/B _9963_/S _9963_/Y vdd gnd MUX2X1
XFILL_1__14038_ vdd gnd FILL
XFILL_2__13589_ vdd gnd FILL
XFILL_0__14768_ vdd gnd FILL
XFILL_0__9266_ vdd gnd FILL
X_8914_ _8914_/D _8914_/CLK _8914_/Q vdd gnd DFFPOSX1
X_9894_ _9894_/A _9894_/B _9894_/Y vdd gnd NAND2X1
XFILL_0__13719_ vdd gnd FILL
XFILL_0__8217_ vdd gnd FILL
XFILL_0__14699_ vdd gnd FILL
XFILL_0__9197_ vdd gnd FILL
X_8845_ _8845_/D _8845_/CLK _8845_/Q vdd gnd DFFPOSX1
XFILL_0__8148_ vdd gnd FILL
X_8776_ _8776_/A _8776_/B _8776_/Y vdd gnd NAND2X1
X_7727_ _7727_/A _7727_/B _7727_/C _7727_/Y vdd gnd OAI21X1
XFILL_0__8079_ vdd gnd FILL
XFILL_1__8961_ vdd gnd FILL
XFILL_1__7912_ vdd gnd FILL
X_7658_ _7658_/A _7658_/B _7658_/C _7658_/Y vdd gnd NAND3X1
XFILL_1__7843_ vdd gnd FILL
X_7589_ _7589_/A _7589_/B _7589_/Y vdd gnd NOR2X1
X_9328_ _9328_/A _9328_/B _9328_/Y vdd gnd AND2X2
XFILL_1__7774_ vdd gnd FILL
X_10210_ _10210_/A _10210_/B _10210_/Y vdd gnd NAND2X1
XFILL_1__9513_ vdd gnd FILL
X_11190_ _11190_/A _11190_/B _11190_/Y vdd gnd NAND2X1
X_9259_ _9259_/A _9259_/B _9259_/C _9259_/Y vdd gnd AOI21X1
X_10141_ _10141_/A _10141_/B _10141_/C _10141_/Y vdd gnd OAI21X1
XFILL_1__9444_ vdd gnd FILL
X_10072_ _10072_/A _10072_/Y vdd gnd INVX1
XFILL_1__9375_ vdd gnd FILL
X_13900_ _13900_/A _13900_/B _13900_/C _13900_/Y vdd gnd AOI21X1
X_14880_ _14880_/D _14880_/CLK _14880_/Q vdd gnd DFFPOSX1
XFILL_1__8326_ vdd gnd FILL
X_13831_ _13831_/A _13831_/B _13831_/C _13831_/D _13831_/Y vdd gnd AOI22X1
XFILL_1__8257_ vdd gnd FILL
XFILL_1__7208_ vdd gnd FILL
X_13762_ _13762_/A _13762_/Y vdd gnd INVX1
X_10974_ _10974_/A _10974_/B _10974_/C _10974_/D _10974_/Y vdd gnd AOI22X1
XFILL_1__8188_ vdd gnd FILL
X_12713_ _12713_/A _12713_/B _12713_/Y vdd gnd NAND2X1
XFILL_1__7139_ vdd gnd FILL
X_13693_ _13693_/A _13693_/B _13693_/C _13693_/Y vdd gnd OAI21X1
X_12644_ _12644_/A _12644_/B _12644_/C _12644_/Y vdd gnd AOI21X1
XFILL_0__10380_ vdd gnd FILL
X_12575_ _12575_/D _12575_/CLK _12575_/Q vdd gnd DFFPOSX1
X_14314_ _14314_/A _14314_/B _14314_/Y vdd gnd NAND2X1
X_11526_ _11526_/A _11526_/B _11526_/C _11526_/Y vdd gnd OAI21X1
XFILL_2__9622_ vdd gnd FILL
XFILL_1__10621_ vdd gnd FILL
XFILL_0__12050_ vdd gnd FILL
XFILL_2__12960_ vdd gnd FILL
X_14245_ _14245_/A _14245_/B _14245_/C _14245_/Y vdd gnd OAI21X1
X_11457_ _11457_/A _11457_/B _11457_/C _11457_/D _11457_/Y vdd gnd OAI22X1
XFILL_0__11001_ vdd gnd FILL
XFILL_2__9553_ vdd gnd FILL
XFILL_1__13340_ vdd gnd FILL
XFILL_1__10552_ vdd gnd FILL
XFILL_2__12891_ vdd gnd FILL
X_10408_ _10408_/A _10408_/B _10408_/Y vdd gnd OR2X2
X_14176_ _14176_/D _14176_/CLK _14176_/Q vdd gnd DFFPOSX1
X_11388_ _11388_/A _11388_/B _11388_/C _11388_/Y vdd gnd OAI21X1
XFILL_2__9484_ vdd gnd FILL
XFILL_1__13271_ vdd gnd FILL
XFILL_1__10483_ vdd gnd FILL
X_13127_ _13127_/A _13127_/B _13127_/Y vdd gnd AND2X2
X_10339_ _10339_/A _10339_/B _10339_/Y vdd gnd NAND2X1
XFILL_1__12222_ vdd gnd FILL
XFILL_0__12952_ vdd gnd FILL
XFILL_0__7450_ vdd gnd FILL
X_13058_ _13058_/A _13058_/B _13058_/C _13058_/Y vdd gnd AOI21X1
XFILL_0__11903_ vdd gnd FILL
XFILL_2__14492_ vdd gnd FILL
XFILL_1__12153_ vdd gnd FILL
X_12009_ _12009_/A _12009_/B _12009_/Y vdd gnd AND2X2
XFILL_0__12883_ vdd gnd FILL
XFILL_0__7381_ vdd gnd FILL
XFILL_1__11104_ vdd gnd FILL
XFILL_2__7317_ vdd gnd FILL
XFILL_0__14622_ vdd gnd FILL
XFILL_0__9120_ vdd gnd FILL
XFILL_0__11834_ vdd gnd FILL
XFILL_1__12084_ vdd gnd FILL
XFILL_2__7248_ vdd gnd FILL
XFILL_1__11035_ vdd gnd FILL
XFILL_2__13374_ vdd gnd FILL
XFILL_0__9051_ vdd gnd FILL
XFILL_0__11765_ vdd gnd FILL
XFILL_2__12325_ vdd gnd FILL
XFILL_2__7179_ vdd gnd FILL
XFILL_0__13504_ vdd gnd FILL
XFILL_0__8002_ vdd gnd FILL
XFILL_0__14484_ vdd gnd FILL
X_8630_ _8630_/A _8630_/B _8630_/Y vdd gnd NAND2X1
XFILL_0__11696_ vdd gnd FILL
XFILL_1__12986_ vdd gnd FILL
XFILL_0__10647_ vdd gnd FILL
X_8561_ _8561_/A _8561_/B _8561_/C _8561_/Y vdd gnd OAI21X1
XFILL_1__14725_ vdd gnd FILL
XFILL_1__11937_ vdd gnd FILL
XFILL_0__13366_ vdd gnd FILL
X_7512_ _7512_/A _7512_/B _7512_/S _7512_/Y vdd gnd MUX2X1
XFILL_0__10578_ vdd gnd FILL
XFILL_0__9953_ vdd gnd FILL
X_8492_ _8492_/A _8492_/B _8492_/Y vdd gnd NOR2X1
XFILL_0__12317_ vdd gnd FILL
XFILL_1__14656_ vdd gnd FILL
XFILL_1__11868_ vdd gnd FILL
XFILL_0__13297_ vdd gnd FILL
X_7443_ _7443_/A _7443_/B _7443_/Y vdd gnd NAND2X1
XFILL_0__9884_ vdd gnd FILL
XFILL_1__10819_ vdd gnd FILL
XFILL_1__13607_ vdd gnd FILL
XFILL_1__14587_ vdd gnd FILL
XFILL_0__12248_ vdd gnd FILL
XFILL_1__11799_ vdd gnd FILL
XFILL_0__8835_ vdd gnd FILL
X_7374_ _7374_/A _7374_/B _7374_/C _7374_/Y vdd gnd NAND3X1
XFILL_1__13538_ vdd gnd FILL
X_9113_ _9113_/A _9113_/B _9113_/C _9113_/Y vdd gnd OAI21X1
XFILL_0__12179_ vdd gnd FILL
XFILL_2_CLKBUF1_insert70 vdd gnd FILL
XFILL_0__8766_ vdd gnd FILL
X_9044_ _9044_/A _9044_/B _9044_/C _9044_/Y vdd gnd AOI21X1
XFILL_0__7717_ vdd gnd FILL
XFILL_1__7490_ vdd gnd FILL
XFILL_0__8697_ vdd gnd FILL
XFILL_0__7648_ vdd gnd FILL
XFILL_1__9160_ vdd gnd FILL
XFILL_0__7579_ vdd gnd FILL
XFILL_1__8111_ vdd gnd FILL
XFILL_0__9318_ vdd gnd FILL
XFILL_1__9091_ vdd gnd FILL
X_9946_ _9946_/A _9946_/B _9946_/C _9946_/Y vdd gnd OAI21X1
XFILL_1__8042_ vdd gnd FILL
XFILL_0__9249_ vdd gnd FILL
X_9877_ _9877_/A _9877_/Y vdd gnd INVX1
X_8828_ _8828_/A _8828_/B _8828_/Y vdd gnd NAND2X1
X_10690_ _10690_/D _10690_/CLK _10690_/Q vdd gnd DFFPOSX1
X_8759_ _8759_/A _8759_/B _8759_/Y vdd gnd NAND2X1
XFILL_1__9993_ vdd gnd FILL
XFILL_1__8944_ vdd gnd FILL
X_12360_ _12360_/A _12360_/B _12360_/C _12360_/Y vdd gnd OAI21X1
X_11311_ _11311_/A _11311_/B _11311_/Y vdd gnd NOR2X1
X_12291_ _12291_/A _12291_/B _12291_/Y vdd gnd AND2X2
XFILL_1__7826_ vdd gnd FILL
X_14030_ _14030_/A _14030_/Y vdd gnd INVX1
X_11242_ _11242_/A _11242_/B _11242_/Y vdd gnd NAND2X1
XFILL_1__7757_ vdd gnd FILL
X_11173_ _11173_/A _11173_/B _11173_/C _11173_/Y vdd gnd AOI21X1
XFILL_1__7688_ vdd gnd FILL
X_10124_ _10124_/A _10124_/B _10124_/C _10124_/Y vdd gnd OAI21X1
XFILL_1__9427_ vdd gnd FILL
X_10055_ _10055_/A _10055_/Y vdd gnd INVX1
XFILL_1__9358_ vdd gnd FILL
X_14863_ _14863_/A _14863_/B _14863_/C _14863_/Y vdd gnd AOI21X1
XFILL_1__8309_ vdd gnd FILL
XFILL_1__9289_ vdd gnd FILL
X_13814_ _13814_/A _13814_/B _13814_/Y vdd gnd NAND2X1
X_14794_ _14794_/A _14794_/B _14794_/Y vdd gnd NOR2X1
XFILL_0__11550_ vdd gnd FILL
XFILL_2__12110_ vdd gnd FILL
X_13745_ _13745_/A _13745_/B _13745_/Y vdd gnd NOR2X1
X_10957_ _10957_/A _10957_/B _10957_/C _10957_/Y vdd gnd OAI21X1
XFILL_0__10501_ vdd gnd FILL
XFILL_1__12840_ vdd gnd FILL
XFILL_0__11481_ vdd gnd FILL
XFILL_2__12041_ vdd gnd FILL
X_13676_ _13676_/A _13676_/B _13676_/Y vdd gnd NAND2X1
XFILL_0__13220_ vdd gnd FILL
X_10888_ _10888_/A _10888_/B _10888_/S _10888_/Y vdd gnd MUX2X1
XFILL_0__10432_ vdd gnd FILL
XFILL_1__12771_ vdd gnd FILL
X_12627_ _12627_/A _12627_/Y vdd gnd INVX1
XFILL_1__11722_ vdd gnd FILL
XFILL_0__13151_ vdd gnd FILL
XFILL_0__10363_ vdd gnd FILL
X_12558_ _12558_/D _12558_/CLK _12558_/Q vdd gnd DFFPOSX1
XFILL_1__14441_ vdd gnd FILL
XFILL_0__12102_ vdd gnd FILL
XFILL_0__13082_ vdd gnd FILL
XFILL_2__13992_ vdd gnd FILL
XFILL_0__10294_ vdd gnd FILL
X_11509_ _11509_/A _11509_/B _11509_/Y vdd gnd NAND2X1
XFILL_2__9605_ vdd gnd FILL
XFILL_1__10604_ vdd gnd FILL
X_12489_ _12489_/A _12489_/B _12489_/C _12489_/Y vdd gnd OAI21X1
XFILL_2__12943_ vdd gnd FILL
XFILL_0__12033_ vdd gnd FILL
XFILL_1__14372_ vdd gnd FILL
XFILL_1__11584_ vdd gnd FILL
X_14228_ _14228_/A _14228_/Y vdd gnd INVX1
XFILL_0__8620_ vdd gnd FILL
XFILL_2__9536_ vdd gnd FILL
XFILL_1__13323_ vdd gnd FILL
XFILL_1__10535_ vdd gnd FILL
XFILL_2__12874_ vdd gnd FILL
XFILL_0__8551_ vdd gnd FILL
X_14159_ _14159_/D _14159_/CLK _14159_/Q vdd gnd DFFPOSX1
X_7090_ _7090_/A _7090_/Y vdd gnd INVX1
XFILL_2__9467_ vdd gnd FILL
XFILL_1__13254_ vdd gnd FILL
XFILL_1__10466_ vdd gnd FILL
XFILL256350x223350 vdd gnd FILL
XFILL_0__13984_ vdd gnd FILL
XFILL_0__7502_ vdd gnd FILL
XFILL_0__8482_ vdd gnd FILL
XFILL_1__12205_ vdd gnd FILL
XFILL_1__13185_ vdd gnd FILL
XFILL_0__12935_ vdd gnd FILL
XFILL_2__9398_ vdd gnd FILL
XFILL_0__7433_ vdd gnd FILL
XFILL_1__10397_ vdd gnd FILL
XFILL_1__12136_ vdd gnd FILL
XFILL_2__14475_ vdd gnd FILL
XFILL_0__12866_ vdd gnd FILL
XFILL_0__7364_ vdd gnd FILL
X_9800_ _9800_/D _9800_/CLK _9800_/Q vdd gnd DFFPOSX1
XFILL_0__14605_ vdd gnd FILL
X_7992_ _7992_/D _7992_/CLK _7992_/Q vdd gnd DFFPOSX1
XFILL_0__11817_ vdd gnd FILL
XFILL_1__12067_ vdd gnd FILL
XFILL_0__9103_ vdd gnd FILL
XFILL_0__12797_ vdd gnd FILL
XFILL_0__7295_ vdd gnd FILL
X_9731_ _9731_/A _9731_/B _9731_/C _9731_/Y vdd gnd OAI21X1
XFILL_1__11018_ vdd gnd FILL
XFILL_0__9034_ vdd gnd FILL
XFILL_0__11748_ vdd gnd FILL
X_9662_ _9662_/A _9662_/B _9662_/Y vdd gnd AND2X2
XFILL_2__12308_ vdd gnd FILL
XFILL_0__14467_ vdd gnd FILL
X_8613_ _8613_/A _8613_/B _8613_/Y vdd gnd NAND2X1
X_9593_ _9593_/A _9593_/B _9593_/Y vdd gnd AND2X2
XFILL_2__12239_ vdd gnd FILL
XFILL_0__13418_ vdd gnd FILL
XFILL_1__12969_ vdd gnd FILL
XFILL_0__14398_ vdd gnd FILL
X_8544_ _8544_/A _8544_/B _8544_/Y vdd gnd NOR2X1
XFILL_1__14708_ vdd gnd FILL
XFILL_0__13349_ vdd gnd FILL
XFILL_0__9936_ vdd gnd FILL
X_8475_ _8475_/A _8475_/Y vdd gnd INVX1
XFILL_1__14639_ vdd gnd FILL
X_7426_ _7426_/A _7426_/B _7426_/Y vdd gnd NAND2X1
XFILL_0__9867_ vdd gnd FILL
XFILL_1__8660_ vdd gnd FILL
XFILL_1__7611_ vdd gnd FILL
XFILL_0__8818_ vdd gnd FILL
X_7357_ _7357_/A _7357_/B _7357_/C _7357_/Y vdd gnd OAI21X1
XFILL_1__8591_ vdd gnd FILL
XFILL_1__7542_ vdd gnd FILL
XFILL_0__8749_ vdd gnd FILL
X_7288_ _7288_/A _7288_/B _7288_/C _7288_/Y vdd gnd NOR3X1
X_9027_ _9027_/A _9027_/Y vdd gnd INVX1
XFILL_1__7473_ vdd gnd FILL
XFILL_1__9212_ vdd gnd FILL
XFILL_1__9143_ vdd gnd FILL
XFILL_1__9074_ vdd gnd FILL
X_11860_ _11860_/A _11860_/B _11860_/Y vdd gnd NAND2X1
X_9929_ _9929_/A _9929_/Y vdd gnd INVX8
X_10811_ _10811_/A _10811_/B _10811_/C _10811_/Y vdd gnd OAI21X1
XFILL_1__8025_ vdd gnd FILL
X_11791_ _11791_/A _11791_/Y vdd gnd INVX8
X_13530_ _13530_/A _13530_/B _13530_/C _13530_/Y vdd gnd AOI21X1
X_10742_ _10742_/D _10742_/CLK _10742_/Q vdd gnd DFFPOSX1
X_10673_ _10673_/A _10673_/B _10673_/C _10673_/Y vdd gnd OAI21X1
X_13461_ _13461_/D _13461_/CLK _13461_/Q vdd gnd DFFPOSX1
XFILL_1__9976_ vdd gnd FILL
X_12412_ _12412_/A _12412_/B _12412_/C _12412_/Y vdd gnd AOI21X1
XFILL_1__8927_ vdd gnd FILL
XFILL_2__7720_ vdd gnd FILL
X_13392_ _13392_/A _13392_/B _13392_/Y vdd gnd NAND2X1
X_12343_ _12343_/A _12343_/Y vdd gnd INVX1
XFILL257250x198150 vdd gnd FILL
XFILL_2__7651_ vdd gnd FILL
X_12274_ _12274_/A _12274_/Y vdd gnd INVX1
XFILL_1__7809_ vdd gnd FILL
XFILL_2__7582_ vdd gnd FILL
XFILL_1__8789_ vdd gnd FILL
X_14013_ _14013_/A _14013_/Y vdd gnd INVX1
X_11225_ _11225_/A _11225_/B _11225_/C _11225_/Y vdd gnd AOI21X1
XFILL_1__10320_ vdd gnd FILL
X_11156_ _11156_/A _11156_/B _11156_/C _11156_/Y vdd gnd OAI21X1
XFILL_1__10251_ vdd gnd FILL
X_10107_ _10107_/A _10107_/Y vdd gnd INVX1
XFILL_0__10981_ vdd gnd FILL
X_11087_ _11087_/A _11087_/B _11087_/C _11087_/Y vdd gnd OAI21X1
XFILL_2__8203_ vdd gnd FILL
XFILL_2__9183_ vdd gnd FILL
XFILL_0__12720_ vdd gnd FILL
XFILL_1__10182_ vdd gnd FILL
X_14915_ _14915_/A _14915_/Y vdd gnd BUFX2
X_10038_ _10038_/A _10038_/Y vdd gnd INVX2
XFILL_2__8134_ vdd gnd FILL
XFILL_2__11472_ vdd gnd FILL
XFILL_0__12651_ vdd gnd FILL
X_14846_ _14846_/A _14846_/B _14846_/Y vdd gnd NOR2X1
XFILL_2__10423_ vdd gnd FILL
XFILL_0__11602_ vdd gnd FILL
XFILL_1__13941_ vdd gnd FILL
XFILL_0_BUFX2_insert0 vdd gnd FILL
XFILL_0__7080_ vdd gnd FILL
X_14777_ _14777_/A _14777_/Y vdd gnd INVX1
X_11989_ _11989_/A _11989_/B _11989_/C _11989_/Y vdd gnd OAI21X1
XFILL_0__14321_ vdd gnd FILL
XFILL_0__11533_ vdd gnd FILL
XFILL_1__13872_ vdd gnd FILL
X_13728_ _13728_/A _13728_/B _13728_/C _13728_/Y vdd gnd AOI21X1
XFILL_0__14252_ vdd gnd FILL
XFILL_1__12823_ vdd gnd FILL
XFILL_0__11464_ vdd gnd FILL
X_13659_ _13659_/A _13659_/B _13659_/C _13659_/Y vdd gnd OAI21X1
XFILL_2__12024_ vdd gnd FILL
XFILL_0__13203_ vdd gnd FILL
XFILL_2__8967_ vdd gnd FILL
XFILL_0__10415_ vdd gnd FILL
XFILL_1__12754_ vdd gnd FILL
XFILL_0_BUFX2_insert340 vdd gnd FILL
XFILL_0__11395_ vdd gnd FILL
XFILL_0_BUFX2_insert351 vdd gnd FILL
XFILL_0_BUFX2_insert362 vdd gnd FILL
XFILL_0_BUFX2_insert373 vdd gnd FILL
XFILL_1__11705_ vdd gnd FILL
XFILL_0__13134_ vdd gnd FILL
XFILL_0__10346_ vdd gnd FILL
XFILL_1__12685_ vdd gnd FILL
XFILL_0__9721_ vdd gnd FILL
X_8260_ _8260_/A _8260_/B _8260_/C _8260_/Y vdd gnd OAI21X1
XFILL_2__7849_ vdd gnd FILL
XFILL_1__14424_ vdd gnd FILL
XFILL_2__13975_ vdd gnd FILL
XFILL_0__13065_ vdd gnd FILL
X_7211_ _7211_/A _7211_/B _7211_/S _7211_/Y vdd gnd MUX2X1
XFILL_0__10277_ vdd gnd FILL
XFILL_0__9652_ vdd gnd FILL
X_8191_ _8191_/A _8191_/B _8191_/C _8191_/Y vdd gnd OAI21X1
XFILL_2__12926_ vdd gnd FILL
XFILL_0__12016_ vdd gnd FILL
XFILL_1__14355_ vdd gnd FILL
XFILL_1__11567_ vdd gnd FILL
XFILL_0__8603_ vdd gnd FILL
X_7142_ _7142_/A _7142_/B _7142_/Y vdd gnd NAND2X1
XFILL_2__9519_ vdd gnd FILL
XFILL_0__9583_ vdd gnd FILL
XFILL_1__13306_ vdd gnd FILL
XFILL_1__10518_ vdd gnd FILL
XFILL_1__14286_ vdd gnd FILL
XFILL_2__12857_ vdd gnd FILL
XFILL_1__11498_ vdd gnd FILL
XFILL_0__8534_ vdd gnd FILL
X_7073_ _7073_/A _7073_/Y vdd gnd INVX2
XFILL_1__13237_ vdd gnd FILL
XFILL_1__10449_ vdd gnd FILL
XFILL_0__13967_ vdd gnd FILL
XFILL_2__12788_ vdd gnd FILL
XFILL_0__8465_ vdd gnd FILL
XFILL_1__13168_ vdd gnd FILL
XFILL_0__12918_ vdd gnd FILL
XFILL_0__7416_ vdd gnd FILL
XFILL_0__13898_ vdd gnd FILL
XFILL_0__8396_ vdd gnd FILL
XFILL_1__12119_ vdd gnd FILL
XFILL_1__13099_ vdd gnd FILL
XFILL_0__12849_ vdd gnd FILL
XFILL_0__7347_ vdd gnd FILL
X_7975_ _7975_/D _7975_/CLK _7975_/Q vdd gnd DFFPOSX1
XFILL_0__7278_ vdd gnd FILL
X_9714_ _9714_/A _9714_/B _9714_/Y vdd gnd NAND2X1
XFILL_0__9017_ vdd gnd FILL
X_9645_ _9645_/A _9645_/B _9645_/C _9645_/Y vdd gnd NAND3X1
X_9576_ _9576_/A _9576_/B _9576_/C _9576_/Y vdd gnd OAI21X1
X_8527_ _8527_/A _8527_/Y vdd gnd INVX1
XFILL_1__9761_ vdd gnd FILL
XFILL_0__9919_ vdd gnd FILL
XFILL_1__8712_ vdd gnd FILL
X_8458_ _8458_/A _8458_/B _8458_/Y vdd gnd NAND2X1
XFILL_1__9692_ vdd gnd FILL
X_7409_ _7409_/A _7409_/B _7409_/C _7409_/Y vdd gnd AOI21X1
XFILL_1__8643_ vdd gnd FILL
X_8389_ _8389_/A _8389_/B _8389_/Y vdd gnd NAND2X1
XFILL_1__8574_ vdd gnd FILL
X_11010_ _11010_/A _11010_/B _11010_/C _11010_/Y vdd gnd AOI21X1
XFILL_1__7525_ vdd gnd FILL
XFILL_1__7456_ vdd gnd FILL
X_12961_ _12961_/A _12961_/Y vdd gnd INVX1
XFILL_1__7387_ vdd gnd FILL
X_14700_ _14700_/A _14700_/B _14700_/C _14700_/Y vdd gnd OAI21X1
X_11912_ _11912_/A _11912_/B _11912_/C _11912_/Y vdd gnd AOI21X1
XFILL_1__9126_ vdd gnd FILL
X_12892_ _12892_/A _12892_/Y vdd gnd INVX1
X_14631_ _14631_/A _14631_/B _14631_/Y vdd gnd NOR2X1
X_11843_ _11843_/A _11843_/B _11843_/Y vdd gnd OR2X2
XFILL_1__9057_ vdd gnd FILL
X_14562_ _14562_/A _14562_/B _14562_/Y vdd gnd NAND2X1
XFILL_1__8008_ vdd gnd FILL
X_11774_ _11774_/A _11774_/Y vdd gnd INVX2
X_13513_ _13513_/A _13513_/Y vdd gnd INVX1
X_10725_ _10725_/D _10725_/CLK _10725_/Q vdd gnd DFFPOSX1
X_14493_ _14493_/A _14493_/B _14493_/C _14493_/Y vdd gnd OAI21X1
XFILL_2__10070_ vdd gnd FILL
X_13444_ _13444_/D _13444_/CLK _13444_/Q vdd gnd DFFPOSX1
X_10656_ _10656_/A _10656_/B _10656_/C _10656_/Y vdd gnd OAI21X1
XFILL_1__9959_ vdd gnd FILL
XFILL_0__10200_ vdd gnd FILL
XFILL_0__11180_ vdd gnd FILL
XFILL_2__7703_ vdd gnd FILL
X_10587_ _10587_/A _10587_/B _10587_/C _10587_/Y vdd gnd OAI21X1
X_13375_ _13375_/A _13375_/B _13375_/C _13375_/Y vdd gnd OAI21X1
XFILL_0__10131_ vdd gnd FILL
XFILL_1__12470_ vdd gnd FILL
X_12326_ _12326_/A _12326_/B _12326_/Y vdd gnd NAND2X1
XFILL_2__7634_ vdd gnd FILL
XFILL_1__11421_ vdd gnd FILL
XFILL_2__10972_ vdd gnd FILL
XFILL_0__10062_ vdd gnd FILL
X_12257_ _12257_/A _12257_/B _12257_/C _12257_/Y vdd gnd OAI21X1
XFILL_1__14140_ vdd gnd FILL
XFILL_2__7565_ vdd gnd FILL
XFILL_1__11352_ vdd gnd FILL
X_11208_ _11208_/A _11208_/B _11208_/S _11208_/Y vdd gnd MUX2X1
X_12188_ _12188_/A _12188_/B _12188_/Y vdd gnd NOR2X1
XFILL_1__10303_ vdd gnd FILL
XFILL_1_BUFX2_insert18 vdd gnd FILL
XFILL_1__14071_ vdd gnd FILL
XFILL_0__13821_ vdd gnd FILL
XFILL_2__7496_ vdd gnd FILL
XFILL_1__11283_ vdd gnd FILL
X_11139_ _11139_/A _11139_/B _11139_/Y vdd gnd NAND2X1
XFILL_1__13022_ vdd gnd FILL
XFILL_1__10234_ vdd gnd FILL
XFILL_0__13752_ vdd gnd FILL
XFILL_0__10964_ vdd gnd FILL
XFILL_0__8250_ vdd gnd FILL
XFILL_0__12703_ vdd gnd FILL
XFILL_1__10165_ vdd gnd FILL
XFILL_0__7201_ vdd gnd FILL
XFILL_0__13683_ vdd gnd FILL
XFILL_0__8181_ vdd gnd FILL
XFILL_0__10895_ vdd gnd FILL
XFILL_2__8117_ vdd gnd FILL
XFILL_0__12634_ vdd gnd FILL
XFILL_0__7132_ vdd gnd FILL
XFILL_1__10096_ vdd gnd FILL
X_14829_ _14829_/A _14829_/B _14829_/Y vdd gnd NAND2X1
X_7760_ _7760_/A _7760_/B _7760_/Y vdd gnd NAND2X1
XFILL_2__10406_ vdd gnd FILL
XFILL_2__8048_ vdd gnd FILL
XFILL_1__13924_ vdd gnd FILL
XFILL_2__10337_ vdd gnd FILL
X_7691_ _7691_/A _7691_/B _7691_/Y vdd gnd NAND2X1
XFILL_0__14304_ vdd gnd FILL
XFILL_0__11516_ vdd gnd FILL
XFILL_1__13855_ vdd gnd FILL
X_9430_ _9430_/A _9430_/B _9430_/Y vdd gnd NAND2X1
XFILL_0__12496_ vdd gnd FILL
XFILL_2__10268_ vdd gnd FILL
XFILL_0__14235_ vdd gnd FILL
XFILL_1__12806_ vdd gnd FILL
XFILL_0__11447_ vdd gnd FILL
XFILL_1__10998_ vdd gnd FILL
XFILL_1__13786_ vdd gnd FILL
X_9361_ _9361_/A _9361_/B _9361_/Y vdd gnd NOR2X1
XFILL_2__10199_ vdd gnd FILL
XFILL_0_BUFX2_insert170 vdd gnd FILL
XFILL_1__12737_ vdd gnd FILL
XFILL_0_BUFX2_insert181 vdd gnd FILL
X_8312_ _8312_/A _8312_/B _8312_/C _8312_/Y vdd gnd NAND3X1
XFILL_0__11378_ vdd gnd FILL
XFILL_0_BUFX2_insert192 vdd gnd FILL
X_9292_ _9292_/A _9292_/B _9292_/C _9292_/Y vdd gnd OAI21X1
XFILL_0__13117_ vdd gnd FILL
XFILL_0__10329_ vdd gnd FILL
XFILL_1__12668_ vdd gnd FILL
XFILL_0__9704_ vdd gnd FILL
XFILL_0__14097_ vdd gnd FILL
X_8243_ _8243_/A _8243_/B _8243_/C _8243_/Y vdd gnd OAI21X1
XFILL_0__7896_ vdd gnd FILL
XFILL_1__14407_ vdd gnd FILL
XFILL_2__13958_ vdd gnd FILL
XFILL_0__13048_ vdd gnd FILL
XFILL_0__9635_ vdd gnd FILL
X_8174_ _8174_/A _8174_/B _8174_/C _8174_/Y vdd gnd NAND3X1
XFILL_1__14338_ vdd gnd FILL
XFILL_2__13889_ vdd gnd FILL
X_7125_ _7125_/A _7125_/B _7125_/C _7125_/Y vdd gnd OAI21X1
XFILL_0__9566_ vdd gnd FILL
XFILL_1__14269_ vdd gnd FILL
XFILL_1__7310_ vdd gnd FILL
XFILL_0__8517_ vdd gnd FILL
XFILL_0__9497_ vdd gnd FILL
XFILL_1__8290_ vdd gnd FILL
XFILL_1__7241_ vdd gnd FILL
XFILL_0__8448_ vdd gnd FILL
XFILL_1__7172_ vdd gnd FILL
XFILL_0__8379_ vdd gnd FILL
X_7958_ _7958_/D _7958_/CLK _7958_/Q vdd gnd DFFPOSX1
X_7889_ _7889_/A _7889_/B _7889_/C _7889_/Y vdd gnd OAI21X1
X_9628_ _9628_/A _9628_/B _9628_/C _9628_/Y vdd gnd OAI21X1
X_10510_ _10510_/A _10510_/B _10510_/C _10510_/Y vdd gnd AOI21X1
X_11490_ _11490_/A _11490_/B _11490_/Y vdd gnd NAND2X1
XBUFX2_insert10 BUFX2_insert10/A BUFX2_insert10/Y vdd gnd BUFX2
X_9559_ _9559_/A _9559_/B _9559_/C _9559_/Y vdd gnd OAI21X1
XBUFX2_insert21 BUFX2_insert21/A BUFX2_insert21/Y vdd gnd BUFX2
X_10441_ _10441_/A _10441_/B _10441_/C _10441_/Y vdd gnd OAI21X1
XFILL_1__9744_ vdd gnd FILL
X_13160_ _13160_/A _13160_/B _13160_/C _13160_/Y vdd gnd NAND3X1
X_10372_ _10372_/A _10372_/Y vdd gnd INVX1
XFILL_1__9675_ vdd gnd FILL
X_12111_ _12111_/A _12111_/B _12111_/C _12111_/Y vdd gnd OAI21X1
X_13091_ _13091_/A _13091_/B _13091_/Y vdd gnd NOR2X1
XFILL_1__8626_ vdd gnd FILL
X_12042_ _12042_/A _12042_/B _12042_/Y vdd gnd NAND2X1
XFILL_1__8557_ vdd gnd FILL
XFILL_1__7508_ vdd gnd FILL
XFILL_2__7281_ vdd gnd FILL
XFILL_1__8488_ vdd gnd FILL
XFILL_2_BUFX2_insert210 vdd gnd FILL
XFILL_1__7439_ vdd gnd FILL
X_13993_ _13993_/A _13993_/Y vdd gnd INVX1
XFILL_2_BUFX2_insert232 vdd gnd FILL
X_12944_ _12944_/A _12944_/B _12944_/Y vdd gnd NAND2X1
XFILL_2_BUFX2_insert265 vdd gnd FILL
XFILL_0__10680_ vdd gnd FILL
XFILL_2_BUFX2_insert287 vdd gnd FILL
XFILL_1__9109_ vdd gnd FILL
X_12875_ _12875_/A _12875_/B _12875_/C _12875_/Y vdd gnd NAND3X1
XFILL_1__11970_ vdd gnd FILL
X_14614_ _14614_/A _14614_/B _14614_/Y vdd gnd NAND2X1
X_11826_ _11826_/A _11826_/B _11826_/C _11826_/Y vdd gnd OAI21X1
XFILL_1__10921_ vdd gnd FILL
XFILL_0__12350_ vdd gnd FILL
X_14545_ _14545_/D _14545_/CLK _14545_/Q vdd gnd DFFPOSX1
XFILL_2__10122_ vdd gnd FILL
X_11757_ _11757_/A _11757_/Y vdd gnd INVX1
XBUFX2_insert220 BUFX2_insert220/A BUFX2_insert220/Y vdd gnd BUFX2
XFILL_0__11301_ vdd gnd FILL
XFILL_1__13640_ vdd gnd FILL
XBUFX2_insert231 BUFX2_insert231/A BUFX2_insert231/Y vdd gnd BUFX2
XFILL_1__10852_ vdd gnd FILL
XFILL_0__12281_ vdd gnd FILL
XBUFX2_insert242 BUFX2_insert242/A BUFX2_insert242/Y vdd gnd BUFX2
X_10708_ _10708_/D _10708_/CLK _10708_/Q vdd gnd DFFPOSX1
XBUFX2_insert253 BUFX2_insert253/A BUFX2_insert253/Y vdd gnd BUFX2
X_14476_ _14476_/A _14476_/Y vdd gnd INVX1
XBUFX2_insert264 BUFX2_insert264/A BUFX2_insert264/Y vdd gnd BUFX2
XFILL_2__10053_ vdd gnd FILL
X_11688_ _11688_/D _11688_/CLK _11688_/Q vdd gnd DFFPOSX1
XFILL_0__14020_ vdd gnd FILL
XBUFX2_insert275 BUFX2_insert275/A BUFX2_insert275/Y vdd gnd BUFX2
XFILL_1__13571_ vdd gnd FILL
XFILL_0__11232_ vdd gnd FILL
XBUFX2_insert286 BUFX2_insert286/A BUFX2_insert286/Y vdd gnd BUFX2
XFILL_1__10783_ vdd gnd FILL
XBUFX2_insert297 BUFX2_insert297/A BUFX2_insert297/Y vdd gnd BUFX2
X_13427_ _13427_/A _13427_/B _13427_/C _13427_/Y vdd gnd OAI21X1
X_10639_ _10639_/A _10639_/B _10639_/C _10639_/Y vdd gnd OAI21X1
XFILL_1__12522_ vdd gnd FILL
XFILL_0__11163_ vdd gnd FILL
XFILL_0__7750_ vdd gnd FILL
X_13358_ _13358_/A _13358_/B _13358_/Y vdd gnd NAND2X1
XFILL_0__10114_ vdd gnd FILL
XFILL_1__12453_ vdd gnd FILL
XFILL_0__11094_ vdd gnd FILL
X_12309_ _12309_/A _12309_/B _12309_/Y vdd gnd NAND2X1
XFILL_0__7681_ vdd gnd FILL
XFILL_2__7617_ vdd gnd FILL
XFILL_1__11404_ vdd gnd FILL
X_13289_ _13289_/A _13289_/B _13289_/C _13289_/Y vdd gnd OAI21X1
XFILL_0__10045_ vdd gnd FILL
XFILL_1__12384_ vdd gnd FILL
XFILL_2__10955_ vdd gnd FILL
XFILL_0__9420_ vdd gnd FILL
XFILL_2__7548_ vdd gnd FILL
XFILL_1__11335_ vdd gnd FILL
XFILL_1__14123_ vdd gnd FILL
XFILL_0__14853_ vdd gnd FILL
XFILL_2__10886_ vdd gnd FILL
XFILL_0__9351_ vdd gnd FILL
XFILL_1__14054_ vdd gnd FILL
XFILL_2__7479_ vdd gnd FILL
XFILL_1__11266_ vdd gnd FILL
XFILL_0__13804_ vdd gnd FILL
XFILL_0__14784_ vdd gnd FILL
XFILL_0__8302_ vdd gnd FILL
XFILL_0__11996_ vdd gnd FILL
XFILL_0__9282_ vdd gnd FILL
X_8930_ _8930_/A _8930_/B _8930_/C _8930_/D _8930_/Y vdd gnd AOI22X1
XFILL_1__13005_ vdd gnd FILL
XFILL_1__10217_ vdd gnd FILL
XFILL_0__13735_ vdd gnd FILL
XFILL_1__11197_ vdd gnd FILL
XFILL_0__10947_ vdd gnd FILL
XFILL_0__8233_ vdd gnd FILL
X_8861_ _8861_/D _8861_/CLK _8861_/Q vdd gnd DFFPOSX1
XFILL_1__10148_ vdd gnd FILL
XFILL_0__13666_ vdd gnd FILL
XFILL_2__12487_ vdd gnd FILL
XFILL_0__10878_ vdd gnd FILL
X_7812_ _7812_/A _7812_/B _7812_/Y vdd gnd NAND2X1
XFILL_0__8164_ vdd gnd FILL
X_8792_ _8792_/A _8792_/Y vdd gnd INVX1
XFILL_0__12617_ vdd gnd FILL
XFILL_1__10079_ vdd gnd FILL
XFILL_0__13597_ vdd gnd FILL
XFILL_0__7115_ vdd gnd FILL
X_7743_ _7743_/A _7743_/B _7743_/Y vdd gnd NAND2X1
XFILL_0__8095_ vdd gnd FILL
XFILL_1__13907_ vdd gnd FILL
XFILL_2__13108_ vdd gnd FILL
X_7674_ _7674_/A _7674_/B _7674_/C _7674_/D _7674_/Y vdd gnd AOI22X1
XFILL_1__13838_ vdd gnd FILL
XFILL_0__12479_ vdd gnd FILL
X_9413_ _9413_/A _9413_/Y vdd gnd INVX1
XFILL_0__14218_ vdd gnd FILL
XFILL_1__13769_ vdd gnd FILL
X_9344_ _9344_/A _9344_/Y vdd gnd INVX1
XFILL_0__8997_ vdd gnd FILL
XFILL_1__7790_ vdd gnd FILL
XFILL_0__14149_ vdd gnd FILL
X_9275_ _9275_/A _9275_/B _9275_/Y vdd gnd NAND2X1
X_8226_ _8226_/A _8226_/B _8226_/C _8226_/Y vdd gnd AOI21X1
XFILL_1__9460_ vdd gnd FILL
XFILL_0__7879_ vdd gnd FILL
XFILL_0__9618_ vdd gnd FILL
XFILL_1__8411_ vdd gnd FILL
X_8157_ _8157_/A _8157_/B _8157_/C _8157_/Y vdd gnd OAI21X1
XFILL_1__9391_ vdd gnd FILL
X_7108_ _7108_/A _7108_/Y vdd gnd INVX1
XFILL_0__9549_ vdd gnd FILL
XFILL_1__8342_ vdd gnd FILL
X_8088_ _8088_/A _8088_/B _8088_/Y vdd gnd NAND2X1
XFILL_1__8273_ vdd gnd FILL
XFILL_1__7224_ vdd gnd FILL
X_10990_ _10990_/A _10990_/B _10990_/Y vdd gnd NAND2X1
XFILL_1_BUFX2_insert206 vdd gnd FILL
XFILL_1__7155_ vdd gnd FILL
XFILL_1_BUFX2_insert217 vdd gnd FILL
XFILL_1_BUFX2_insert228 vdd gnd FILL
XFILL_1_BUFX2_insert239 vdd gnd FILL
X_12660_ _12660_/A _12660_/Y vdd gnd INVX1
XFILL_1__7086_ vdd gnd FILL
X_11611_ _11611_/A _11611_/B _11611_/C _11611_/Y vdd gnd OAI21X1
X_12591_ _12591_/D _12591_/CLK _12591_/Q vdd gnd DFFPOSX1
X_14330_ _14330_/A _14330_/B _14330_/Y vdd gnd NAND2X1
X_11542_ _11542_/A _11542_/B _11542_/Y vdd gnd NAND2X1
XFILL_0_CLKBUF1_insert387 vdd gnd FILL
X_14261_ _14261_/A _14261_/B _14261_/Y vdd gnd NAND2X1
X_11473_ _11473_/A _11473_/B _11473_/Y vdd gnd NOR2X1
X_13212_ _13212_/A _13212_/B _13212_/Y vdd gnd NAND2X1
X_10424_ _10424_/A _10424_/B _10424_/C _10424_/Y vdd gnd OAI21X1
XFILL_1__9727_ vdd gnd FILL
XFILL_2__8520_ vdd gnd FILL
X_14192_ _14192_/D _14192_/CLK _14192_/Q vdd gnd DFFPOSX1
X_13143_ _13143_/A _13143_/Y vdd gnd INVX1
X_10355_ _10355_/A _10355_/B _10355_/C _10355_/Y vdd gnd NAND3X1
XFILL_1__9658_ vdd gnd FILL
X_10286_ _10286_/A _10286_/B _10286_/Y vdd gnd NAND2X1
XFILL_1__8609_ vdd gnd FILL
X_13074_ _13074_/A _13074_/B _13074_/C _13074_/Y vdd gnd NAND3X1
XFILL_1__9589_ vdd gnd FILL
X_12025_ _12025_/A _12025_/B _12025_/Y vdd gnd NAND2X1
XFILL_1__11120_ vdd gnd FILL
XFILL_0__11850_ vdd gnd FILL
XFILL_2__12410_ vdd gnd FILL
XFILL_1__11051_ vdd gnd FILL
XFILL_0__10801_ vdd gnd FILL
XFILL_0__11781_ vdd gnd FILL
X_13976_ _13976_/A _13976_/B _13976_/C _13976_/Y vdd gnd OAI21X1
XFILL_1__10002_ vdd gnd FILL
XFILL_2__12341_ vdd gnd FILL
XFILL_0__13520_ vdd gnd FILL
X_12927_ _12927_/A _12927_/B _12927_/Y vdd gnd AND2X2
XFILL_1__14810_ vdd gnd FILL
XFILL_2__12272_ vdd gnd FILL
XFILL_0__10663_ vdd gnd FILL
XFILL_2__14011_ vdd gnd FILL
X_12858_ _12858_/A _12858_/Y vdd gnd INVX1
XFILL_0__12402_ vdd gnd FILL
XFILL_1__14741_ vdd gnd FILL
XFILL_1__11953_ vdd gnd FILL
XFILL_0__13382_ vdd gnd FILL
XFILL_0__10594_ vdd gnd FILL
X_11809_ _11809_/A _11809_/B _11809_/S _11809_/Y vdd gnd MUX2X1
XFILL_2__9905_ vdd gnd FILL
X_12789_ _12789_/A _12789_/Y vdd gnd INVX1
XFILL_0__12333_ vdd gnd FILL
XFILL_1__10904_ vdd gnd FILL
XFILL_1__14672_ vdd gnd FILL
XFILL_0__8920_ vdd gnd FILL
XFILL_1__11884_ vdd gnd FILL
X_14528_ _14528_/D _14528_/CLK _14528_/Q vdd gnd DFFPOSX1
XFILL_1__13623_ vdd gnd FILL
XFILL_0__12264_ vdd gnd FILL
XFILL_1__10835_ vdd gnd FILL
X_14459_ _14459_/A _14459_/B _14459_/Y vdd gnd NAND2X1
X_7390_ _7390_/A _7390_/B _7390_/Y vdd gnd AND2X2
XFILL_2__10036_ vdd gnd FILL
XFILL_0__14003_ vdd gnd FILL
XFILL_0__11215_ vdd gnd FILL
XFILL_1__13554_ vdd gnd FILL
XFILL_0__7802_ vdd gnd FILL
XFILL_0__12195_ vdd gnd FILL
XFILL_0__8782_ vdd gnd FILL
XFILL_2__14844_ vdd gnd FILL
XFILL_1__12505_ vdd gnd FILL
XFILL_2__9698_ vdd gnd FILL
XFILL_0__11146_ vdd gnd FILL
X_9060_ _9060_/A _9060_/B _9060_/Y vdd gnd NAND2X1
XFILL_0__7733_ vdd gnd FILL
XFILL_1__12436_ vdd gnd FILL
XFILL_0__11077_ vdd gnd FILL
X_8011_ _8011_/A _8011_/Y vdd gnd INVX1
XFILL_0__7664_ vdd gnd FILL
XFILL_0__10028_ vdd gnd FILL
XFILL_1__12367_ vdd gnd FILL
XFILL_0__9403_ vdd gnd FILL
XFILL_0__7595_ vdd gnd FILL
XFILL_1__11318_ vdd gnd FILL
XFILL_1__14106_ vdd gnd FILL
XFILL_0__14836_ vdd gnd FILL
XFILL_1__12298_ vdd gnd FILL
XFILL_0__9334_ vdd gnd FILL
X_9962_ _9962_/A _9962_/B _9962_/S _9962_/Y vdd gnd MUX2X1
XFILL_1__11249_ vdd gnd FILL
XFILL_1__14037_ vdd gnd FILL
XFILL_0__14767_ vdd gnd FILL
XFILL_0__11979_ vdd gnd FILL
XFILL_0__9265_ vdd gnd FILL
X_8913_ _8913_/D _8913_/CLK _8913_/Q vdd gnd DFFPOSX1
X_9893_ _9893_/A _9893_/B _9893_/C _9893_/D _9893_/Y vdd gnd AOI22X1
XFILL_0__13718_ vdd gnd FILL
XFILL_0__8216_ vdd gnd FILL
XFILL_0__14698_ vdd gnd FILL
XFILL_0__9196_ vdd gnd FILL
X_8844_ _8844_/D _8844_/CLK _8844_/Q vdd gnd DFFPOSX1
XFILL_0__13649_ vdd gnd FILL
XFILL_0__8147_ vdd gnd FILL
X_8775_ _8775_/A _8775_/B _8775_/Y vdd gnd AND2X2
XFILL_1__8960_ vdd gnd FILL
X_7726_ _7726_/A _7726_/B _7726_/C _7726_/Y vdd gnd OAI21X1
XFILL_0__8078_ vdd gnd FILL
XFILL_1__7911_ vdd gnd FILL
X_7657_ _7657_/A _7657_/B _7657_/Y vdd gnd NOR2X1
XFILL_1__7842_ vdd gnd FILL
X_7588_ _7588_/A _7588_/B _7588_/Y vdd gnd NAND2X1
X_9327_ _9327_/A _9327_/B _9327_/C _9327_/Y vdd gnd NAND3X1
XFILL256050x144150 vdd gnd FILL
XFILL_1__7773_ vdd gnd FILL
XFILL_1__9512_ vdd gnd FILL
X_9258_ _9258_/A _9258_/B _9258_/C _9258_/Y vdd gnd NAND3X1
X_10140_ _10140_/A _10140_/B _10140_/C _10140_/Y vdd gnd AOI21X1
XFILL_1__9443_ vdd gnd FILL
X_8209_ _8209_/A _8209_/B _8209_/Y vdd gnd NAND2X1
X_9189_ _9189_/A _9189_/B _9189_/C _9189_/Y vdd gnd NAND3X1
X_10071_ _10071_/A _10071_/Y vdd gnd INVX1
XFILL_1__9374_ vdd gnd FILL
XFILL_1__8325_ vdd gnd FILL
X_13830_ _13830_/A _13830_/B _13830_/Y vdd gnd OR2X2
XFILL_1__8256_ vdd gnd FILL
XFILL_1__7207_ vdd gnd FILL
X_13761_ _13761_/A _13761_/B _13761_/C _13761_/Y vdd gnd OAI21X1
X_10973_ _10973_/A _10973_/B _10973_/C _10973_/Y vdd gnd OAI21X1
XFILL_1__8187_ vdd gnd FILL
X_12712_ _12712_/A _12712_/Y vdd gnd INVX1
XFILL_1__7138_ vdd gnd FILL
X_13692_ _13692_/A _13692_/B _13692_/C _13692_/D _13692_/Y vdd gnd AOI22X1
X_12643_ _12643_/A _12643_/B _12643_/C _12643_/Y vdd gnd OAI21X1
XFILL257550x64950 vdd gnd FILL
X_12574_ _12574_/D _12574_/CLK _12574_/Q vdd gnd DFFPOSX1
XFILL_2__7882_ vdd gnd FILL
X_14313_ _14313_/A _14313_/B _14313_/Y vdd gnd OR2X2
X_11525_ _11525_/A _11525_/B _11525_/Y vdd gnd NAND2X1
XFILL_1__10620_ vdd gnd FILL
X_14244_ _14244_/A _14244_/B _14244_/Y vdd gnd NAND2X1
X_11456_ _11456_/A _11456_/B _11456_/Y vdd gnd NAND2X1
XFILL_0__11000_ vdd gnd FILL
XFILL_2__11910_ vdd gnd FILL
XFILL_1__10551_ vdd gnd FILL
X_10407_ _10407_/A _10407_/Y vdd gnd INVX1
XFILL_2__8503_ vdd gnd FILL
X_14175_ _14175_/D _14175_/CLK _14175_/Q vdd gnd DFFPOSX1
X_11387_ _11387_/A _11387_/B _11387_/Y vdd gnd NAND2X1
XFILL_2__11841_ vdd gnd FILL
XFILL_1__13270_ vdd gnd FILL
XFILL_1__10482_ vdd gnd FILL
X_13126_ _13126_/A _13126_/B _13126_/Y vdd gnd NOR2X1
X_10338_ _10338_/A _10338_/B _10338_/C _10338_/Y vdd gnd NAND3X1
XFILL_2__8434_ vdd gnd FILL
XFILL_1__12221_ vdd gnd FILL
XFILL_2__14560_ vdd gnd FILL
XFILL_2__11772_ vdd gnd FILL
XFILL_0__12951_ vdd gnd FILL
X_13057_ _13057_/A _13057_/B _13057_/C _13057_/Y vdd gnd OAI21X1
X_10269_ _10269_/A _10269_/B _10269_/C _10269_/Y vdd gnd NAND3X1
XFILL_1__12152_ vdd gnd FILL
XFILL_2__8365_ vdd gnd FILL
XFILL_0__11902_ vdd gnd FILL
X_12008_ _12008_/A _12008_/B _12008_/C _12008_/Y vdd gnd NAND3X1
XFILL_0__12882_ vdd gnd FILL
XFILL_0__7380_ vdd gnd FILL
XFILL_1__11103_ vdd gnd FILL
XFILL_0__14621_ vdd gnd FILL
XFILL_2__10654_ vdd gnd FILL
XFILL_1__12083_ vdd gnd FILL
XFILL_0__11833_ vdd gnd FILL
XFILL_2__8296_ vdd gnd FILL
XFILL_1__11034_ vdd gnd FILL
XFILL_2__10585_ vdd gnd FILL
XFILL_0__11764_ vdd gnd FILL
XFILL_0__9050_ vdd gnd FILL
X_13959_ _13959_/A _13959_/B _13959_/C _13959_/Y vdd gnd NAND3X1
XFILL_0__13503_ vdd gnd FILL
XFILL_0__8001_ vdd gnd FILL
XFILL_0__14483_ vdd gnd FILL
XFILL_0__11695_ vdd gnd FILL
XFILL_2__12255_ vdd gnd FILL
XFILL_0__10646_ vdd gnd FILL
XFILL_1__12985_ vdd gnd FILL
XFILL_2__11206_ vdd gnd FILL
X_8560_ _8560_/A _8560_/B _8560_/Y vdd gnd OR2X2
XFILL_1__14724_ vdd gnd FILL
XFILL_1__11936_ vdd gnd FILL
XFILL_2__12186_ vdd gnd FILL
XFILL_0__13365_ vdd gnd FILL
XFILL_0__10577_ vdd gnd FILL
X_7511_ _7511_/A _7511_/B _7511_/C _7511_/Y vdd gnd OAI21X1
XFILL_0__9952_ vdd gnd FILL
X_8491_ _8491_/A _8491_/B _8491_/Y vdd gnd NAND2X1
XFILL_0__12316_ vdd gnd FILL
XFILL_1__14655_ vdd gnd FILL
XFILL_1__11867_ vdd gnd FILL
XFILL_0__13296_ vdd gnd FILL
X_7442_ _7442_/A _7442_/B _7442_/C _7442_/Y vdd gnd NAND3X1
XFILL_0__9883_ vdd gnd FILL
XFILL_1__13606_ vdd gnd FILL
XFILL_0__12247_ vdd gnd FILL
XFILL_1__10818_ vdd gnd FILL
XFILL_1__14586_ vdd gnd FILL
XFILL_0__8834_ vdd gnd FILL
XFILL_1__11798_ vdd gnd FILL
X_7373_ _7373_/A _7373_/B _7373_/Y vdd gnd AND2X2
XFILL_1__13537_ vdd gnd FILL
XFILL_0__12178_ vdd gnd FILL
X_9112_ _9112_/A _9112_/B _9112_/Y vdd gnd NAND2X1
XFILL_0__8765_ vdd gnd FILL
XFILL_2__14827_ vdd gnd FILL
XFILL_2_CLKBUF1_insert60 vdd gnd FILL
XFILL_0__11129_ vdd gnd FILL
XFILL_2_CLKBUF1_insert82 vdd gnd FILL
X_9043_ _9043_/A _9043_/B _9043_/C _9043_/Y vdd gnd OAI21X1
XFILL_0__7716_ vdd gnd FILL
XFILL_0__8696_ vdd gnd FILL
XFILL_2__14758_ vdd gnd FILL
XFILL_1__12419_ vdd gnd FILL
XFILL_1__13399_ vdd gnd FILL
XFILL_0__7647_ vdd gnd FILL
XFILL_2__14689_ vdd gnd FILL
XFILL_0__7578_ vdd gnd FILL
XFILL_0__14819_ vdd gnd FILL
XFILL_0__9317_ vdd gnd FILL
XFILL_0_BUFX2_insert20 vdd gnd FILL
XFILL_1__8110_ vdd gnd FILL
X_9945_ _9945_/A _9945_/B _9945_/Y vdd gnd NAND2X1
XFILL_1__9090_ vdd gnd FILL
XFILL_0__9248_ vdd gnd FILL
XFILL_1__8041_ vdd gnd FILL
X_9876_ _9876_/A _9876_/B _9876_/Y vdd gnd NAND2X1
XFILL_0__9179_ vdd gnd FILL
X_8827_ _8827_/A _8827_/B _8827_/C _8827_/Y vdd gnd OAI21X1
XFILL_1__9992_ vdd gnd FILL
X_8758_ _8758_/A _8758_/B _8758_/Y vdd gnd NOR2X1
XFILL_1__8943_ vdd gnd FILL
X_7709_ _7709_/A _7709_/B _7709_/C _7709_/Y vdd gnd OAI21X1
X_8689_ _8689_/A _8689_/B _8689_/C _8689_/Y vdd gnd OAI21X1
X_11310_ _11310_/A _11310_/B _11310_/C _11310_/Y vdd gnd OAI21X1
XFILL_1__7825_ vdd gnd FILL
X_12290_ _12290_/A _12290_/B _12290_/Y vdd gnd NAND2X1
X_11241_ _11241_/A _11241_/B _11241_/C _11241_/Y vdd gnd NAND3X1
XFILL_1__7756_ vdd gnd FILL
X_11172_ _11172_/A _11172_/B _11172_/C _11172_/Y vdd gnd OAI21X1
XFILL_1__7687_ vdd gnd FILL
X_10123_ _10123_/A _10123_/Y vdd gnd INVX1
XFILL_1__9426_ vdd gnd FILL
X_10054_ _10054_/A _10054_/B _10054_/Y vdd gnd NAND2X1
XFILL_1__9357_ vdd gnd FILL
XFILL_2__8150_ vdd gnd FILL
X_14862_ _14862_/A _14862_/B _14862_/C _14862_/Y vdd gnd OAI21X1
XFILL_1__8308_ vdd gnd FILL
XFILL_1__9288_ vdd gnd FILL
XFILL_2__8081_ vdd gnd FILL
X_13813_ _13813_/A _13813_/B _13813_/Y vdd gnd NAND2X1
X_14793_ _14793_/A _14793_/B _14793_/Y vdd gnd AND2X2
XFILL_1__8239_ vdd gnd FILL
XFILL_2__10370_ vdd gnd FILL
X_13744_ _13744_/A _13744_/Y vdd gnd INVX1
X_10956_ _10956_/A _10956_/B _10956_/Y vdd gnd NAND2X1
XFILL_0__10500_ vdd gnd FILL
XFILL_0__11480_ vdd gnd FILL
X_13675_ _13675_/A _13675_/B _13675_/C _13675_/Y vdd gnd OAI21X1
X_10887_ _10887_/A _10887_/B _10887_/S _10887_/Y vdd gnd MUX2X1
XFILL_2__8983_ vdd gnd FILL
XFILL_0__10431_ vdd gnd FILL
XFILL_1__12770_ vdd gnd FILL
X_12626_ _12626_/A _12626_/B _12626_/C _12626_/Y vdd gnd AOI21X1
XFILL_0__13150_ vdd gnd FILL
XFILL_1__11721_ vdd gnd FILL
XFILL_0__10362_ vdd gnd FILL
X_12557_ _12557_/D _12557_/CLK _12557_/Q vdd gnd DFFPOSX1
XFILL_0__12101_ vdd gnd FILL
XFILL_2__7865_ vdd gnd FILL
XFILL_1__14440_ vdd gnd FILL
XFILL_0__13081_ vdd gnd FILL
XFILL_0__10293_ vdd gnd FILL
X_11508_ _11508_/A _11508_/B _11508_/Y vdd gnd NAND2X1
X_12488_ _12488_/A _12488_/Y vdd gnd INVX1
XFILL_1__10603_ vdd gnd FILL
XFILL_0__12032_ vdd gnd FILL
XFILL_2__7796_ vdd gnd FILL
XFILL_1__14371_ vdd gnd FILL
XFILL_1__11583_ vdd gnd FILL
X_14227_ _14227_/A _14227_/B _14227_/C _14227_/Y vdd gnd OAI21X1
X_11439_ _11439_/A _11439_/B _11439_/Y vdd gnd NAND2X1
XFILL_1__10534_ vdd gnd FILL
XFILL_1__13322_ vdd gnd FILL
XFILL_0__8550_ vdd gnd FILL
X_14158_ _14158_/A _14158_/B _14158_/C _14158_/Y vdd gnd OAI21X1
XFILL_2__14612_ vdd gnd FILL
XFILL_2__11824_ vdd gnd FILL
XFILL_1__10465_ vdd gnd FILL
XFILL_1__13253_ vdd gnd FILL
X_13109_ _13109_/A _13109_/Y vdd gnd INVX1
XFILL_0__7501_ vdd gnd FILL
XFILL_0__13983_ vdd gnd FILL
XFILL_0__8481_ vdd gnd FILL
XFILL_2__8417_ vdd gnd FILL
X_14089_ _14089_/A _14089_/B _14089_/Y vdd gnd NAND2X1
XFILL_1__12204_ vdd gnd FILL
XFILL_1__13184_ vdd gnd FILL
XFILL_2__11755_ vdd gnd FILL
XFILL_0__12934_ vdd gnd FILL
XFILL_1__10396_ vdd gnd FILL
XFILL_0__7432_ vdd gnd FILL
XFILL_2__8348_ vdd gnd FILL
XFILL_1__12135_ vdd gnd FILL
XFILL_0__12865_ vdd gnd FILL
XFILL_0__7363_ vdd gnd FILL
XFILL_2__13425_ vdd gnd FILL
XFILL_0__14604_ vdd gnd FILL
XFILL_2__10637_ vdd gnd FILL
X_7991_ _7991_/D _7991_/CLK _7991_/Q vdd gnd DFFPOSX1
XFILL_2__8279_ vdd gnd FILL
XFILL_1__12066_ vdd gnd FILL
XFILL_0__9102_ vdd gnd FILL
XFILL_0__11816_ vdd gnd FILL
XFILL_0__12796_ vdd gnd FILL
X_9730_ _9730_/A _9730_/B _9730_/C _9730_/Y vdd gnd OAI21X1
XFILL_0__7294_ vdd gnd FILL
XFILL_1__11017_ vdd gnd FILL
XFILL_2__10568_ vdd gnd FILL
XFILL_0__9033_ vdd gnd FILL
XFILL_0__11747_ vdd gnd FILL
X_9661_ _9661_/A _9661_/B _9661_/Y vdd gnd NAND2X1
XFILL_2__10499_ vdd gnd FILL
XFILL_0__14466_ vdd gnd FILL
X_8612_ _8612_/A _8612_/B _8612_/Y vdd gnd NOR2X1
X_9592_ _9592_/A _9592_/B _9592_/C _9592_/Y vdd gnd AOI21X1
XFILL_0__10629_ vdd gnd FILL
XFILL_0__13417_ vdd gnd FILL
XFILL_1__12968_ vdd gnd FILL
XFILL_0__14397_ vdd gnd FILL
X_8543_ _8543_/A _8543_/B _8543_/C _8543_/Y vdd gnd OAI21X1
XFILL_1__14707_ vdd gnd FILL
XFILL_1__11919_ vdd gnd FILL
XFILL_0__13348_ vdd gnd FILL
XFILL_0__9935_ vdd gnd FILL
XFILL_1__12899_ vdd gnd FILL
X_8474_ _8474_/A _8474_/B _8474_/C _8474_/D _8474_/Y vdd gnd AOI22X1
XFILL_1__14638_ vdd gnd FILL
XFILL_0__13279_ vdd gnd FILL
X_7425_ _7425_/A _7425_/B _7425_/Y vdd gnd NAND2X1
XFILL_0__9866_ vdd gnd FILL
XFILL_1__14569_ vdd gnd FILL
XFILL_1__7610_ vdd gnd FILL
XFILL_0__8817_ vdd gnd FILL
X_7356_ _7356_/A _7356_/B _7356_/Y vdd gnd OR2X2
XFILL_1__8590_ vdd gnd FILL
XFILL_1__7541_ vdd gnd FILL
XFILL_0__8748_ vdd gnd FILL
X_7287_ _7287_/A _7287_/B _7287_/C _7287_/Y vdd gnd NAND3X1
X_9026_ _9026_/A _9026_/B _9026_/S _9026_/Y vdd gnd MUX2X1
XFILL_1__7472_ vdd gnd FILL
XFILL_0__8679_ vdd gnd FILL
XFILL_1__9211_ vdd gnd FILL
XFILL_1__9142_ vdd gnd FILL
XFILL_1__9073_ vdd gnd FILL
X_9928_ _9928_/A _9928_/B _9928_/C _9928_/Y vdd gnd OAI21X1
X_10810_ _10810_/A _10810_/Y vdd gnd INVX1
XFILL_1__8024_ vdd gnd FILL
X_11790_ _11790_/A _11790_/Y vdd gnd INVX1
X_9859_ _9859_/A _9859_/Y vdd gnd INVX1
X_10741_ _10741_/D _10741_/CLK _10741_/Q vdd gnd DFFPOSX1
X_13460_ _13460_/D _13460_/CLK _13460_/Q vdd gnd DFFPOSX1
X_10672_ _10672_/A _10672_/B _10672_/Y vdd gnd NAND2X1
XFILL_1__9975_ vdd gnd FILL
X_12411_ _12411_/A _12411_/B _12411_/Y vdd gnd OR2X2
XFILL_1__8926_ vdd gnd FILL
X_13391_ _13391_/A _13391_/B _13391_/C _13391_/Y vdd gnd OAI21X1
X_12342_ _12342_/A _12342_/B _12342_/Y vdd gnd NAND2X1
XFILL_1__7808_ vdd gnd FILL
X_12273_ _12273_/A _12273_/B _12273_/C _12273_/Y vdd gnd OAI21X1
XFILL_1__8788_ vdd gnd FILL
X_14012_ _14012_/A _14012_/B _14012_/C _14012_/Y vdd gnd OAI21X1
X_11224_ _11224_/A _11224_/B _11224_/C _11224_/D _11224_/Y vdd gnd AOI22X1
XFILL_1__7739_ vdd gnd FILL
X_11155_ _11155_/A _11155_/B _11155_/Y vdd gnd NAND2X1
XFILL_1__10250_ vdd gnd FILL
XFILL_0__10980_ vdd gnd FILL
X_10106_ _10106_/A _10106_/B _10106_/C _10106_/Y vdd gnd NAND3X1
XFILL_1__9409_ vdd gnd FILL
X_11086_ _11086_/A _11086_/B _11086_/Y vdd gnd AND2X2
XFILL257250x86550 vdd gnd FILL
XFILL_1__10181_ vdd gnd FILL
X_10037_ _10037_/A _10037_/B _10037_/C _10037_/Y vdd gnd OAI21X1
X_14914_ _14914_/A _14914_/Y vdd gnd BUFX2
XFILL_0__12650_ vdd gnd FILL
XFILL_2__13210_ vdd gnd FILL
X_14845_ _14845_/A _14845_/B _14845_/C _14845_/Y vdd gnd OAI21X1
XFILL_2__8064_ vdd gnd FILL
XFILL_1__13940_ vdd gnd FILL
XFILL_0__11601_ vdd gnd FILL
X_14776_ _14776_/A _14776_/B _14776_/C _14776_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert1 vdd gnd FILL
XFILL_2__13141_ vdd gnd FILL
X_11988_ _11988_/A _11988_/B _11988_/C _11988_/Y vdd gnd AOI21X1
XFILL_2__10353_ vdd gnd FILL
XFILL_0__14320_ vdd gnd FILL
XFILL_0__11532_ vdd gnd FILL
XFILL_1__13871_ vdd gnd FILL
X_13727_ _13727_/A _13727_/B _13727_/Y vdd gnd NAND2X1
X_10939_ _10939_/A _10939_/B _10939_/Y vdd gnd NOR2X1
XFILL_0__14251_ vdd gnd FILL
XFILL_1__12822_ vdd gnd FILL
XFILL_2__13072_ vdd gnd FILL
XFILL_2__10284_ vdd gnd FILL
XFILL_0__11463_ vdd gnd FILL
X_13658_ _13658_/A _13658_/B _13658_/C _13658_/D _13658_/Y vdd gnd AOI22X1
XFILL_0__13202_ vdd gnd FILL
XFILL_0__10414_ vdd gnd FILL
XFILL_1__12753_ vdd gnd FILL
XFILL_0_BUFX2_insert330 vdd gnd FILL
XFILL_0_BUFX2_insert341 vdd gnd FILL
X_12609_ _12609_/D _12609_/CLK _12609_/Q vdd gnd DFFPOSX1
XFILL_0__11394_ vdd gnd FILL
XFILL_0_BUFX2_insert352 vdd gnd FILL
X_13589_ _13589_/A _13589_/Y vdd gnd INVX1
XFILL_0__13133_ vdd gnd FILL
XFILL_0_BUFX2_insert363 vdd gnd FILL
XFILL_1__11704_ vdd gnd FILL
XFILL_0__10345_ vdd gnd FILL
XFILL_0_BUFX2_insert374 vdd gnd FILL
XFILL_0__9720_ vdd gnd FILL
XFILL_1__12684_ vdd gnd FILL
XFILL_1__14423_ vdd gnd FILL
XFILL_0__13064_ vdd gnd FILL
XFILL_0__10276_ vdd gnd FILL
X_7210_ _7210_/A _7210_/B _7210_/S _7210_/Y vdd gnd MUX2X1
XFILL_0__9651_ vdd gnd FILL
X_8190_ _8190_/A _8190_/Y vdd gnd INVX2
XFILL_0__12015_ vdd gnd FILL
XFILL_2__7779_ vdd gnd FILL
XFILL_1__14354_ vdd gnd FILL
XFILL_0__8602_ vdd gnd FILL
XFILL_1__11566_ vdd gnd FILL
X_7141_ _7141_/A _7141_/Y vdd gnd INVX1
XFILL_0__9582_ vdd gnd FILL
XFILL_1__13305_ vdd gnd FILL
XFILL_1__10517_ vdd gnd FILL
XFILL_1__14285_ vdd gnd FILL
XFILL_0__8533_ vdd gnd FILL
XFILL_1__11497_ vdd gnd FILL
X_7072_ _7072_/A _7072_/Y vdd gnd INVX1
XFILL_2__11807_ vdd gnd FILL
XFILL_1__13236_ vdd gnd FILL
XFILL_1__10448_ vdd gnd FILL
XFILL_0__13966_ vdd gnd FILL
XFILL_0__8464_ vdd gnd FILL
XFILL256950x252150 vdd gnd FILL
XFILL_2__11738_ vdd gnd FILL
XFILL_1__13167_ vdd gnd FILL
XFILL257550x237750 vdd gnd FILL
XFILL_1__10379_ vdd gnd FILL
XFILL_0__12917_ vdd gnd FILL
XFILL_0__7415_ vdd gnd FILL
XFILL_0__13897_ vdd gnd FILL
XFILL_0__8395_ vdd gnd FILL
XFILL_1__12118_ vdd gnd FILL
XFILL_0__12848_ vdd gnd FILL
XFILL_1__13098_ vdd gnd FILL
XFILL_0__7346_ vdd gnd FILL
XFILL_2__13408_ vdd gnd FILL
X_7974_ _7974_/D _7974_/CLK _7974_/Q vdd gnd DFFPOSX1
XFILL_1__12049_ vdd gnd FILL
X_9713_ _9713_/A _9713_/B _9713_/C _9713_/Y vdd gnd OAI21X1
XFILL_0__12779_ vdd gnd FILL
XFILL_0__7277_ vdd gnd FILL
XFILL_2__13339_ vdd gnd FILL
XFILL_0__9016_ vdd gnd FILL
X_9644_ _9644_/A _9644_/Y vdd gnd INVX1
XFILL_0__14449_ vdd gnd FILL
X_9575_ _9575_/A _9575_/B _9575_/C _9575_/Y vdd gnd OAI21X1
XFILL_1__9760_ vdd gnd FILL
X_8526_ _8526_/A _8526_/B _8526_/Y vdd gnd NOR2X1
XFILL_1__8711_ vdd gnd FILL
XFILL_0__9918_ vdd gnd FILL
XFILL_1__9691_ vdd gnd FILL
X_8457_ _8457_/A _8457_/B _8457_/C _8457_/Y vdd gnd OAI21X1
X_7408_ _7408_/A _7408_/B _7408_/C _7408_/Y vdd gnd AOI21X1
XFILL_1__8642_ vdd gnd FILL
XFILL_0__9849_ vdd gnd FILL
X_8388_ _8388_/A _8388_/B _8388_/Y vdd gnd NAND2X1
X_7339_ _7339_/A _7339_/B _7339_/C _7339_/Y vdd gnd NAND3X1
XFILL_1__8573_ vdd gnd FILL
XFILL_1__7524_ vdd gnd FILL
X_9009_ _9009_/A _9009_/B _9009_/S _9009_/Y vdd gnd MUX2X1
XFILL_1__7455_ vdd gnd FILL
XFILL257550x147750 vdd gnd FILL
X_12960_ _12960_/A _12960_/B _12960_/Y vdd gnd NAND2X1
XFILL_1__7386_ vdd gnd FILL
X_11911_ _11911_/A _11911_/B _11911_/C _11911_/Y vdd gnd NAND3X1
XFILL_1__9125_ vdd gnd FILL
XFILL257250x18150 vdd gnd FILL
X_12891_ _12891_/A _12891_/B _12891_/C _12891_/Y vdd gnd AOI21X1
X_14630_ _14630_/A _14630_/B _14630_/C _14630_/Y vdd gnd OAI21X1
X_11842_ _11842_/A _11842_/Y vdd gnd INVX1
XFILL_1__9056_ vdd gnd FILL
X_14561_ _14561_/A _14561_/Y vdd gnd INVX1
XFILL_1__8007_ vdd gnd FILL
X_11773_ _11773_/A _11773_/B _11773_/C _11773_/Y vdd gnd OAI21X1
XFILL257550x190950 vdd gnd FILL
X_13512_ _13512_/A _13512_/B _13512_/C _13512_/Y vdd gnd AOI21X1
X_10724_ _10724_/D _10724_/CLK _10724_/Q vdd gnd DFFPOSX1
XFILL_2__8820_ vdd gnd FILL
X_14492_ _14492_/A _14492_/B _14492_/C _14492_/Y vdd gnd OAI21X1
XFILL257250x61350 vdd gnd FILL
X_13443_ _13443_/D _13443_/CLK _13443_/Q vdd gnd DFFPOSX1
X_10655_ _10655_/A _10655_/B _10655_/C _10655_/Y vdd gnd OAI21X1
XFILL_2__8751_ vdd gnd FILL
XFILL_1__9958_ vdd gnd FILL
X_13374_ _13374_/A _13374_/B _13374_/Y vdd gnd NAND2X1
X_10586_ _10586_/A _10586_/B _10586_/Y vdd gnd AND2X2
XFILL_0__10130_ vdd gnd FILL
XFILL_2__8682_ vdd gnd FILL
XFILL_1__9889_ vdd gnd FILL
X_12325_ _12325_/A _12325_/B _12325_/Y vdd gnd NAND2X1
XFILL_1__11420_ vdd gnd FILL
XFILL_0__10061_ vdd gnd FILL
X_12256_ _12256_/A _12256_/B _12256_/Y vdd gnd OR2X2
XFILL_2__12710_ vdd gnd FILL
XFILL_1__11351_ vdd gnd FILL
X_11207_ _11207_/A _11207_/B _11207_/C _11207_/Y vdd gnd OAI21X1
XFILL_2__9303_ vdd gnd FILL
X_12187_ _12187_/A _12187_/B _12187_/Y vdd gnd NAND2X1
XFILL_1__10302_ vdd gnd FILL
XFILL_1_BUFX2_insert19 vdd gnd FILL
XFILL_1__14070_ vdd gnd FILL
XFILL_0__13820_ vdd gnd FILL
XFILL_1__11282_ vdd gnd FILL
X_11138_ _11138_/A _11138_/B _11138_/C _11138_/Y vdd gnd NAND3X1
XFILL_2__9234_ vdd gnd FILL
XFILL_1__10233_ vdd gnd FILL
XFILL_1__13021_ vdd gnd FILL
XFILL_0__13751_ vdd gnd FILL
XFILL_0__10963_ vdd gnd FILL
X_11069_ _11069_/A _11069_/B _11069_/Y vdd gnd AND2X2
XFILL_2__14311_ vdd gnd FILL
XFILL_1__10164_ vdd gnd FILL
XFILL_0__12702_ vdd gnd FILL
XFILL_0__7200_ vdd gnd FILL
XFILL_0__10894_ vdd gnd FILL
XFILL_0__13682_ vdd gnd FILL
XFILL_0__8180_ vdd gnd FILL
XFILL_2__14242_ vdd gnd FILL
XFILL_0__12633_ vdd gnd FILL
XFILL_1__10095_ vdd gnd FILL
XFILL_0__7131_ vdd gnd FILL
X_14828_ _14828_/A _14828_/B _14828_/C _14828_/Y vdd gnd OAI21X1
XFILL_1__13923_ vdd gnd FILL
XFILL_2__13124_ vdd gnd FILL
X_14759_ _14759_/A _14759_/B _14759_/Y vdd gnd NOR2X1
X_7690_ _7690_/A _7690_/B _7690_/Y vdd gnd NAND2X1
XFILL_0__14303_ vdd gnd FILL
XFILL_1__13854_ vdd gnd FILL
XFILL_0__11515_ vdd gnd FILL
XFILL_0__12495_ vdd gnd FILL
XFILL_2__13055_ vdd gnd FILL
XFILL_1__12805_ vdd gnd FILL
XFILL_0__14234_ vdd gnd FILL
XFILL_0__11446_ vdd gnd FILL
XFILL_1__13785_ vdd gnd FILL
XFILL_1__10997_ vdd gnd FILL
X_9360_ _9360_/A _9360_/B _9360_/S _9360_/Y vdd gnd MUX2X1
XFILL_0_BUFX2_insert160 vdd gnd FILL
XFILL_1__12736_ vdd gnd FILL
XFILL257550x212550 vdd gnd FILL
XFILL_0_BUFX2_insert171 vdd gnd FILL
XFILL_0__11377_ vdd gnd FILL
X_8311_ _8311_/A _8311_/B _8311_/C _8311_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert182 vdd gnd FILL
X_9291_ _9291_/A _9291_/B _9291_/Y vdd gnd NAND2X1
XFILL_0_BUFX2_insert193 vdd gnd FILL
XFILL_0__13116_ vdd gnd FILL
XFILL_0__10328_ vdd gnd FILL
XFILL_0__14096_ vdd gnd FILL
XFILL_1__12667_ vdd gnd FILL
XFILL_0__9703_ vdd gnd FILL
X_8242_ _8242_/A _8242_/B _8242_/C _8242_/Y vdd gnd AOI21X1
XFILL_0__7895_ vdd gnd FILL
XFILL_1__14406_ vdd gnd FILL
XFILL_0__13047_ vdd gnd FILL
XFILL_0__10259_ vdd gnd FILL
XFILL_0__9634_ vdd gnd FILL
X_8173_ _8173_/A _8173_/B _8173_/C _8173_/Y vdd gnd OAI21X1
XFILL_1__14337_ vdd gnd FILL
XFILL_1__11549_ vdd gnd FILL
X_7124_ _7124_/A _7124_/B _7124_/Y vdd gnd NOR2X1
XFILL_0__9565_ vdd gnd FILL
XFILL_1__14268_ vdd gnd FILL
XFILL_0__8516_ vdd gnd FILL
XFILL_0__9496_ vdd gnd FILL
XFILL_1__13219_ vdd gnd FILL
XFILL_0__13949_ vdd gnd FILL
XFILL_1__7240_ vdd gnd FILL
XFILL_0__8447_ vdd gnd FILL
XFILL_1__7171_ vdd gnd FILL
XFILL_0__8378_ vdd gnd FILL
XFILL_0__7329_ vdd gnd FILL
X_7957_ _7957_/D _7957_/CLK _7957_/Q vdd gnd DFFPOSX1
X_7888_ _7888_/A _7888_/B _7888_/Y vdd gnd NAND2X1
X_9627_ _9627_/A _9627_/B _9627_/Y vdd gnd NAND2X1
X_9558_ _9558_/A _9558_/B _9558_/C _9558_/Y vdd gnd OAI21X1
XBUFX2_insert11 BUFX2_insert11/A BUFX2_insert11/Y vdd gnd BUFX2
XFILL257550x122550 vdd gnd FILL
XBUFX2_insert22 BUFX2_insert22/A BUFX2_insert22/Y vdd gnd BUFX2
X_10440_ _10440_/A _10440_/B _10440_/Y vdd gnd NOR2X1
X_8509_ _8509_/A _8509_/B _8509_/C _8509_/Y vdd gnd AOI21X1
XFILL_1__9743_ vdd gnd FILL
X_9489_ _9489_/A _9489_/B _9489_/Y vdd gnd NOR2X1
X_10371_ _10371_/A _10371_/Y vdd gnd INVX1
XFILL_1__9674_ vdd gnd FILL
X_12110_ _12110_/A _12110_/B _12110_/Y vdd gnd NAND2X1
X_13090_ _13090_/A _13090_/B _13090_/Y vdd gnd NAND2X1
XFILL_1__8625_ vdd gnd FILL
X_12041_ _12041_/A _12041_/Y vdd gnd INVX1
XFILL_1__8556_ vdd gnd FILL
XFILL_1__7507_ vdd gnd FILL
XFILL_1__8487_ vdd gnd FILL
X_13992_ _13992_/A _13992_/B _13992_/C _13992_/Y vdd gnd NOR3X1
XFILL_1__7438_ vdd gnd FILL
XFILL_2_BUFX2_insert222 vdd gnd FILL
X_12943_ _12943_/A _12943_/B _12943_/C _12943_/Y vdd gnd NAND3X1
XFILL_2_BUFX2_insert244 vdd gnd FILL
XFILL_1__7369_ vdd gnd FILL
XFILL_2_BUFX2_insert277 vdd gnd FILL
XFILL_1__9108_ vdd gnd FILL
X_12874_ _12874_/A _12874_/B _12874_/Y vdd gnd NAND2X1
XFILL_2_BUFX2_insert299 vdd gnd FILL
X_14613_ _14613_/A _14613_/Y vdd gnd INVX1
X_11825_ _11825_/A _11825_/B _11825_/Y vdd gnd NAND2X1
XFILL_1__9039_ vdd gnd FILL
XFILL_2__9921_ vdd gnd FILL
XFILL_2__11170_ vdd gnd FILL
XFILL_1__10920_ vdd gnd FILL
X_14544_ _14544_/D _14544_/CLK _14544_/Q vdd gnd DFFPOSX1
X_11756_ _11756_/A _11756_/B _11756_/C _11756_/Y vdd gnd OAI21X1
XFILL_0__11300_ vdd gnd FILL
XBUFX2_insert210 BUFX2_insert210/A BUFX2_insert210/Y vdd gnd BUFX2
XFILL_2__9852_ vdd gnd FILL
XBUFX2_insert221 BUFX2_insert221/A BUFX2_insert221/Y vdd gnd BUFX2
XFILL_0__12280_ vdd gnd FILL
XFILL_1__10851_ vdd gnd FILL
X_10707_ _10707_/D _10707_/CLK _10707_/Q vdd gnd DFFPOSX1
XBUFX2_insert232 BUFX2_insert232/A BUFX2_insert232/Y vdd gnd BUFX2
XBUFX2_insert243 BUFX2_insert243/A BUFX2_insert243/Y vdd gnd BUFX2
X_14475_ _14475_/A _14475_/B _14475_/C _14475_/Y vdd gnd OAI21X1
XBUFX2_insert254 BUFX2_insert254/A BUFX2_insert254/Y vdd gnd BUFX2
XFILL_2__8803_ vdd gnd FILL
X_11687_ _11687_/D _11687_/CLK _11687_/Q vdd gnd DFFPOSX1
XFILL_0__11231_ vdd gnd FILL
XBUFX2_insert265 BUFX2_insert265/A BUFX2_insert265/Y vdd gnd BUFX2
XFILL_1__13570_ vdd gnd FILL
XBUFX2_insert276 BUFX2_insert276/A BUFX2_insert276/Y vdd gnd BUFX2
XFILL_1__10782_ vdd gnd FILL
X_13426_ _13426_/A _13426_/B _13426_/Y vdd gnd NAND2X1
X_10638_ _10638_/A _10638_/B _10638_/Y vdd gnd NAND2X1
XBUFX2_insert287 BUFX2_insert287/A BUFX2_insert287/Y vdd gnd BUFX2
XBUFX2_insert298 BUFX2_insert298/A BUFX2_insert298/Y vdd gnd BUFX2
XFILL_2__14860_ vdd gnd FILL
XFILL_2__8734_ vdd gnd FILL
XFILL_1__12521_ vdd gnd FILL
XFILL_0__11162_ vdd gnd FILL
X_13357_ _13357_/A _13357_/B _13357_/C _13357_/Y vdd gnd OAI21X1
X_10569_ _10569_/A _10569_/B _10569_/C _10569_/Y vdd gnd NAND3X1
XFILL_2__13811_ vdd gnd FILL
XFILL_0__10113_ vdd gnd FILL
XFILL_2__8665_ vdd gnd FILL
XFILL_2__14791_ vdd gnd FILL
XFILL_1__12452_ vdd gnd FILL
XFILL_0__11093_ vdd gnd FILL
X_12308_ _12308_/A _12308_/B _12308_/Y vdd gnd NOR2X1
XFILL_0__7680_ vdd gnd FILL
X_13288_ _13288_/A _13288_/B _13288_/Y vdd gnd NAND2X1
XFILL_1__11403_ vdd gnd FILL
XFILL_2__13742_ vdd gnd FILL
XFILL_0__10044_ vdd gnd FILL
XFILL_2__8596_ vdd gnd FILL
XFILL_1__12383_ vdd gnd FILL
X_12239_ _12239_/A _12239_/B _12239_/C _12239_/Y vdd gnd OAI21X1
XFILL_1__14122_ vdd gnd FILL
XFILL_1__11334_ vdd gnd FILL
XFILL_0__14852_ vdd gnd FILL
XFILL_0__9350_ vdd gnd FILL
XFILL_2__12624_ vdd gnd FILL
XFILL_1__14053_ vdd gnd FILL
XFILL_0__13803_ vdd gnd FILL
XFILL_0__8301_ vdd gnd FILL
XFILL_1__11265_ vdd gnd FILL
XFILL_0__14783_ vdd gnd FILL
XFILL_0__9281_ vdd gnd FILL
XFILL_2__9217_ vdd gnd FILL
XFILL_0__11995_ vdd gnd FILL
XFILL_1__13004_ vdd gnd FILL
XFILL_1__10216_ vdd gnd FILL
XFILL_0__13734_ vdd gnd FILL
XFILL_1__11196_ vdd gnd FILL
XFILL_0__8232_ vdd gnd FILL
XFILL_0__10946_ vdd gnd FILL
XFILL_2__9148_ vdd gnd FILL
X_8860_ _8860_/D _8860_/CLK _8860_/Q vdd gnd DFFPOSX1
XFILL_2__11506_ vdd gnd FILL
XFILL_1__10147_ vdd gnd FILL
XFILL_0__13665_ vdd gnd FILL
X_7811_ _7811_/A _7811_/B _7811_/Y vdd gnd OR2X2
XFILL_0__8163_ vdd gnd FILL
XFILL_0__10877_ vdd gnd FILL
XFILL_2__14225_ vdd gnd FILL
XFILL_2__9079_ vdd gnd FILL
X_8791_ _8791_/A _8791_/B _8791_/C _8791_/Y vdd gnd OAI21X1
XFILL_2__11437_ vdd gnd FILL
XFILL_1__10078_ vdd gnd FILL
XFILL_0__12616_ vdd gnd FILL
XFILL_0__7114_ vdd gnd FILL
XFILL_0__13596_ vdd gnd FILL
X_7742_ _7742_/A _7742_/B _7742_/Y vdd gnd NAND2X1
XFILL_0__8094_ vdd gnd FILL
XFILL_1__13906_ vdd gnd FILL
XFILL_2__14156_ vdd gnd FILL
XFILL_2__11368_ vdd gnd FILL
X_7673_ _7673_/A _7673_/B _7673_/Y vdd gnd NOR2X1
XFILL_2__14087_ vdd gnd FILL
XFILL_1__13837_ vdd gnd FILL
X_9412_ _9412_/A _9412_/B _9412_/C _9412_/Y vdd gnd AOI21X1
XFILL_0__12478_ vdd gnd FILL
XFILL_2__13038_ vdd gnd FILL
XFILL_0__14217_ vdd gnd FILL
XFILL_0__11429_ vdd gnd FILL
XFILL_1__13768_ vdd gnd FILL
X_9343_ _9343_/A _9343_/B _9343_/C _9343_/Y vdd gnd AOI21X1
XFILL_0__8996_ vdd gnd FILL
XFILL_1__12719_ vdd gnd FILL
XFILL_0__14148_ vdd gnd FILL
XFILL_1__13699_ vdd gnd FILL
X_9274_ _9274_/A _9274_/B _9274_/Y vdd gnd NAND2X1
XFILL_0__14079_ vdd gnd FILL
X_8225_ _8225_/A _8225_/B _8225_/C _8225_/Y vdd gnd NAND3X1
XFILL_0__7878_ vdd gnd FILL
XFILL_1__8410_ vdd gnd FILL
XFILL_0__9617_ vdd gnd FILL
XFILL_1__9390_ vdd gnd FILL
X_8156_ _8156_/A _8156_/Y vdd gnd INVX2
X_7107_ _7107_/A _7107_/B _7107_/C _7107_/Y vdd gnd AOI21X1
XFILL_0__9548_ vdd gnd FILL
XFILL_1__8341_ vdd gnd FILL
X_8087_ _8087_/A _8087_/Y vdd gnd INVX2
XFILL_0__9479_ vdd gnd FILL
XFILL_1__8272_ vdd gnd FILL
XFILL_1__7223_ vdd gnd FILL
XFILL_1__7154_ vdd gnd FILL
XFILL_1_BUFX2_insert207 vdd gnd FILL
X_8989_ _8989_/A _8989_/Y vdd gnd INVX1
XFILL_1_BUFX2_insert218 vdd gnd FILL
XFILL_1_BUFX2_insert229 vdd gnd FILL
XFILL_1__7085_ vdd gnd FILL
X_11610_ _11610_/A _11610_/B _11610_/Y vdd gnd NAND2X1
X_12590_ _12590_/D _12590_/CLK _12590_/Q vdd gnd DFFPOSX1
X_11541_ _11541_/A _11541_/B _11541_/C _11541_/Y vdd gnd OAI21X1
XFILL_0_CLKBUF1_insert388 vdd gnd FILL
X_14260_ _14260_/A _14260_/B _14260_/Y vdd gnd NAND2X1
X_11472_ _11472_/A _11472_/Y vdd gnd INVX1
X_13211_ _13211_/A _13211_/B _13211_/C _13211_/D _13211_/Y vdd gnd AOI22X1
X_10423_ _10423_/A _10423_/B _10423_/Y vdd gnd AND2X2
X_14191_ _14191_/D _14191_/CLK _14191_/Q vdd gnd DFFPOSX1
XFILL_1__9726_ vdd gnd FILL
X_13142_ _13142_/A _13142_/B _13142_/C _13142_/Y vdd gnd NAND3X1
X_10354_ _10354_/A _10354_/B _10354_/Y vdd gnd NAND2X1
XFILL_2__8450_ vdd gnd FILL
XFILL_1__9657_ vdd gnd FILL
X_13073_ _13073_/A _13073_/Y vdd gnd INVX1
XFILL_2__7401_ vdd gnd FILL
X_10285_ _10285_/A _10285_/B _10285_/Y vdd gnd NOR2X1
XFILL_1__8608_ vdd gnd FILL
XFILL_1__9588_ vdd gnd FILL
XFILL_2__8381_ vdd gnd FILL
X_12024_ _12024_/A _12024_/B _12024_/Y vdd gnd AND2X2
XFILL_1__8539_ vdd gnd FILL
XFILL_2__10670_ vdd gnd FILL
XFILL_1__11050_ vdd gnd FILL
XFILL_0__10800_ vdd gnd FILL
XFILL_2__9002_ vdd gnd FILL
XFILL_0__11780_ vdd gnd FILL
XFILL_1__10001_ vdd gnd FILL
X_13975_ _13975_/A _13975_/B _13975_/C _13975_/Y vdd gnd NAND3X1
X_12926_ _12926_/A _12926_/B _12926_/Y vdd gnd AND2X2
XFILL_0__10662_ vdd gnd FILL
XFILL_2__11222_ vdd gnd FILL
X_12857_ _12857_/A _12857_/B _12857_/C _12857_/D _12857_/Y vdd gnd AOI22X1
XFILL_1__14740_ vdd gnd FILL
XFILL_0__12401_ vdd gnd FILL
XFILL_1__11952_ vdd gnd FILL
XFILL_0__10593_ vdd gnd FILL
XFILL_0__13381_ vdd gnd FILL
X_11808_ _11808_/A _11808_/B _11808_/S _11808_/Y vdd gnd MUX2X1
X_12788_ _12788_/A _12788_/B _12788_/C _12788_/Y vdd gnd AOI21X1
XFILL_2__11153_ vdd gnd FILL
XFILL_1__10903_ vdd gnd FILL
XFILL_1__14671_ vdd gnd FILL
XFILL_0__12332_ vdd gnd FILL
XFILL_1__11883_ vdd gnd FILL
X_14527_ _14527_/D _14527_/CLK _14527_/Q vdd gnd DFFPOSX1
X_11739_ _11739_/A _11739_/B _11739_/C _11739_/Y vdd gnd OAI21X1
XFILL_1__13622_ vdd gnd FILL
XFILL_2__11084_ vdd gnd FILL
XFILL_0__12263_ vdd gnd FILL
XFILL_1__10834_ vdd gnd FILL
X_14458_ _14458_/A _14458_/B _14458_/C _14458_/Y vdd gnd NAND3X1
XFILL_0__14002_ vdd gnd FILL
XFILL_0__11214_ vdd gnd FILL
XFILL_1__13553_ vdd gnd FILL
XFILL_0__7801_ vdd gnd FILL
XFILL_0__12194_ vdd gnd FILL
X_13409_ _13409_/A _13409_/Y vdd gnd INVX1
X_14389_ _14389_/A _14389_/B _14389_/C _14389_/Y vdd gnd OAI21X1
XFILL_0__8781_ vdd gnd FILL
XFILL_2__8717_ vdd gnd FILL
XFILL_1__12504_ vdd gnd FILL
XFILL_0__11145_ vdd gnd FILL
XFILL_0__7732_ vdd gnd FILL
XFILL_2__14774_ vdd gnd FILL
XFILL_2__8648_ vdd gnd FILL
XFILL_1__12435_ vdd gnd FILL
XFILL_0__11076_ vdd gnd FILL
XFILL_2__11986_ vdd gnd FILL
X_8010_ _8010_/A _8010_/B _8010_/C _8010_/Y vdd gnd OAI21X1
XFILL_0__7663_ vdd gnd FILL
XFILL_0__10027_ vdd gnd FILL
XFILL_2__8579_ vdd gnd FILL
XFILL_2__13725_ vdd gnd FILL
XFILL_0__9402_ vdd gnd FILL
XFILL_1__12366_ vdd gnd FILL
XFILL_0__7594_ vdd gnd FILL
XFILL_1__14105_ vdd gnd FILL
XFILL_2__13656_ vdd gnd FILL
XFILL_1__11317_ vdd gnd FILL
XFILL_0__14835_ vdd gnd FILL
XFILL_0__9333_ vdd gnd FILL
XFILL_1__12297_ vdd gnd FILL
X_9961_ _9961_/A _9961_/B _9961_/S _9961_/Y vdd gnd MUX2X1
XFILL_1__14036_ vdd gnd FILL
XFILL_1__11248_ vdd gnd FILL
XFILL_2__13587_ vdd gnd FILL
XFILL_0__14766_ vdd gnd FILL
XFILL_0__9264_ vdd gnd FILL
XFILL_0__11978_ vdd gnd FILL
X_8912_ _8912_/D _8912_/CLK _8912_/Q vdd gnd DFFPOSX1
X_9892_ _9892_/A _9892_/B _9892_/C _9892_/Y vdd gnd OAI21X1
XFILL_0__13717_ vdd gnd FILL
XFILL_0__8215_ vdd gnd FILL
XFILL_1__11179_ vdd gnd FILL
XFILL_0__10929_ vdd gnd FILL
XFILL_0__14697_ vdd gnd FILL
XFILL_0__9195_ vdd gnd FILL
X_8843_ _8843_/D _8843_/CLK _8843_/Q vdd gnd DFFPOSX1
XFILL_0__13648_ vdd gnd FILL
XFILL_0__8146_ vdd gnd FILL
X_8774_ _8774_/A _8774_/B _8774_/C _8774_/Y vdd gnd OAI21X1
XFILL_0__13579_ vdd gnd FILL
X_7725_ _7725_/A _7725_/B _7725_/Y vdd gnd NOR2X1
XFILL_0__8077_ vdd gnd FILL
XFILL_1__7910_ vdd gnd FILL
X_7656_ _7656_/A _7656_/B _7656_/C _7656_/Y vdd gnd AOI21X1
XFILL_1__7841_ vdd gnd FILL
X_7587_ _7587_/A _7587_/B _7587_/C _7587_/Y vdd gnd OAI21X1
X_9326_ _9326_/A _9326_/Y vdd gnd INVX1
XFILL_1__7772_ vdd gnd FILL
XFILL_0__8979_ vdd gnd FILL
XFILL_1__9511_ vdd gnd FILL
X_9257_ _9257_/A _9257_/B _9257_/C _9257_/Y vdd gnd AOI21X1
XFILL_1__9442_ vdd gnd FILL
X_8208_ _8208_/A _8208_/B _8208_/C _8208_/Y vdd gnd AOI21X1
X_9188_ _9188_/A _9188_/B _9188_/Y vdd gnd NAND2X1
X_10070_ _10070_/A _10070_/B _10070_/C _10070_/Y vdd gnd OAI21X1
XFILL_1__9373_ vdd gnd FILL
X_8139_ _8139_/A _8139_/B _8139_/C _8139_/Y vdd gnd AOI21X1
XFILL_1__8324_ vdd gnd FILL
XFILL_1__8255_ vdd gnd FILL
XFILL_1__7206_ vdd gnd FILL
X_13760_ _13760_/A _13760_/B _13760_/C _13760_/Y vdd gnd OAI21X1
X_10972_ _10972_/A _10972_/B _10972_/C _10972_/Y vdd gnd AOI21X1
XFILL_1__8186_ vdd gnd FILL
X_12711_ _12711_/A _12711_/B _12711_/C _12711_/Y vdd gnd OAI21X1
XFILL_1__7137_ vdd gnd FILL
XFILL256650x198150 vdd gnd FILL
X_13691_ _13691_/A _13691_/B _13691_/C _13691_/Y vdd gnd OAI21X1
X_12642_ _12642_/A _12642_/Y vdd gnd INVX1
X_12573_ _12573_/D _12573_/CLK _12573_/Q vdd gnd DFFPOSX1
X_14312_ _14312_/A _14312_/B _14312_/C _14312_/Y vdd gnd OAI21X1
X_11524_ _11524_/A _11524_/B _11524_/C _11524_/Y vdd gnd OAI21X1
XFILL_2__9620_ vdd gnd FILL
X_14243_ _14243_/A _14243_/Y vdd gnd INVX1
X_11455_ _11455_/A _11455_/B _11455_/Y vdd gnd NAND2X1
XFILL_1__10550_ vdd gnd FILL
X_10406_ _10406_/A _10406_/B _10406_/C _10406_/Y vdd gnd OAI21X1
X_14174_ _14174_/D _14174_/CLK _14174_/Q vdd gnd DFFPOSX1
XFILL_1__9709_ vdd gnd FILL
X_11386_ _11386_/A _11386_/B _11386_/Y vdd gnd NAND2X1
X_13125_ _13125_/A _13125_/B _13125_/Y vdd gnd NAND2X1
XFILL_1__10481_ vdd gnd FILL
X_10337_ _10337_/A _10337_/Y vdd gnd INVX1
XFILL_1__12220_ vdd gnd FILL
XFILL_0__12950_ vdd gnd FILL
X_13056_ _13056_/A _13056_/B _13056_/Y vdd gnd OR2X2
X_10268_ _10268_/A _10268_/Y vdd gnd INVX1
XFILL_2__13510_ vdd gnd FILL
XFILL_0__11901_ vdd gnd FILL
XFILL_1__12151_ vdd gnd FILL
XFILL_2__14490_ vdd gnd FILL
X_12007_ _12007_/A _12007_/B _12007_/C _12007_/Y vdd gnd OAI21X1
XFILL_0__12881_ vdd gnd FILL
XFILL_2__7315_ vdd gnd FILL
X_10199_ _10199_/A _10199_/B _10199_/Y vdd gnd NAND2X1
XFILL_1__11102_ vdd gnd FILL
XFILL_0__14620_ vdd gnd FILL
XFILL_1__12082_ vdd gnd FILL
XFILL_0__11832_ vdd gnd FILL
XFILL_2__7246_ vdd gnd FILL
XFILL_1__11033_ vdd gnd FILL
XFILL_2__13372_ vdd gnd FILL
XFILL_0__11763_ vdd gnd FILL
X_13958_ _13958_/A _13958_/B _13958_/C _13958_/Y vdd gnd OAI21X1
XFILL_2__7177_ vdd gnd FILL
XFILL_0__13502_ vdd gnd FILL
XFILL_0__8000_ vdd gnd FILL
XFILL_0__14482_ vdd gnd FILL
XFILL_0__11694_ vdd gnd FILL
X_12909_ _12909_/A _12909_/B _12909_/Y vdd gnd AND2X2
X_13889_ _13889_/A _13889_/B _13889_/S _13889_/Y vdd gnd MUX2X1
XFILL_0__10645_ vdd gnd FILL
XFILL_1__12984_ vdd gnd FILL
XFILL_1__14723_ vdd gnd FILL
XFILL_1__11935_ vdd gnd FILL
XFILL_0__13364_ vdd gnd FILL
X_7510_ _7510_/A _7510_/B _7510_/Y vdd gnd NAND2X1
XFILL_0__10576_ vdd gnd FILL
XFILL_0__9951_ vdd gnd FILL
X_8490_ _8490_/A _8490_/B _8490_/C _8490_/Y vdd gnd NAND3X1
XFILL_2__11136_ vdd gnd FILL
XFILL_1__14654_ vdd gnd FILL
XFILL_0__12315_ vdd gnd FILL
XFILL_1__11866_ vdd gnd FILL
XFILL_0__13295_ vdd gnd FILL
X_7441_ _7441_/A _7441_/B _7441_/C _7441_/D _7441_/Y vdd gnd AOI22X1
XFILL_0__9882_ vdd gnd FILL
XFILL_1__13605_ vdd gnd FILL
XFILL_2__11067_ vdd gnd FILL
XFILL_1__10817_ vdd gnd FILL
XFILL_1__14585_ vdd gnd FILL
XFILL_0__12246_ vdd gnd FILL
XFILL_1__11797_ vdd gnd FILL
XFILL_0__8833_ vdd gnd FILL
X_7372_ _7372_/A _7372_/B _7372_/Y vdd gnd AND2X2
XFILL_1__13536_ vdd gnd FILL
X_9111_ _9111_/A _9111_/B _9111_/C _9111_/Y vdd gnd OAI21X1
XFILL_0__12177_ vdd gnd FILL
XFILL_0__8764_ vdd gnd FILL
XFILL_0__11128_ vdd gnd FILL
XFILL_2_CLKBUF1_insert72 vdd gnd FILL
XFILL_1__10679_ vdd gnd FILL
X_9042_ _9042_/A _9042_/B _9042_/S _9042_/Y vdd gnd MUX2X1
XFILL_0__7715_ vdd gnd FILL
XFILL257250x248550 vdd gnd FILL
XFILL_2_CLKBUF1_insert94 vdd gnd FILL
XFILL_0__8695_ vdd gnd FILL
XFILL_1__12418_ vdd gnd FILL
XFILL_0__11059_ vdd gnd FILL
XFILL_2__11969_ vdd gnd FILL
XFILL_1__13398_ vdd gnd FILL
XFILL_0__7646_ vdd gnd FILL
XFILL_2__13708_ vdd gnd FILL
XFILL_1__12349_ vdd gnd FILL
XFILL_0__7577_ vdd gnd FILL
XFILL_2__13639_ vdd gnd FILL
XFILL_0__14818_ vdd gnd FILL
XFILL_0_BUFX2_insert10 vdd gnd FILL
XFILL_0__9316_ vdd gnd FILL
X_9944_ _9944_/A _9944_/Y vdd gnd INVX1
XFILL_0_BUFX2_insert21 vdd gnd FILL
XFILL_1__14019_ vdd gnd FILL
XFILL_0__14749_ vdd gnd FILL
XFILL_0__9247_ vdd gnd FILL
XFILL_1__8040_ vdd gnd FILL
X_9875_ _9875_/A _9875_/B _9875_/C _9875_/D _9875_/Y vdd gnd AOI22X1
XFILL_0__9178_ vdd gnd FILL
X_8826_ _8826_/A _8826_/B _8826_/Y vdd gnd NAND2X1
XFILL_0__8129_ vdd gnd FILL
X_8757_ _8757_/A _8757_/B _8757_/Y vdd gnd NAND2X1
XFILL_1__9991_ vdd gnd FILL
X_7708_ _7708_/A _7708_/Y vdd gnd INVX1
XFILL_1__8942_ vdd gnd FILL
X_8688_ _8688_/A _8688_/B _8688_/Y vdd gnd NAND2X1
X_7639_ _7639_/A _7639_/B _7639_/Y vdd gnd NAND2X1
XFILL_1__7824_ vdd gnd FILL
X_11240_ _11240_/A _11240_/B _11240_/C _11240_/Y vdd gnd OAI21X1
X_9309_ _9309_/A _9309_/B _9309_/Y vdd gnd NAND2X1
XFILL_1__7755_ vdd gnd FILL
X_11171_ _11171_/A _11171_/B _11171_/S _11171_/Y vdd gnd MUX2X1
XFILL257250x158550 vdd gnd FILL
XFILL_1__7686_ vdd gnd FILL
X_10122_ _10122_/A _10122_/B _10122_/C _10122_/Y vdd gnd OAI21X1
XFILL_1__9425_ vdd gnd FILL
X_10053_ _10053_/A _10053_/B _10053_/C _10053_/Y vdd gnd NAND3X1
XFILL_1__9356_ vdd gnd FILL
XFILL_2__7100_ vdd gnd FILL
X_14861_ _14861_/A _14861_/B _14861_/C _14861_/Y vdd gnd AOI21X1
XFILL_1__8307_ vdd gnd FILL
XFILL_1__9287_ vdd gnd FILL
XFILL256650x7350 vdd gnd FILL
X_13812_ _13812_/A _13812_/B _13812_/C _13812_/Y vdd gnd NAND3X1
XFILL_1__8238_ vdd gnd FILL
X_14792_ _14792_/A _14792_/B _14792_/C _14792_/Y vdd gnd OAI21X1
XFILL256950x3750 vdd gnd FILL
X_10955_ _10955_/A _10955_/Y vdd gnd INVX1
X_13743_ _13743_/A _13743_/B _13743_/C _13743_/Y vdd gnd NAND3X1
XFILL_1__8169_ vdd gnd FILL
X_10886_ _10886_/A _10886_/B _10886_/S _10886_/Y vdd gnd MUX2X1
X_13674_ _13674_/A _13674_/B _13674_/Y vdd gnd NAND2X1
XFILL_0__10430_ vdd gnd FILL
X_12625_ _12625_/A _12625_/B _12625_/C _12625_/Y vdd gnd OAI21X1
XFILL_1__11720_ vdd gnd FILL
XFILL_0__10361_ vdd gnd FILL
X_12556_ _12556_/D _12556_/CLK _12556_/Q vdd gnd DFFPOSX1
XFILL_0__12100_ vdd gnd FILL
XFILL_0__13080_ vdd gnd FILL
XFILL_0__10292_ vdd gnd FILL
X_11507_ _11507_/A _11507_/B _11507_/Y vdd gnd OR2X2
XFILL_2__9603_ vdd gnd FILL
X_12487_ _12487_/A _12487_/B _12487_/C _12487_/Y vdd gnd OAI21X1
XFILL_1__10602_ vdd gnd FILL
XFILL_2__12941_ vdd gnd FILL
XFILL_0__12031_ vdd gnd FILL
XFILL_1__14370_ vdd gnd FILL
XFILL_1__11582_ vdd gnd FILL
X_14226_ _14226_/A _14226_/B _14226_/Y vdd gnd NAND2X1
X_11438_ _11438_/A _11438_/B _11438_/Y vdd gnd NAND2X1
XFILL_2__9534_ vdd gnd FILL
XFILL_1__13321_ vdd gnd FILL
XFILL_1__10533_ vdd gnd FILL
XFILL_2__12872_ vdd gnd FILL
X_14157_ _14157_/A _14157_/B _14157_/Y vdd gnd NAND2X1
X_11369_ _11369_/A _11369_/B _11369_/Y vdd gnd NOR2X1
XFILL_2__9465_ vdd gnd FILL
XFILL_1__13252_ vdd gnd FILL
XFILL_0__7500_ vdd gnd FILL
XFILL_1__10464_ vdd gnd FILL
X_13108_ _13108_/A _13108_/B _13108_/C _13108_/Y vdd gnd OAI21X1
XFILL_0__13982_ vdd gnd FILL
XFILL_0__8480_ vdd gnd FILL
X_14088_ _14088_/A _14088_/B _14088_/C _14088_/D _14088_/Y vdd gnd AOI22X1
XFILL_1__12203_ vdd gnd FILL
XFILL_1__13183_ vdd gnd FILL
XFILL_0__12933_ vdd gnd FILL
XFILL_2__9396_ vdd gnd FILL
XFILL_1__10395_ vdd gnd FILL
XFILL_0__7431_ vdd gnd FILL
X_13039_ _13039_/A _13039_/B _13039_/C _13039_/Y vdd gnd AOI21X1
XFILL_1__12134_ vdd gnd FILL
XFILL_2__14473_ vdd gnd FILL
XFILL_0__12864_ vdd gnd FILL
XFILL_0__7362_ vdd gnd FILL
XFILL_0__14603_ vdd gnd FILL
X_7990_ _7990_/D _7990_/CLK _7990_/Q vdd gnd DFFPOSX1
XFILL_0__9101_ vdd gnd FILL
XFILL_0__11815_ vdd gnd FILL
XFILL_1__12065_ vdd gnd FILL
XFILL_0__12795_ vdd gnd FILL
XFILL_2__7229_ vdd gnd FILL
XFILL_0__7293_ vdd gnd FILL
XFILL_2__13355_ vdd gnd FILL
XFILL_1__11016_ vdd gnd FILL
XFILL_0__9032_ vdd gnd FILL
XFILL_0__11746_ vdd gnd FILL
X_9660_ _9660_/A _9660_/B _9660_/Y vdd gnd NAND2X1
XFILL_2__13286_ vdd gnd FILL
XFILL_0__14465_ vdd gnd FILL
X_8611_ _8611_/A _8611_/Y vdd gnd INVX1
XFILL257250x223350 vdd gnd FILL
X_9591_ _9591_/A _9591_/B _9591_/Y vdd gnd NAND2X1
XFILL_0__13416_ vdd gnd FILL
XFILL_1__12967_ vdd gnd FILL
XFILL_0__10628_ vdd gnd FILL
XFILL_0__14396_ vdd gnd FILL
X_8542_ _8542_/A _8542_/B _8542_/C _8542_/D _8542_/Y vdd gnd AOI22X1
XFILL_1__14706_ vdd gnd FILL
XFILL_1__11918_ vdd gnd FILL
XFILL_0__13347_ vdd gnd FILL
XFILL_1__12898_ vdd gnd FILL
XFILL_0__10559_ vdd gnd FILL
XFILL_0__9934_ vdd gnd FILL
X_8473_ _8473_/A _8473_/B _8473_/Y vdd gnd NAND2X1
XFILL_1__14637_ vdd gnd FILL
XFILL_1__11849_ vdd gnd FILL
XFILL_0__13278_ vdd gnd FILL
X_7424_ _7424_/A _7424_/Y vdd gnd INVX1
XFILL_0__9865_ vdd gnd FILL
XFILL_1__14568_ vdd gnd FILL
XFILL_0__12229_ vdd gnd FILL
XFILL_0__8816_ vdd gnd FILL
X_7355_ _7355_/A _7355_/Y vdd gnd INVX1
XFILL_1__13519_ vdd gnd FILL
XFILL_1__14499_ vdd gnd FILL
XFILL_1__7540_ vdd gnd FILL
XFILL_0__8747_ vdd gnd FILL
X_7286_ _7286_/A _7286_/B _7286_/C _7286_/Y vdd gnd OAI21X1
X_9025_ _9025_/A _9025_/B _9025_/C _9025_/Y vdd gnd OAI21X1
XFILL_1__7471_ vdd gnd FILL
XFILL_0__8678_ vdd gnd FILL
XFILL_1__9210_ vdd gnd FILL
XFILL_0__7629_ vdd gnd FILL
XFILL_1__9141_ vdd gnd FILL
XFILL_1__9072_ vdd gnd FILL
X_9927_ _9927_/A _9927_/B _9927_/C _9927_/Y vdd gnd OAI21X1
XFILL_1__8023_ vdd gnd FILL
X_9858_ _9858_/A _9858_/B _9858_/C _9858_/Y vdd gnd OAI21X1
X_10740_ _10740_/D _10740_/CLK _10740_/Q vdd gnd DFFPOSX1
XFILL257250x133350 vdd gnd FILL
X_8809_ _8809_/A _8809_/B _8809_/C _8809_/Y vdd gnd OAI21X1
X_9789_ _9789_/D _9789_/CLK _9789_/Q vdd gnd DFFPOSX1
X_10671_ _10671_/A _10671_/B _10671_/C _10671_/Y vdd gnd OAI21X1
XFILL_1__9974_ vdd gnd FILL
X_12410_ _12410_/A _12410_/B _12410_/Y vdd gnd NAND2X1
X_13390_ _13390_/A _13390_/B _13390_/Y vdd gnd NAND2X1
XFILL_1__8925_ vdd gnd FILL
X_12341_ _12341_/A _12341_/B _12341_/Y vdd gnd NOR2X1
X_12272_ _12272_/A _12272_/B _12272_/C _12272_/Y vdd gnd OAI21X1
XFILL_1__7807_ vdd gnd FILL
XFILL_1__8787_ vdd gnd FILL
X_14011_ _14011_/A _14011_/B _14011_/Y vdd gnd NAND2X1
X_11223_ _11223_/A _11223_/B _11223_/Y vdd gnd NAND2X1
XFILL_1__7738_ vdd gnd FILL
X_11154_ _11154_/A _11154_/B _11154_/Y vdd gnd NOR2X1
XFILL_2__9250_ vdd gnd FILL
XFILL_1__7669_ vdd gnd FILL
X_10105_ _10105_/A _10105_/B _10105_/C _10105_/Y vdd gnd OAI21X1
X_11085_ _11085_/A _11085_/B _11085_/Y vdd gnd AND2X2
XFILL_1__9408_ vdd gnd FILL
XFILL_2__9181_ vdd gnd FILL
XFILL_1__10180_ vdd gnd FILL
X_10036_ _10036_/A _10036_/B _10036_/Y vdd gnd NAND2X1
X_14913_ _14913_/A _14913_/Y vdd gnd BUFX2
XFILL_1__9339_ vdd gnd FILL
XFILL_2__11470_ vdd gnd FILL
X_14844_ _14844_/A _14844_/B _14844_/Y vdd gnd NOR2X1
XFILL_0__11600_ vdd gnd FILL
X_14775_ _14775_/A _14775_/B _14775_/C _14775_/Y vdd gnd NAND3X1
X_11987_ _11987_/A _11987_/Y vdd gnd INVX1
XFILL_0_BUFX2_insert2 vdd gnd FILL
XFILL_0__11531_ vdd gnd FILL
XFILL_1__13870_ vdd gnd FILL
X_13726_ _13726_/A _13726_/B _13726_/C _13726_/Y vdd gnd NAND3X1
X_10938_ _10938_/A _10938_/B _10938_/Y vdd gnd NOR2X1
XFILL_1__12821_ vdd gnd FILL
XFILL_0__14250_ vdd gnd FILL
XFILL_0__11462_ vdd gnd FILL
X_13657_ _13657_/A _13657_/B _13657_/Y vdd gnd NOR2X1
XFILL_2__12022_ vdd gnd FILL
X_10869_ _10869_/A _10869_/B _10869_/Y vdd gnd NAND2X1
XFILL_0__13201_ vdd gnd FILL
XFILL_0__10413_ vdd gnd FILL
XFILL_0_BUFX2_insert320 vdd gnd FILL
XFILL_1__12752_ vdd gnd FILL
X_12608_ _12608_/D _12608_/CLK _12608_/Q vdd gnd DFFPOSX1
XFILL_0__11393_ vdd gnd FILL
XFILL_0_BUFX2_insert331 vdd gnd FILL
XFILL_0_BUFX2_insert342 vdd gnd FILL
XFILL_1__11703_ vdd gnd FILL
XFILL_0_BUFX2_insert353 vdd gnd FILL
X_13588_ _13588_/A _13588_/B _13588_/C _13588_/Y vdd gnd OAI21X1
XFILL_0__13132_ vdd gnd FILL
XFILL_0_BUFX2_insert364 vdd gnd FILL
XFILL_0__10344_ vdd gnd FILL
XFILL_0_BUFX2_insert375 vdd gnd FILL
XFILL_1__12683_ vdd gnd FILL
X_12539_ _12539_/D _12539_/CLK _12539_/Q vdd gnd DFFPOSX1
XFILL_1__14422_ vdd gnd FILL
XFILL_2__13973_ vdd gnd FILL
XFILL_0__10275_ vdd gnd FILL
XFILL_0__13063_ vdd gnd FILL
XFILL_0__9650_ vdd gnd FILL
XFILL_0__12014_ vdd gnd FILL
XFILL_1__14353_ vdd gnd FILL
XFILL_2__12924_ vdd gnd FILL
XFILL_1__11565_ vdd gnd FILL
XFILL_0__8601_ vdd gnd FILL
X_14209_ _14209_/D _14209_/CLK _14209_/Q vdd gnd DFFPOSX1
X_7140_ _7140_/A _7140_/B _7140_/S _7140_/Y vdd gnd MUX2X1
XFILL_2__9517_ vdd gnd FILL
XFILL_0__9581_ vdd gnd FILL
XFILL_1__13304_ vdd gnd FILL
XFILL_1__10516_ vdd gnd FILL
XFILL_1__14284_ vdd gnd FILL
XFILL_2__12855_ vdd gnd FILL
XFILL_1__11496_ vdd gnd FILL
XFILL_0__8532_ vdd gnd FILL
XFILL_2__9448_ vdd gnd FILL
XFILL_1__13235_ vdd gnd FILL
XFILL_1__10447_ vdd gnd FILL
XFILL_2__12786_ vdd gnd FILL
XFILL_0__13965_ vdd gnd FILL
XFILL_0__8463_ vdd gnd FILL
XFILL_1__13166_ vdd gnd FILL
XFILL_2__9379_ vdd gnd FILL
XFILL_0__12916_ vdd gnd FILL
XFILL_1__10378_ vdd gnd FILL
XFILL_0__7414_ vdd gnd FILL
XFILL_0__13896_ vdd gnd FILL
XFILL_0__8394_ vdd gnd FILL
XFILL_1__12117_ vdd gnd FILL
XFILL_2__14456_ vdd gnd FILL
XFILL_0__12847_ vdd gnd FILL
XFILL_1__13097_ vdd gnd FILL
XFILL_0__7345_ vdd gnd FILL
X_7973_ _7973_/D _7973_/CLK _7973_/Q vdd gnd DFFPOSX1
XFILL_1__12048_ vdd gnd FILL
XFILL_2__14387_ vdd gnd FILL
XFILL_2__11599_ vdd gnd FILL
X_9712_ _9712_/A _9712_/B _9712_/Y vdd gnd NAND2X1
XFILL_0__12778_ vdd gnd FILL
XFILL_0__7276_ vdd gnd FILL
XFILL_0__9015_ vdd gnd FILL
XFILL_0__11729_ vdd gnd FILL
X_9643_ _9643_/A _9643_/B _9643_/Y vdd gnd NOR2X1
XFILL_0__14448_ vdd gnd FILL
XFILL_1__13999_ vdd gnd FILL
X_9574_ _9574_/A _9574_/B _9574_/C _9574_/Y vdd gnd OAI21X1
XFILL_0__14379_ vdd gnd FILL
X_8525_ _8525_/A _8525_/B _8525_/Y vdd gnd NAND2X1
XFILL_0__9917_ vdd gnd FILL
XFILL_1__8710_ vdd gnd FILL
X_8456_ _8456_/A _8456_/B _8456_/Y vdd gnd NAND2X1
XFILL_1__9690_ vdd gnd FILL
X_7407_ _7407_/A _7407_/B _7407_/Y vdd gnd NAND2X1
XFILL_0__9848_ vdd gnd FILL
XFILL_1__8641_ vdd gnd FILL
X_8387_ _8387_/A _8387_/B _8387_/S _8387_/Y vdd gnd MUX2X1
X_7338_ _7338_/A _7338_/B _7338_/C _7338_/Y vdd gnd NAND3X1
XFILL_1__8572_ vdd gnd FILL
XFILL_2_CLKBUF1_insert106 vdd gnd FILL
XFILL_1__7523_ vdd gnd FILL
X_7269_ _7269_/A _7269_/B _7269_/Y vdd gnd NOR2X1
X_9008_ _9008_/A _9008_/B _9008_/S _9008_/Y vdd gnd MUX2X1
XFILL_1__7454_ vdd gnd FILL
XFILL_1__7385_ vdd gnd FILL
X_11910_ _11910_/A _11910_/B _11910_/C _11910_/Y vdd gnd OAI21X1
XFILL_1__9124_ vdd gnd FILL
X_12890_ _12890_/A _12890_/B _12890_/Y vdd gnd NOR2X1
XFILL_1__9055_ vdd gnd FILL
X_11841_ _11841_/A _11841_/B _11841_/C _11841_/Y vdd gnd NAND3X1
X_14560_ _14560_/A _14560_/Y vdd gnd INVX1
XFILL_1__8006_ vdd gnd FILL
X_11772_ _11772_/A _11772_/B _11772_/Y vdd gnd NAND2X1
X_10723_ _10723_/D _10723_/CLK _10723_/Q vdd gnd DFFPOSX1
X_13511_ _13511_/A _13511_/B _13511_/C _13511_/Y vdd gnd OAI21X1
X_14491_ _14491_/A _14491_/B _14491_/C _14491_/Y vdd gnd OAI21X1
X_10654_ _10654_/A _10654_/B _10654_/C _10654_/Y vdd gnd OAI21X1
X_13442_ _13442_/D _13442_/CLK _13442_/Q vdd gnd DFFPOSX1
XFILL_1__9957_ vdd gnd FILL
X_13373_ _13373_/A _13373_/B _13373_/C _13373_/Y vdd gnd OAI21X1
XFILL_2__7701_ vdd gnd FILL
X_10585_ _10585_/A _10585_/B _10585_/Y vdd gnd NAND2X1
XFILL_1__9888_ vdd gnd FILL
X_12324_ _12324_/A _12324_/B _12324_/Y vdd gnd NOR2X1
XFILL_2__7632_ vdd gnd FILL
XFILL_1__8839_ vdd gnd FILL
XFILL_2__10970_ vdd gnd FILL
XFILL_0__10060_ vdd gnd FILL
X_12255_ _12255_/A _12255_/Y vdd gnd INVX1
XFILL_2__7563_ vdd gnd FILL
XFILL_1__11350_ vdd gnd FILL
X_11206_ _11206_/A _11206_/B _11206_/Y vdd gnd NAND2X1
X_12186_ _12186_/A _12186_/B _12186_/C _12186_/Y vdd gnd NAND3X1
XFILL_1__10301_ vdd gnd FILL
XFILL_2__12640_ vdd gnd FILL
XFILL_2__7494_ vdd gnd FILL
XFILL_1__11281_ vdd gnd FILL
X_11137_ _11137_/A _11137_/B _11137_/C _11137_/D _11137_/Y vdd gnd AOI22X1
XFILL_1__13020_ vdd gnd FILL
XFILL_1__10232_ vdd gnd FILL
XFILL_0__13750_ vdd gnd FILL
XFILL_0__10962_ vdd gnd FILL
X_11068_ _11068_/A _11068_/B _11068_/Y vdd gnd AND2X2
XFILL_2__11522_ vdd gnd FILL
XFILL_2__9164_ vdd gnd FILL
XFILL_0__12701_ vdd gnd FILL
XFILL_1__10163_ vdd gnd FILL
X_10019_ _10019_/A _10019_/Y vdd gnd INVX1
XFILL_0__13681_ vdd gnd FILL
XFILL_0__10893_ vdd gnd FILL
XFILL_2__9095_ vdd gnd FILL
XFILL_2__11453_ vdd gnd FILL
XFILL_0__12632_ vdd gnd FILL
XFILL_0__7130_ vdd gnd FILL
XFILL_1__10094_ vdd gnd FILL
X_14827_ _14827_/A _14827_/B _14827_/C _14827_/Y vdd gnd AOI21X1
XFILL_1__13922_ vdd gnd FILL
XFILL_2__11384_ vdd gnd FILL
X_14758_ _14758_/A _14758_/B _14758_/Y vdd gnd NOR2X1
XFILL_0__14302_ vdd gnd FILL
XFILL_1__13853_ vdd gnd FILL
XFILL_0__11514_ vdd gnd FILL
XFILL256050x219750 vdd gnd FILL
XFILL_0__12494_ vdd gnd FILL
X_13709_ _13709_/A _13709_/B _13709_/Y vdd gnd AND2X2
XFILL256650x64950 vdd gnd FILL
X_14689_ _14689_/A _14689_/Y vdd gnd INVX1
XFILL_0__14233_ vdd gnd FILL
XFILL_1__12804_ vdd gnd FILL
XFILL_2__9997_ vdd gnd FILL
XFILL_0__11445_ vdd gnd FILL
XFILL_1__13784_ vdd gnd FILL
XFILL_1__10996_ vdd gnd FILL
XFILL_2__12005_ vdd gnd FILL
XFILL_2__8948_ vdd gnd FILL
XFILL_1__12735_ vdd gnd FILL
XFILL_0_BUFX2_insert150 vdd gnd FILL
X_8310_ _8310_/A _8310_/B _8310_/C _8310_/Y vdd gnd NAND3X1
XFILL_0_BUFX2_insert161 vdd gnd FILL
XFILL_0__11376_ vdd gnd FILL
XFILL_0_BUFX2_insert172 vdd gnd FILL
X_9290_ _9290_/A _9290_/B _9290_/C _9290_/Y vdd gnd NAND3X1
XFILL_0_BUFX2_insert183 vdd gnd FILL
XFILL_0__13115_ vdd gnd FILL
XFILL_0_BUFX2_insert194 vdd gnd FILL
XFILL_0__10327_ vdd gnd FILL
XFILL_1__12666_ vdd gnd FILL
XFILL_0__9702_ vdd gnd FILL
XFILL_0__14095_ vdd gnd FILL
X_8241_ _8241_/A _8241_/B _8241_/Y vdd gnd NAND2X1
XFILL_0__7894_ vdd gnd FILL
XFILL_1__14405_ vdd gnd FILL
XFILL_2__13956_ vdd gnd FILL
XFILL_0__13046_ vdd gnd FILL
XFILL_0__10258_ vdd gnd FILL
XFILL_0__9633_ vdd gnd FILL
X_8172_ _8172_/A _8172_/Y vdd gnd INVX1
XFILL_2__12907_ vdd gnd FILL
XFILL_1__14336_ vdd gnd FILL
XFILL_1__11548_ vdd gnd FILL
XFILL_2__13887_ vdd gnd FILL
X_7123_ _7123_/A _7123_/Y vdd gnd INVX1
XFILL_0__10189_ vdd gnd FILL
XFILL_0__9564_ vdd gnd FILL
XFILL_1__14267_ vdd gnd FILL
XFILL_2__12838_ vdd gnd FILL
XFILL_1__11479_ vdd gnd FILL
XFILL_0__8515_ vdd gnd FILL
XFILL_1__13218_ vdd gnd FILL
XFILL_0__9495_ vdd gnd FILL
XFILL_0__13948_ vdd gnd FILL
XFILL_2__12769_ vdd gnd FILL
XFILL_0__8446_ vdd gnd FILL
XFILL_1__13149_ vdd gnd FILL
XFILL_0__13879_ vdd gnd FILL
XFILL_1__7170_ vdd gnd FILL
XFILL_0__8377_ vdd gnd FILL
XFILL_0__7328_ vdd gnd FILL
X_7956_ _7956_/D _7956_/CLK _7956_/Q vdd gnd DFFPOSX1
XFILL_0__7259_ vdd gnd FILL
X_7887_ _7887_/A _7887_/B _7887_/C _7887_/Y vdd gnd OAI21X1
X_9626_ _9626_/A _9626_/B _9626_/Y vdd gnd NAND2X1
X_9557_ _9557_/A _9557_/B _9557_/C _9557_/Y vdd gnd OAI21X1
XBUFX2_insert12 BUFX2_insert12/A BUFX2_insert12/Y vdd gnd BUFX2
XBUFX2_insert23 BUFX2_insert23/A BUFX2_insert23/Y vdd gnd BUFX2
X_8508_ _8508_/A _8508_/B _8508_/Y vdd gnd NAND2X1
XFILL_1__9742_ vdd gnd FILL
X_9488_ _9488_/A _9488_/B _9488_/Y vdd gnd NOR2X1
X_10370_ _10370_/A _10370_/B _10370_/C _10370_/Y vdd gnd OAI21X1
X_8439_ _8439_/A _8439_/B _8439_/Y vdd gnd NAND2X1
XFILL_1__9673_ vdd gnd FILL
XFILL_1__8624_ vdd gnd FILL
X_12040_ _12040_/A _12040_/B _12040_/Y vdd gnd NAND2X1
XFILL_1__8555_ vdd gnd FILL
XFILL_1__7506_ vdd gnd FILL
XFILL_1__8486_ vdd gnd FILL
XFILL_1__7437_ vdd gnd FILL
XFILL_2_BUFX2_insert201 vdd gnd FILL
X_13991_ _13991_/A _13991_/B _13991_/C _13991_/Y vdd gnd NAND3X1
X_12942_ _12942_/A _12942_/B _12942_/Y vdd gnd NAND2X1
XFILL_2_BUFX2_insert234 vdd gnd FILL
XFILL_1__7368_ vdd gnd FILL
XFILL_2_BUFX2_insert256 vdd gnd FILL
XFILL_1__9107_ vdd gnd FILL
XFILL_2_BUFX2_insert289 vdd gnd FILL
X_12873_ _12873_/A _12873_/B _12873_/C _12873_/Y vdd gnd OAI21X1
XFILL_1__7299_ vdd gnd FILL
X_14612_ _14612_/A _14612_/B _14612_/Y vdd gnd NOR2X1
X_11824_ _11824_/A _11824_/Y vdd gnd INVX1
XFILL_1__9038_ vdd gnd FILL
X_14543_ _14543_/D _14543_/CLK _14543_/Q vdd gnd DFFPOSX1
XFILL_2__10120_ vdd gnd FILL
X_11755_ _11755_/A _11755_/B _11755_/Y vdd gnd NAND2X1
XBUFX2_insert200 BUFX2_insert200/A BUFX2_insert200/Y vdd gnd BUFX2
XBUFX2_insert211 BUFX2_insert211/A BUFX2_insert211/Y vdd gnd BUFX2
XFILL_1__10850_ vdd gnd FILL
XBUFX2_insert222 BUFX2_insert222/A BUFX2_insert222/Y vdd gnd BUFX2
X_10706_ _10706_/D _10706_/CLK _10706_/Q vdd gnd DFFPOSX1
XBUFX2_insert233 BUFX2_insert233/A BUFX2_insert233/Y vdd gnd BUFX2
X_14474_ _14474_/A _14474_/B _14474_/Y vdd gnd NAND2X1
XBUFX2_insert244 BUFX2_insert244/A BUFX2_insert244/Y vdd gnd BUFX2
XFILL_2__10051_ vdd gnd FILL
X_11686_ _11686_/D _11686_/CLK _11686_/Q vdd gnd DFFPOSX1
XFILL_0__11230_ vdd gnd FILL
XBUFX2_insert255 BUFX2_insert255/A BUFX2_insert255/Y vdd gnd BUFX2
XBUFX2_insert266 BUFX2_insert266/A BUFX2_insert266/Y vdd gnd BUFX2
XFILL_1__10781_ vdd gnd FILL
XBUFX2_insert277 BUFX2_insert277/A BUFX2_insert277/Y vdd gnd BUFX2
X_13425_ _13425_/A _13425_/B _13425_/C _13425_/Y vdd gnd OAI21X1
X_10637_ _10637_/A _10637_/B _10637_/C _10637_/Y vdd gnd OAI21X1
XBUFX2_insert288 BUFX2_insert288/A BUFX2_insert288/Y vdd gnd BUFX2
XFILL_1__12520_ vdd gnd FILL
XBUFX2_insert299 BUFX2_insert299/A BUFX2_insert299/Y vdd gnd BUFX2
XFILL_0__11161_ vdd gnd FILL
X_10568_ _10568_/A _10568_/Y vdd gnd INVX1
X_13356_ _13356_/A _13356_/B _13356_/C _13356_/Y vdd gnd OAI21X1
XFILL_0__10112_ vdd gnd FILL
XFILL_1__12451_ vdd gnd FILL
XFILL_0__11092_ vdd gnd FILL
X_12307_ _12307_/A _12307_/Y vdd gnd INVX1
XFILL_2__7615_ vdd gnd FILL
X_10499_ _10499_/A _10499_/B _10499_/C _10499_/Y vdd gnd OAI21X1
XFILL_1__11402_ vdd gnd FILL
X_13287_ _13287_/A _13287_/Y vdd gnd INVX1
XFILL_0__14920_ vdd gnd FILL
XFILL_0__10043_ vdd gnd FILL
XFILL_1__12382_ vdd gnd FILL
XFILL_2__10953_ vdd gnd FILL
X_12238_ _12238_/A _12238_/B _12238_/C _12238_/D _12238_/Y vdd gnd AOI22X1
XFILL_1__14121_ vdd gnd FILL
XFILL_2__7546_ vdd gnd FILL
XFILL_1__11333_ vdd gnd FILL
XFILL_2__13672_ vdd gnd FILL
XFILL_0__14851_ vdd gnd FILL
XFILL_2__10884_ vdd gnd FILL
X_12169_ _12169_/A _12169_/B _12169_/Y vdd gnd NAND2X1
XFILL_1__14052_ vdd gnd FILL
XFILL_0__13802_ vdd gnd FILL
XFILL_2__7477_ vdd gnd FILL
XFILL_1__11264_ vdd gnd FILL
XFILL_0__14782_ vdd gnd FILL
XFILL_0__8300_ vdd gnd FILL
XFILL_0__9280_ vdd gnd FILL
XFILL_0__11994_ vdd gnd FILL
XFILL_1__13003_ vdd gnd FILL
XFILL_1__10215_ vdd gnd FILL
XFILL_0__13733_ vdd gnd FILL
XFILL_0__8231_ vdd gnd FILL
XFILL_1__11195_ vdd gnd FILL
XFILL_0__10945_ vdd gnd FILL
XFILL_1__10146_ vdd gnd FILL
XFILL_0__13664_ vdd gnd FILL
X_7810_ _7810_/A _7810_/B _7810_/C _7810_/Y vdd gnd AOI21X1
XFILL_0__8162_ vdd gnd FILL
XFILL_0__10876_ vdd gnd FILL
X_8790_ _8790_/A _8790_/B _8790_/Y vdd gnd NAND2X1
XFILL_0__7113_ vdd gnd FILL
XFILL_1__10077_ vdd gnd FILL
XFILL_0__13595_ vdd gnd FILL
X_7741_ _7741_/A _7741_/B _7741_/Y vdd gnd OR2X2
XFILL_0__8093_ vdd gnd FILL
XFILL_2__8029_ vdd gnd FILL
XFILL_1__13905_ vdd gnd FILL
XFILL_2__10318_ vdd gnd FILL
X_7672_ _7672_/A _7672_/B _7672_/Y vdd gnd NOR2X1
XFILL_2__11298_ vdd gnd FILL
XFILL_1__13836_ vdd gnd FILL
X_9411_ _9411_/A _9411_/B _9411_/Y vdd gnd NAND2X1
XFILL_0__12477_ vdd gnd FILL
XFILL_2__10249_ vdd gnd FILL
XFILL_0__14216_ vdd gnd FILL
XFILL_0__11428_ vdd gnd FILL
XFILL_1__10979_ vdd gnd FILL
XFILL_1__13767_ vdd gnd FILL
X_9342_ _9342_/A _9342_/B _9342_/Y vdd gnd NAND2X1
XFILL_0__8995_ vdd gnd FILL
XFILL_1__12718_ vdd gnd FILL
XFILL_0__14147_ vdd gnd FILL
XFILL_0__11359_ vdd gnd FILL
XFILL_1__13698_ vdd gnd FILL
X_9273_ _9273_/A _9273_/B _9273_/Y vdd gnd NAND2X1
XFILL_1__12649_ vdd gnd FILL
XFILL_0__14078_ vdd gnd FILL
X_8224_ _8224_/A _8224_/Y vdd gnd INVX1
XFILL_0__7877_ vdd gnd FILL
XFILL_2__13939_ vdd gnd FILL
XFILL_0__13029_ vdd gnd FILL
XFILL_0__9616_ vdd gnd FILL
X_8155_ _8155_/A _8155_/Y vdd gnd INVX1
XFILL_1__14319_ vdd gnd FILL
X_7106_ _7106_/A _7106_/B _7106_/C _7106_/Y vdd gnd OAI21X1
XFILL_0__9547_ vdd gnd FILL
XFILL_1__8340_ vdd gnd FILL
X_8086_ _8086_/A _8086_/B _8086_/S _8086_/Y vdd gnd MUX2X1
XFILL_1__8271_ vdd gnd FILL
XFILL_0__9478_ vdd gnd FILL
XFILL_1__7222_ vdd gnd FILL
XFILL_0__8429_ vdd gnd FILL
XFILL_1__7153_ vdd gnd FILL
X_8988_ _8988_/A _8988_/B _8988_/S _8988_/Y vdd gnd MUX2X1
XFILL_1_BUFX2_insert208 vdd gnd FILL
XFILL_1_BUFX2_insert219 vdd gnd FILL
XFILL_1__7084_ vdd gnd FILL
X_7939_ _7939_/D _7939_/CLK _7939_/Q vdd gnd DFFPOSX1
X_11540_ _11540_/A _11540_/B _11540_/C _11540_/Y vdd gnd OAI21X1
X_9609_ _9609_/A _9609_/B _9609_/C _9609_/D _9609_/Y vdd gnd OAI22X1
XFILL_0_CLKBUF1_insert389 vdd gnd FILL
X_11471_ _11471_/A _11471_/B _11471_/Y vdd gnd NAND2X1
X_13210_ _13210_/A _13210_/B _13210_/Y vdd gnd NOR2X1
X_10422_ _10422_/A _10422_/B _10422_/Y vdd gnd NAND2X1
XFILL_1__9725_ vdd gnd FILL
X_14190_ _14190_/D _14190_/CLK _14190_/Q vdd gnd DFFPOSX1
X_13141_ _13141_/A _13141_/B _13141_/C _13141_/Y vdd gnd OAI21X1
X_10353_ _10353_/A _10353_/B _10353_/Y vdd gnd NAND2X1
XFILL_1__9656_ vdd gnd FILL
X_13072_ _13072_/A _13072_/B _13072_/C _13072_/Y vdd gnd OAI21X1
X_10284_ _10284_/A _10284_/B _10284_/S _10284_/Y vdd gnd MUX2X1
XFILL_1__8607_ vdd gnd FILL
XFILL_1__9587_ vdd gnd FILL
X_12023_ _12023_/A _12023_/Y vdd gnd INVX1
XFILL_2__7331_ vdd gnd FILL
XFILL_1__8538_ vdd gnd FILL
XFILL_2__7262_ vdd gnd FILL
XFILL_1__8469_ vdd gnd FILL
X_13974_ _13974_/A _13974_/B _13974_/Y vdd gnd NOR2X1
XFILL_1__10000_ vdd gnd FILL
XFILL_2__7193_ vdd gnd FILL
X_12925_ _12925_/A _12925_/B _12925_/C _12925_/Y vdd gnd NAND3X1
XFILL_2__12270_ vdd gnd FILL
XFILL_0__10661_ vdd gnd FILL
X_12856_ _12856_/A _12856_/B _12856_/C _12856_/Y vdd gnd OAI21X1
XFILL_0__12400_ vdd gnd FILL
XFILL_1__11951_ vdd gnd FILL
XFILL_0__13380_ vdd gnd FILL
XFILL_0__10592_ vdd gnd FILL
X_11807_ _11807_/A _11807_/B _11807_/C _11807_/Y vdd gnd NAND3X1
XFILL_1__10902_ vdd gnd FILL
X_12787_ _12787_/A _12787_/B _12787_/C _12787_/Y vdd gnd NAND3X1
XFILL_0__12331_ vdd gnd FILL
XFILL_1__14670_ vdd gnd FILL
XFILL_1__11882_ vdd gnd FILL
X_14526_ _14526_/D _14526_/CLK _14526_/Q vdd gnd DFFPOSX1
XFILL_2__10103_ vdd gnd FILL
X_11738_ _11738_/A _11738_/B _11738_/Y vdd gnd NAND2X1
XFILL_1__13621_ vdd gnd FILL
XFILL_1__10833_ vdd gnd FILL
XFILL_0__12262_ vdd gnd FILL
X_14457_ _14457_/A _14457_/Y vdd gnd INVX1
XFILL_0__14001_ vdd gnd FILL
XFILL_2__14911_ vdd gnd FILL
XFILL_2__10034_ vdd gnd FILL
X_11669_ _11669_/D _11669_/CLK _11669_/Q vdd gnd DFFPOSX1
XFILL_0__11213_ vdd gnd FILL
XFILL_1__13552_ vdd gnd FILL
XFILL_0__7800_ vdd gnd FILL
XFILL_0__12193_ vdd gnd FILL
X_13408_ _13408_/A _13408_/B _13408_/C _13408_/Y vdd gnd OAI21X1
X_14388_ _14388_/A _14388_/B _14388_/C _14388_/Y vdd gnd NAND3X1
XFILL_0__8780_ vdd gnd FILL
XFILL_1__12503_ vdd gnd FILL
XFILL_0__11144_ vdd gnd FILL
XFILL_2__9696_ vdd gnd FILL
XFILL_0__7731_ vdd gnd FILL
X_13339_ _13339_/A _13339_/B _13339_/Y vdd gnd NAND2X1
XFILL_1__12434_ vdd gnd FILL
XFILL_0__11075_ vdd gnd FILL
XFILL_0__7662_ vdd gnd FILL
XFILL_2__10936_ vdd gnd FILL
XFILL_0__10026_ vdd gnd FILL
XFILL_1__12365_ vdd gnd FILL
XFILL_0__9401_ vdd gnd FILL
XFILL_0__7593_ vdd gnd FILL
XFILL_1__14104_ vdd gnd FILL
XFILL_2__7529_ vdd gnd FILL
XFILL_1__11316_ vdd gnd FILL
XFILL_0__14834_ vdd gnd FILL
XFILL_1__12296_ vdd gnd FILL
XFILL_2__10867_ vdd gnd FILL
XFILL_0__9332_ vdd gnd FILL
X_9960_ _9960_/A _9960_/B _9960_/S _9960_/Y vdd gnd MUX2X1
XFILL_1__14035_ vdd gnd FILL
XFILL_1__11247_ vdd gnd FILL
XFILL_0__14765_ vdd gnd FILL
XFILL_2__10798_ vdd gnd FILL
XFILL_0__11977_ vdd gnd FILL
XFILL_0__9263_ vdd gnd FILL
X_8911_ _8911_/D _8911_/CLK _8911_/Q vdd gnd DFFPOSX1
X_9891_ _9891_/A _9891_/B _9891_/C _9891_/Y vdd gnd OAI21X1
XFILL_0__13716_ vdd gnd FILL
XFILL_0__10928_ vdd gnd FILL
XFILL_1__11178_ vdd gnd FILL
XFILL_0__14696_ vdd gnd FILL
XFILL_0__8214_ vdd gnd FILL
XFILL_0__9194_ vdd gnd FILL
X_8842_ _8842_/D _8842_/CLK _8842_/Q vdd gnd DFFPOSX1
XFILL_1__10129_ vdd gnd FILL
XFILL_0__13647_ vdd gnd FILL
XFILL_2__12468_ vdd gnd FILL
XFILL_0__10859_ vdd gnd FILL
XFILL_0__8145_ vdd gnd FILL
X_8773_ _8773_/A _8773_/B _8773_/Y vdd gnd NAND2X1
XFILL_0__13578_ vdd gnd FILL
X_7724_ _7724_/A _7724_/Y vdd gnd INVX1
XFILL_0__8076_ vdd gnd FILL
XFILL_0__12529_ vdd gnd FILL
XFILL_1__14868_ vdd gnd FILL
X_7655_ _7655_/A _7655_/Y vdd gnd INVX1
XFILL_1__13819_ vdd gnd FILL
XFILL_1__14799_ vdd gnd FILL
XFILL_1__7840_ vdd gnd FILL
X_7586_ _7586_/A _7586_/B _7586_/Y vdd gnd NOR2X1
X_9325_ _9325_/A _9325_/B _9325_/C _9325_/Y vdd gnd AOI21X1
XFILL_1__7771_ vdd gnd FILL
XFILL_0__8978_ vdd gnd FILL
XFILL_1__9510_ vdd gnd FILL
X_9256_ _9256_/A _9256_/B _9256_/C _9256_/Y vdd gnd AOI21X1
X_8207_ _8207_/A _8207_/Y vdd gnd INVX1
XFILL_1__9441_ vdd gnd FILL
X_9187_ _9187_/A _9187_/B _9187_/C _9187_/Y vdd gnd NAND3X1
X_8138_ _8138_/A _8138_/B _8138_/C _8138_/Y vdd gnd AOI21X1
XFILL_1__9372_ vdd gnd FILL
XFILL_1__8323_ vdd gnd FILL
X_8069_ _8069_/A _8069_/B _8069_/Y vdd gnd NAND2X1
XFILL_1__8254_ vdd gnd FILL
XFILL_1__7205_ vdd gnd FILL
X_10971_ _10971_/A _10971_/B _10971_/Y vdd gnd NAND2X1
XFILL_1__8185_ vdd gnd FILL
X_12710_ _12710_/A _12710_/B _12710_/Y vdd gnd NAND2X1
XFILL_1__7136_ vdd gnd FILL
X_13690_ _13690_/A _13690_/B _13690_/C _13690_/Y vdd gnd AOI21X1
X_12641_ _12641_/A _12641_/B _12641_/Y vdd gnd NAND2X1
X_12572_ _12572_/D _12572_/CLK _12572_/Q vdd gnd DFFPOSX1
XFILL_2__7880_ vdd gnd FILL
X_14311_ _14311_/A _14311_/B _14311_/Y vdd gnd NAND2X1
X_11523_ _11523_/A _11523_/B _11523_/C _11523_/Y vdd gnd OAI21X1
X_14242_ _14242_/A _14242_/B _14242_/C _14242_/Y vdd gnd OAI21X1
X_11454_ _11454_/A _11454_/B _11454_/Y vdd gnd NOR2X1
XFILL_2__9550_ vdd gnd FILL
X_10405_ _10405_/A _10405_/B _10405_/C _10405_/Y vdd gnd AOI21X1
XFILL_1__9708_ vdd gnd FILL
XFILL_2__8501_ vdd gnd FILL
X_11385_ _11385_/A _11385_/B _11385_/Y vdd gnd NAND2X1
X_14173_ _14173_/D _14173_/CLK _14173_/Q vdd gnd DFFPOSX1
XFILL_2__9481_ vdd gnd FILL
XFILL_1__10480_ vdd gnd FILL
X_13124_ _13124_/A _13124_/B _13124_/C _13124_/Y vdd gnd OAI21X1
X_10336_ _10336_/A _10336_/B _10336_/C _10336_/Y vdd gnd AOI21X1
XFILL_1__9639_ vdd gnd FILL
X_13055_ _13055_/A _13055_/B _13055_/C _13055_/Y vdd gnd OAI21X1
X_10267_ _10267_/A _10267_/B _10267_/C _10267_/Y vdd gnd AOI21X1
XFILL_1__12150_ vdd gnd FILL
XFILL_0__11900_ vdd gnd FILL
X_12006_ _12006_/A _12006_/B _12006_/C _12006_/Y vdd gnd NAND3X1
XFILL_0__12880_ vdd gnd FILL
X_10198_ _10198_/A _10198_/B _10198_/Y vdd gnd NAND2X1
XFILL_1__11101_ vdd gnd FILL
XFILL_1__12081_ vdd gnd FILL
XFILL_0__11831_ vdd gnd FILL
XFILL_1__11032_ vdd gnd FILL
XFILL_0__11762_ vdd gnd FILL
X_13957_ _13957_/A _13957_/B _13957_/Y vdd gnd OR2X2
XFILL_2__12322_ vdd gnd FILL
XFILL_0__14481_ vdd gnd FILL
XFILL_0__11693_ vdd gnd FILL
X_12908_ _12908_/A _12908_/B _12908_/Y vdd gnd NAND2X1
X_13888_ _13888_/A _13888_/B _13888_/S _13888_/Y vdd gnd MUX2X1
XFILL_2__12253_ vdd gnd FILL
XFILL_0__10644_ vdd gnd FILL
XFILL_1__12983_ vdd gnd FILL
X_12839_ _12839_/A _12839_/B _12839_/C _12839_/Y vdd gnd AOI21X1
XFILL_1__14722_ vdd gnd FILL
XFILL_2__12184_ vdd gnd FILL
XFILL_1__11934_ vdd gnd FILL
XFILL_0__13363_ vdd gnd FILL
XFILL_0__10575_ vdd gnd FILL
XFILL_0__9950_ vdd gnd FILL
XFILL_0__12314_ vdd gnd FILL
XFILL_1__14653_ vdd gnd FILL
XFILL_1__11865_ vdd gnd FILL
X_14509_ _14509_/D _14509_/CLK _14509_/Q vdd gnd DFFPOSX1
XFILL_0__13294_ vdd gnd FILL
X_7440_ _7440_/A _7440_/B _7440_/Y vdd gnd NOR2X1
XFILL_0__9881_ vdd gnd FILL
XFILL_1__13604_ vdd gnd FILL
XFILL_0__12245_ vdd gnd FILL
XFILL_1__10816_ vdd gnd FILL
XFILL_1__14584_ vdd gnd FILL
XFILL_1__11796_ vdd gnd FILL
XFILL_0__8832_ vdd gnd FILL
X_7371_ _7371_/A _7371_/B _7371_/Y vdd gnd NAND2X1
XFILL_2__10017_ vdd gnd FILL
XFILL_2__9748_ vdd gnd FILL
XFILL_1__13535_ vdd gnd FILL
X_9110_ _9110_/A _9110_/B _9110_/Y vdd gnd NAND2X1
XFILL_0__12176_ vdd gnd FILL
XFILL256950x237750 vdd gnd FILL
XFILL_0__8763_ vdd gnd FILL
XFILL_2__14825_ vdd gnd FILL
XFILL_2__9679_ vdd gnd FILL
XFILL_2_CLKBUF1_insert51 vdd gnd FILL
XFILL_0__11127_ vdd gnd FILL
XFILL_1__10678_ vdd gnd FILL
X_9041_ _9041_/A _9041_/B _9041_/S _9041_/Y vdd gnd MUX2X1
XFILL_0__7714_ vdd gnd FILL
XFILL_2_CLKBUF1_insert84 vdd gnd FILL
XFILL_0__8694_ vdd gnd FILL
XFILL_1__12417_ vdd gnd FILL
XFILL_0__11058_ vdd gnd FILL
XFILL_1__13397_ vdd gnd FILL
XFILL_0__7645_ vdd gnd FILL
XFILL_0__10009_ vdd gnd FILL
XFILL_1__12348_ vdd gnd FILL
XFILL_0__7576_ vdd gnd FILL
XFILL_0__14817_ vdd gnd FILL
XFILL_1__12279_ vdd gnd FILL
XFILL_0__9315_ vdd gnd FILL
XFILL_0_BUFX2_insert11 vdd gnd FILL
X_9943_ _9943_/A _9943_/Y vdd gnd INVX8
XFILL_0_BUFX2_insert22 vdd gnd FILL
XFILL_1__14018_ vdd gnd FILL
XFILL_0__14748_ vdd gnd FILL
XFILL_0__9246_ vdd gnd FILL
X_9874_ _9874_/A _9874_/B _9874_/C _9874_/Y vdd gnd OAI21X1
XFILL_0__14679_ vdd gnd FILL
XFILL_0__9177_ vdd gnd FILL
X_8825_ _8825_/A _8825_/B _8825_/C _8825_/Y vdd gnd OAI21X1
XFILL_0__8128_ vdd gnd FILL
XFILL_1__9990_ vdd gnd FILL
X_8756_ _8756_/A _8756_/B _8756_/Y vdd gnd NAND2X1
XFILL_1__8941_ vdd gnd FILL
X_7707_ _7707_/A _7707_/B _7707_/C _7707_/Y vdd gnd OAI21X1
XFILL_0__8059_ vdd gnd FILL
X_8687_ _8687_/A _8687_/Y vdd gnd INVX1
X_7638_ _7638_/A _7638_/B _7638_/C _7638_/D _7638_/Y vdd gnd OAI22X1
XFILL_1__7823_ vdd gnd FILL
X_7569_ _7569_/A _7569_/B _7569_/Y vdd gnd AND2X2
XFILL256950x147750 vdd gnd FILL
X_9308_ _9308_/A _9308_/B _9308_/C _9308_/Y vdd gnd OAI21X1
XFILL_1__7754_ vdd gnd FILL
X_11170_ _11170_/A _11170_/B _11170_/S _11170_/Y vdd gnd MUX2X1
X_9239_ _9239_/A _9239_/B _9239_/C _9239_/Y vdd gnd OAI21X1
XFILL_1__7685_ vdd gnd FILL
X_10121_ _10121_/A _10121_/B _10121_/C _10121_/Y vdd gnd OAI21X1
XFILL_1__9424_ vdd gnd FILL
X_10052_ _10052_/A _10052_/Y vdd gnd INVX1
XFILL_1__9355_ vdd gnd FILL
X_14860_ _14860_/A _14860_/B _14860_/C _14860_/Y vdd gnd OAI21X1
XFILL_1__8306_ vdd gnd FILL
XFILL_1__9286_ vdd gnd FILL
X_13811_ _13811_/A _13811_/B _13811_/C _13811_/Y vdd gnd AOI21X1
X_14791_ _14791_/A _14791_/B _14791_/C _14791_/Y vdd gnd AOI21X1
XFILL_1__8237_ vdd gnd FILL
XFILL257250x46950 vdd gnd FILL
X_13742_ _13742_/A _13742_/Y vdd gnd INVX1
X_10954_ _10954_/A _10954_/Y vdd gnd INVX1
XFILL_1__8168_ vdd gnd FILL
XFILL_1__7119_ vdd gnd FILL
X_13673_ _13673_/A _13673_/Y vdd gnd INVX1
X_10885_ _10885_/A _10885_/B _10885_/S _10885_/Y vdd gnd MUX2X1
XFILL_2__8981_ vdd gnd FILL
XFILL_1__8099_ vdd gnd FILL
X_12624_ _12624_/A _12624_/Y vdd gnd INVX1
XFILL_0__10360_ vdd gnd FILL
X_12555_ _12555_/D _12555_/CLK _12555_/Q vdd gnd DFFPOSX1
XFILL_2__7863_ vdd gnd FILL
XFILL_0__10291_ vdd gnd FILL
X_11506_ _11506_/A _11506_/B _11506_/C _11506_/Y vdd gnd AOI21X1
XFILL_1__10601_ vdd gnd FILL
X_12486_ _12486_/A _12486_/B _12486_/Y vdd gnd NAND2X1
XFILL_0__12030_ vdd gnd FILL
XFILL_2__7794_ vdd gnd FILL
XFILL_1__11581_ vdd gnd FILL
X_14225_ _14225_/A _14225_/Y vdd gnd INVX1
X_11437_ _11437_/A _11437_/B _11437_/Y vdd gnd OR2X2
XFILL_1__10532_ vdd gnd FILL
XFILL_1__13320_ vdd gnd FILL
X_14156_ _14156_/A _14156_/B _14156_/C _14156_/Y vdd gnd OAI21X1
XFILL_2__14610_ vdd gnd FILL
X_11368_ _11368_/A _11368_/B _11368_/Y vdd gnd NOR2X1
XFILL_2__11822_ vdd gnd FILL
XFILL_1__13251_ vdd gnd FILL
XFILL_1__10463_ vdd gnd FILL
X_13107_ _13107_/A _13107_/B _13107_/C _13107_/Y vdd gnd OAI21X1
XFILL_0__13981_ vdd gnd FILL
X_10319_ _10319_/A _10319_/B _10319_/Y vdd gnd OR2X2
XFILL_2__8415_ vdd gnd FILL
XFILL_1__12202_ vdd gnd FILL
X_14087_ _14087_/A _14087_/B _14087_/Y vdd gnd NOR2X1
X_11299_ _11299_/A _11299_/Y vdd gnd INVX1
XFILL_1__13182_ vdd gnd FILL
XFILL_2__11753_ vdd gnd FILL
XFILL_1__10394_ vdd gnd FILL
XFILL_0__12932_ vdd gnd FILL
XFILL_0__7430_ vdd gnd FILL
X_13038_ _13038_/A _13038_/Y vdd gnd INVX1
XFILL_2__8346_ vdd gnd FILL
XFILL_1__12133_ vdd gnd FILL
XFILL_0__12863_ vdd gnd FILL
XFILL_0__7361_ vdd gnd FILL
XFILL_0__14602_ vdd gnd FILL
XFILL_2__10635_ vdd gnd FILL
XFILL_1__12064_ vdd gnd FILL
XFILL_0__11814_ vdd gnd FILL
XFILL_2__8277_ vdd gnd FILL
XFILL_0__9100_ vdd gnd FILL
XFILL_0__12794_ vdd gnd FILL
XFILL_0__7292_ vdd gnd FILL
XFILL_1__11015_ vdd gnd FILL
XFILL_2__10566_ vdd gnd FILL
XFILL_0__11745_ vdd gnd FILL
XFILL_0__9031_ vdd gnd FILL
XFILL_2__12305_ vdd gnd FILL
XFILL_0__14464_ vdd gnd FILL
X_8610_ _8610_/A _8610_/B _8610_/C _8610_/Y vdd gnd OAI21X1
X_9590_ _9590_/A _9590_/B _9590_/Y vdd gnd NAND2X1
XFILL_2__12236_ vdd gnd FILL
XFILL_0__13415_ vdd gnd FILL
XFILL_0__10627_ vdd gnd FILL
XFILL_1__12966_ vdd gnd FILL
XFILL_0__14395_ vdd gnd FILL
XFILL_1_BUFX2_insert380 vdd gnd FILL
X_8541_ _8541_/A _8541_/B _8541_/C _8541_/Y vdd gnd AOI21X1
XFILL_1__14705_ vdd gnd FILL
XFILL_1__11917_ vdd gnd FILL
XFILL_2__12167_ vdd gnd FILL
XFILL_0__13346_ vdd gnd FILL
XFILL_0__10558_ vdd gnd FILL
XFILL_1__12897_ vdd gnd FILL
XFILL_0__9933_ vdd gnd FILL
X_8472_ _8472_/A _8472_/B _8472_/Y vdd gnd NAND2X1
XFILL_1__14636_ vdd gnd FILL
XFILL_2__12098_ vdd gnd FILL
XFILL_1__11848_ vdd gnd FILL
XFILL_0__13277_ vdd gnd FILL
X_7423_ _7423_/A _7423_/B _7423_/Y vdd gnd NAND2X1
XFILL_0__10489_ vdd gnd FILL
XFILL_0__9864_ vdd gnd FILL
XFILL_0__12228_ vdd gnd FILL
XFILL_1__14567_ vdd gnd FILL
XFILL_0__8815_ vdd gnd FILL
XFILL_1__11779_ vdd gnd FILL
X_7354_ _7354_/A _7354_/B _7354_/C _7354_/Y vdd gnd AOI21X1
XFILL_1__13518_ vdd gnd FILL
XFILL257250x7350 vdd gnd FILL
XFILL_0__12159_ vdd gnd FILL
XFILL_1__14498_ vdd gnd FILL
XFILL_0__8746_ vdd gnd FILL
X_7285_ _7285_/A _7285_/B _7285_/Y vdd gnd NAND2X1
XFILL_2__14808_ vdd gnd FILL
X_9024_ _9024_/A _9024_/B _9024_/Y vdd gnd NAND2X1
XFILL257550x3750 vdd gnd FILL
XFILL_1__7470_ vdd gnd FILL
XFILL_0__8677_ vdd gnd FILL
XFILL_2__14739_ vdd gnd FILL
XFILL_0__7628_ vdd gnd FILL
XFILL_1__9140_ vdd gnd FILL
XFILL_0__7559_ vdd gnd FILL
XFILL_1__9071_ vdd gnd FILL
X_9926_ _9926_/A _9926_/Y vdd gnd INVX2
XFILL256950x122550 vdd gnd FILL
XFILL_0__9229_ vdd gnd FILL
XFILL_1__8022_ vdd gnd FILL
X_9857_ _9857_/A _9857_/B _9857_/C _9857_/D _9857_/Y vdd gnd AOI22X1
X_8808_ _8808_/A _8808_/B _8808_/C _8808_/Y vdd gnd OAI21X1
X_9788_ _9788_/D _9788_/CLK _9788_/Q vdd gnd DFFPOSX1
X_10670_ _10670_/A _10670_/B _10670_/C _10670_/Y vdd gnd OAI21X1
XFILL_1__9973_ vdd gnd FILL
X_8739_ _8739_/A _8739_/B _8739_/C _8739_/Y vdd gnd OAI21X1
XFILL_1__8924_ vdd gnd FILL
X_12340_ _12340_/A _12340_/B _12340_/C _12340_/D _12340_/Y vdd gnd OAI22X1
XFILL_1__7806_ vdd gnd FILL
X_12271_ _12271_/A _12271_/B _12271_/Y vdd gnd AND2X2
XFILL257250x21750 vdd gnd FILL
XFILL_1__8786_ vdd gnd FILL
X_14010_ _14010_/A _14010_/B _14010_/C _14010_/Y vdd gnd OAI21X1
X_11222_ _11222_/A _11222_/B _11222_/Y vdd gnd NAND2X1
XFILL_1__7737_ vdd gnd FILL
X_11153_ _11153_/A _11153_/B _11153_/Y vdd gnd NAND2X1
XFILL_1__7668_ vdd gnd FILL
X_10104_ _10104_/A _10104_/Y vdd gnd INVX1
X_11084_ _11084_/A _11084_/B _11084_/C _11084_/Y vdd gnd NAND3X1
XFILL_1__9407_ vdd gnd FILL
XFILL_2__8200_ vdd gnd FILL
XFILL_1__7599_ vdd gnd FILL
X_10035_ _10035_/A _10035_/B _10035_/C _10035_/Y vdd gnd OAI21X1
X_14912_ _14912_/A _14912_/Y vdd gnd BUFX2
XFILL_1__9338_ vdd gnd FILL
XFILL_2__8131_ vdd gnd FILL
X_14843_ _14843_/A _14843_/B _14843_/C _14843_/D _14843_/Y vdd gnd AOI22X1
XFILL_1__9269_ vdd gnd FILL
XFILL_2__8062_ vdd gnd FILL
XFILL_2__10420_ vdd gnd FILL
X_14774_ _14774_/A _14774_/B _14774_/Y vdd gnd NOR2X1
XFILL_2__10351_ vdd gnd FILL
X_11986_ _11986_/A _11986_/B _11986_/Y vdd gnd AND2X2
XFILL_0_BUFX2_insert3 vdd gnd FILL
XFILL_0__11530_ vdd gnd FILL
X_13725_ _13725_/A _13725_/B _13725_/Y vdd gnd NAND2X1
X_10937_ _10937_/A _10937_/B _10937_/C _10937_/Y vdd gnd OAI21X1
XFILL_2__10282_ vdd gnd FILL
XFILL_1__12820_ vdd gnd FILL
XFILL_0__11461_ vdd gnd FILL
X_13656_ _13656_/A _13656_/B _13656_/Y vdd gnd NOR2X1
XFILL_0__13200_ vdd gnd FILL
X_10868_ _10868_/A _10868_/Y vdd gnd INVX1
XFILL_0__10412_ vdd gnd FILL
XFILL_2__8964_ vdd gnd FILL
XFILL_0_BUFX2_insert310 vdd gnd FILL
XFILL_1__12751_ vdd gnd FILL
XFILL_0_BUFX2_insert321 vdd gnd FILL
X_12607_ _12607_/D _12607_/CLK _12607_/Q vdd gnd DFFPOSX1
XFILL_0__11392_ vdd gnd FILL
XFILL_0_BUFX2_insert332 vdd gnd FILL
XFILL_0_BUFX2_insert343 vdd gnd FILL
XFILL_2__7915_ vdd gnd FILL
X_13587_ _13587_/A _13587_/B _13587_/Y vdd gnd NAND2X1
XFILL_0__13131_ vdd gnd FILL
XFILL_1__11702_ vdd gnd FILL
X_10799_ _10799_/A _10799_/B _10799_/C _10799_/D _10799_/Y vdd gnd AOI22X1
XFILL_0_BUFX2_insert354 vdd gnd FILL
XFILL_0__10343_ vdd gnd FILL
XFILL_1__12682_ vdd gnd FILL
XFILL_0_BUFX2_insert365 vdd gnd FILL
XFILL_0_BUFX2_insert376 vdd gnd FILL
X_12538_ _12538_/D _12538_/CLK _12538_/Q vdd gnd DFFPOSX1
XFILL_2__7846_ vdd gnd FILL
XFILL_1__14421_ vdd gnd FILL
XFILL_0__13062_ vdd gnd FILL
XFILL_0__10274_ vdd gnd FILL
X_12469_ _12469_/A _12469_/B _12469_/Y vdd gnd NAND2X1
XFILL_0__12013_ vdd gnd FILL
XFILL_2__7777_ vdd gnd FILL
XFILL_1__14352_ vdd gnd FILL
XFILL_1__11564_ vdd gnd FILL
XFILL_0__8600_ vdd gnd FILL
X_14208_ _14208_/D _14208_/CLK _14208_/Q vdd gnd DFFPOSX1
XFILL_0__9580_ vdd gnd FILL
XFILL_1__10515_ vdd gnd FILL
XFILL_1__13303_ vdd gnd FILL
XFILL_1__14283_ vdd gnd FILL
XFILL_1__11495_ vdd gnd FILL
XFILL_0__8531_ vdd gnd FILL
X_14139_ _14139_/A _14139_/B _14139_/C _14139_/Y vdd gnd OAI21X1
XFILL_2__11805_ vdd gnd FILL
XFILL_1__10446_ vdd gnd FILL
XFILL_1__13234_ vdd gnd FILL
XFILL_0__13964_ vdd gnd FILL
XFILL_0__8462_ vdd gnd FILL
XFILL_1__13165_ vdd gnd FILL
XFILL_2__11736_ vdd gnd FILL
XFILL_1__10377_ vdd gnd FILL
XFILL_0__12915_ vdd gnd FILL
XFILL_0__7413_ vdd gnd FILL
XFILL_0__13895_ vdd gnd FILL
XFILL_2__8329_ vdd gnd FILL
XFILL_1__12116_ vdd gnd FILL
XFILL_0__8393_ vdd gnd FILL
XFILL_1__13096_ vdd gnd FILL
XFILL_0__12846_ vdd gnd FILL
XFILL_0__7344_ vdd gnd FILL
X_7972_ _7972_/D _7972_/CLK _7972_/Q vdd gnd DFFPOSX1
XFILL_2__10618_ vdd gnd FILL
XFILL_1__12047_ vdd gnd FILL
XFILL_0__12777_ vdd gnd FILL
X_9711_ _9711_/A _9711_/B _9711_/C _9711_/Y vdd gnd OAI21X1
XFILL_0__7275_ vdd gnd FILL
XFILL_2__10549_ vdd gnd FILL
XFILL_0__11728_ vdd gnd FILL
XFILL_0__9014_ vdd gnd FILL
X_9642_ _9642_/A _9642_/B _9642_/Y vdd gnd NAND2X1
XFILL_0__14447_ vdd gnd FILL
XFILL_1__13998_ vdd gnd FILL
X_9573_ _9573_/A _9573_/B _9573_/Y vdd gnd NOR2X1
XFILL_1__12949_ vdd gnd FILL
XFILL_0__14378_ vdd gnd FILL
X_8524_ _8524_/A _8524_/Y vdd gnd INVX1
XFILL_0__13329_ vdd gnd FILL
XFILL_0__9916_ vdd gnd FILL
X_8455_ _8455_/A _8455_/B _8455_/C _8455_/Y vdd gnd OAI21X1
XFILL_1__14619_ vdd gnd FILL
X_7406_ _7406_/A _7406_/B _7406_/C _7406_/Y vdd gnd NAND3X1
XFILL_0__9847_ vdd gnd FILL
XFILL_1__8640_ vdd gnd FILL
X_8386_ _8386_/A _8386_/B _8386_/C _8386_/Y vdd gnd OAI21X1
X_7337_ _7337_/A _7337_/B _7337_/Y vdd gnd NAND2X1
XFILL_1__8571_ vdd gnd FILL
XFILL_1__7522_ vdd gnd FILL
XFILL_0__8729_ vdd gnd FILL
X_7268_ _7268_/A _7268_/B _7268_/Y vdd gnd OR2X2
X_9007_ _9007_/A _9007_/B _9007_/Y vdd gnd NOR2X1
XFILL_1__7453_ vdd gnd FILL
X_7199_ _7199_/A _7199_/B _7199_/Y vdd gnd AND2X2
XFILL_1__7384_ vdd gnd FILL
XFILL_1__9123_ vdd gnd FILL
X_11840_ _11840_/A _11840_/B _11840_/C _11840_/Y vdd gnd AOI21X1
X_9909_ _9909_/A _9909_/Y vdd gnd INVX1
XFILL_1__9054_ vdd gnd FILL
XFILL_1__8005_ vdd gnd FILL
X_11771_ _11771_/A _11771_/Y vdd gnd INVX1
X_13510_ _13510_/A _13510_/Y vdd gnd INVX1
X_10722_ _10722_/D _10722_/CLK _10722_/Q vdd gnd DFFPOSX1
X_14490_ _14490_/A _14490_/B _14490_/C _14490_/Y vdd gnd OAI21X1
X_13441_ _13441_/D _13441_/CLK _13441_/Q vdd gnd DFFPOSX1
X_10653_ _10653_/A _10653_/B _10653_/C _10653_/Y vdd gnd OAI21X1
XFILL_1__9956_ vdd gnd FILL
X_13372_ _13372_/A _13372_/B _13372_/Y vdd gnd NAND2X1
X_10584_ _10584_/A _10584_/B _10584_/Y vdd gnd NAND2X1
XFILL_1__9887_ vdd gnd FILL
X_12323_ _12323_/A _12323_/B _12323_/Y vdd gnd NAND2X1
XFILL_1__8838_ vdd gnd FILL
X_12254_ _12254_/A _12254_/B _12254_/C _12254_/Y vdd gnd OAI21X1
XFILL_1__8769_ vdd gnd FILL
X_11205_ _11205_/A _11205_/Y vdd gnd INVX1
XFILL_1__10300_ vdd gnd FILL
X_12185_ _12185_/A _12185_/Y vdd gnd INVX1
XFILL_1__11280_ vdd gnd FILL
X_11136_ _11136_/A _11136_/B _11136_/Y vdd gnd NOR2X1
XFILL_1__10231_ vdd gnd FILL
XFILL_0__10961_ vdd gnd FILL
X_11067_ _11067_/A _11067_/B _11067_/Y vdd gnd NAND2X1
XFILL_1__10162_ vdd gnd FILL
XFILL_0__12700_ vdd gnd FILL
XFILL_0__13680_ vdd gnd FILL
X_10018_ _10018_/A _10018_/B _10018_/C _10018_/Y vdd gnd NAND3X1
XFILL_0__10892_ vdd gnd FILL
XFILL_2__8114_ vdd gnd FILL
XFILL_0__12631_ vdd gnd FILL
XFILL_1__10093_ vdd gnd FILL
X_14826_ _14826_/A _14826_/Y vdd gnd INVX1
XFILL_2__10403_ vdd gnd FILL
XFILL_2__8045_ vdd gnd FILL
XFILL_1__13921_ vdd gnd FILL
X_14757_ _14757_/A _14757_/B _14757_/C _14757_/Y vdd gnd AOI21X1
XFILL_2__13122_ vdd gnd FILL
X_11969_ _11969_/A _11969_/B _11969_/C _11969_/Y vdd gnd OAI21X1
XFILL_2__10334_ vdd gnd FILL
XFILL_0__14301_ vdd gnd FILL
XFILL_0__11513_ vdd gnd FILL
XFILL_1__13852_ vdd gnd FILL
XFILL_0__12493_ vdd gnd FILL
X_13708_ _13708_/A _13708_/B _13708_/Y vdd gnd NAND2X1
X_14688_ _14688_/A _14688_/B _14688_/C _14688_/Y vdd gnd OAI21X1
XFILL_2__10265_ vdd gnd FILL
XFILL_0__14232_ vdd gnd FILL
XFILL_1__12803_ vdd gnd FILL
XFILL_2__13053_ vdd gnd FILL
XFILL_0__11444_ vdd gnd FILL
XFILL_1__13783_ vdd gnd FILL
X_13639_ _13639_/A _13639_/Y vdd gnd INVX1
XFILL_1__10995_ vdd gnd FILL
XFILL_0_BUFX2_insert140 vdd gnd FILL
XFILL_2__10196_ vdd gnd FILL
XFILL_1__12734_ vdd gnd FILL
XFILL_0_BUFX2_insert151 vdd gnd FILL
XFILL_0__11375_ vdd gnd FILL
XFILL_0_BUFX2_insert162 vdd gnd FILL
XFILL_0__13114_ vdd gnd FILL
XFILL_0_BUFX2_insert173 vdd gnd FILL
XFILL_0__10326_ vdd gnd FILL
XFILL_0_BUFX2_insert184 vdd gnd FILL
XFILL_0__9701_ vdd gnd FILL
XFILL_0__14094_ vdd gnd FILL
XFILL_0_BUFX2_insert195 vdd gnd FILL
XFILL_1__12665_ vdd gnd FILL
X_8240_ _8240_/A _8240_/B _8240_/C _8240_/Y vdd gnd OAI21X1
XFILL_0__7893_ vdd gnd FILL
XFILL_1__14404_ vdd gnd FILL
XFILL_0__13045_ vdd gnd FILL
XFILL_0__10257_ vdd gnd FILL
XFILL_0__9632_ vdd gnd FILL
X_8171_ _8171_/A _8171_/Y vdd gnd INVX1
XFILL_1__14335_ vdd gnd FILL
XFILL_1__11547_ vdd gnd FILL
X_7122_ _7122_/A _7122_/B _7122_/Y vdd gnd NAND2X1
XFILL_0__10188_ vdd gnd FILL
XFILL_0__9563_ vdd gnd FILL
XFILL_1__14266_ vdd gnd FILL
XFILL_1__11478_ vdd gnd FILL
XFILL_0__8514_ vdd gnd FILL
XFILL_0__9494_ vdd gnd FILL
XFILL_1__13217_ vdd gnd FILL
XFILL_1__10429_ vdd gnd FILL
XFILL_0__13947_ vdd gnd FILL
XFILL_0__8445_ vdd gnd FILL
XFILL_2__11719_ vdd gnd FILL
XFILL_1__13148_ vdd gnd FILL
XFILL_0__13878_ vdd gnd FILL
XFILL_0__8376_ vdd gnd FILL
XFILL_1__13079_ vdd gnd FILL
XFILL_0__12829_ vdd gnd FILL
XFILL_0__7327_ vdd gnd FILL
X_7955_ _7955_/D _7955_/CLK _7955_/Q vdd gnd DFFPOSX1
XFILL_0__7258_ vdd gnd FILL
X_7886_ _7886_/A _7886_/B _7886_/Y vdd gnd NAND2X1
X_9625_ _9625_/A _9625_/B _9625_/Y vdd gnd NOR2X1
XFILL_0__7189_ vdd gnd FILL
X_9556_ _9556_/A _9556_/Y vdd gnd INVX1
XBUFX2_insert13 BUFX2_insert13/A BUFX2_insert13/Y vdd gnd BUFX2
XFILL_1__9741_ vdd gnd FILL
XBUFX2_insert24 BUFX2_insert24/A BUFX2_insert24/Y vdd gnd BUFX2
X_8507_ _8507_/A _8507_/B _8507_/C _8507_/Y vdd gnd NAND3X1
X_9487_ _9487_/A _9487_/B _9487_/Y vdd gnd NAND2X1
XFILL_1__9672_ vdd gnd FILL
X_8438_ _8438_/A _8438_/B _8438_/Y vdd gnd NAND2X1
XFILL_1__8623_ vdd gnd FILL
X_8369_ _8369_/A _8369_/B _8369_/Y vdd gnd NAND2X1
XFILL_1__8554_ vdd gnd FILL
XFILL_1__7505_ vdd gnd FILL
XFILL_1__8485_ vdd gnd FILL
XFILL_1__7436_ vdd gnd FILL
X_13990_ _13990_/A _13990_/B _13990_/C _13990_/Y vdd gnd OAI21X1
XFILL_2_BUFX2_insert213 vdd gnd FILL
X_12941_ _12941_/A _12941_/B _12941_/Y vdd gnd AND2X2
XFILL_1__7367_ vdd gnd FILL
XFILL_2_BUFX2_insert246 vdd gnd FILL
XFILL_1__9106_ vdd gnd FILL
XFILL_2_BUFX2_insert268 vdd gnd FILL
X_12872_ _12872_/A _12872_/Y vdd gnd INVX1
XFILL_2_BUFX2_insert279 vdd gnd FILL
XFILL_1__7298_ vdd gnd FILL
X_14611_ _14611_/A _14611_/B _14611_/Y vdd gnd OR2X2
X_11823_ _11823_/A _11823_/B _11823_/C _11823_/Y vdd gnd OAI21X1
XFILL_1__9037_ vdd gnd FILL
X_14542_ _14542_/D _14542_/CLK _14542_/Q vdd gnd DFFPOSX1
X_11754_ _11754_/A _11754_/Y vdd gnd INVX1
XFILL_2__9850_ vdd gnd FILL
XBUFX2_insert201 BUFX2_insert201/A BUFX2_insert201/Y vdd gnd BUFX2
X_10705_ _10705_/D _10705_/CLK _10705_/Q vdd gnd DFFPOSX1
XBUFX2_insert212 BUFX2_insert212/A BUFX2_insert212/Y vdd gnd BUFX2
XBUFX2_insert223 BUFX2_insert223/A BUFX2_insert223/Y vdd gnd BUFX2
XFILL_2__8801_ vdd gnd FILL
X_14473_ _14473_/A _14473_/B _14473_/C _14473_/Y vdd gnd OAI21X1
XBUFX2_insert234 BUFX2_insert234/A BUFX2_insert234/Y vdd gnd BUFX2
X_11685_ _11685_/D _11685_/CLK _11685_/Q vdd gnd DFFPOSX1
XBUFX2_insert245 BUFX2_insert245/A BUFX2_insert245/Y vdd gnd BUFX2
XBUFX2_insert256 BUFX2_insert256/A BUFX2_insert256/Y vdd gnd BUFX2
XFILL_1__10780_ vdd gnd FILL
X_13424_ _13424_/A _13424_/B _13424_/Y vdd gnd NAND2X1
XBUFX2_insert267 BUFX2_insert267/A BUFX2_insert267/Y vdd gnd BUFX2
X_10636_ _10636_/A _10636_/B _10636_/Y vdd gnd NAND2X1
XBUFX2_insert278 BUFX2_insert278/A BUFX2_insert278/Y vdd gnd BUFX2
XFILL_2__8732_ vdd gnd FILL
XFILL_1__9939_ vdd gnd FILL
XFILL257550x90150 vdd gnd FILL
XBUFX2_insert289 BUFX2_insert289/A BUFX2_insert289/Y vdd gnd BUFX2
XFILL_0__11160_ vdd gnd FILL
X_13355_ _13355_/A _13355_/Y vdd gnd INVX1
X_10567_ _10567_/A _10567_/B _10567_/Y vdd gnd NOR2X1
XFILL_0__10111_ vdd gnd FILL
XFILL_2__8663_ vdd gnd FILL
XFILL_1__12450_ vdd gnd FILL
XFILL_0__11091_ vdd gnd FILL
X_12306_ _12306_/A _12306_/B _12306_/C _12306_/Y vdd gnd OAI21X1
X_13286_ _13286_/A _13286_/B _13286_/C _13286_/D _13286_/Y vdd gnd OAI22X1
X_10498_ _10498_/A _10498_/B _10498_/C _10498_/Y vdd gnd OAI21X1
XFILL_1__11401_ vdd gnd FILL
XFILL_0__10042_ vdd gnd FILL
XFILL_1__12381_ vdd gnd FILL
X_12237_ _12237_/A _12237_/B _12237_/C _12237_/Y vdd gnd AOI21X1
XFILL_1__11332_ vdd gnd FILL
XFILL_1__14120_ vdd gnd FILL
XFILL_0__14850_ vdd gnd FILL
X_12168_ _12168_/A _12168_/B _12168_/Y vdd gnd NAND2X1
XFILL_1__14051_ vdd gnd FILL
XFILL_1__11263_ vdd gnd FILL
XFILL_0__13801_ vdd gnd FILL
XFILL_0__14781_ vdd gnd FILL
XFILL_0__11993_ vdd gnd FILL
X_11119_ _11119_/A _11119_/B _11119_/Y vdd gnd NAND2X1
XFILL_1__10214_ vdd gnd FILL
X_12099_ _12099_/A _12099_/B _12099_/C _12099_/Y vdd gnd NAND3X1
XFILL_1__13002_ vdd gnd FILL
XFILL_0__10944_ vdd gnd FILL
XFILL_0__13732_ vdd gnd FILL
XFILL_1__11194_ vdd gnd FILL
XFILL_0__8230_ vdd gnd FILL
XFILL_1__10145_ vdd gnd FILL
XFILL_2__12484_ vdd gnd FILL
XFILL_0__13663_ vdd gnd FILL
XFILL_0__10875_ vdd gnd FILL
XFILL_0__8161_ vdd gnd FILL
XFILL_2__14223_ vdd gnd FILL
XFILL_1__10076_ vdd gnd FILL
XFILL_0__13594_ vdd gnd FILL
XFILL_0__7112_ vdd gnd FILL
X_14809_ _14809_/A _14809_/B _14809_/C _14809_/Y vdd gnd AOI21X1
X_7740_ _7740_/A _7740_/B _7740_/C _7740_/Y vdd gnd OAI21X1
XFILL_0__8092_ vdd gnd FILL
XFILL_1__13904_ vdd gnd FILL
XFILL_2__14154_ vdd gnd FILL
XFILL_2__13105_ vdd gnd FILL
X_7671_ _7671_/A _7671_/B _7671_/Y vdd gnd AND2X2
XFILL_2__14085_ vdd gnd FILL
XFILL_1__13835_ vdd gnd FILL
XFILL_0__12476_ vdd gnd FILL
X_9410_ _9410_/A _9410_/B _9410_/C _9410_/Y vdd gnd OAI21X1
XFILL256650x248550 vdd gnd FILL
XFILL_2__13036_ vdd gnd FILL
XFILL_0__11427_ vdd gnd FILL
XFILL_1__13766_ vdd gnd FILL
XFILL_1__10978_ vdd gnd FILL
X_9341_ _9341_/A _9341_/B _9341_/Y vdd gnd NAND2X1
XFILL_0__8994_ vdd gnd FILL
XFILL_1__12717_ vdd gnd FILL
XFILL_2__10179_ vdd gnd FILL
XFILL_0__11358_ vdd gnd FILL
XFILL_0__14146_ vdd gnd FILL
XFILL_1__13697_ vdd gnd FILL
X_9272_ _9272_/A _9272_/Y vdd gnd INVX1
XFILL_0__10309_ vdd gnd FILL
XFILL_0__14077_ vdd gnd FILL
XFILL_1__12648_ vdd gnd FILL
XFILL_0__11289_ vdd gnd FILL
X_8223_ _8223_/A _8223_/Y vdd gnd INVX1
XFILL_0__7876_ vdd gnd FILL
XFILL_0__13028_ vdd gnd FILL
XFILL_0__9615_ vdd gnd FILL
X_8154_ _8154_/A _8154_/B _8154_/C _8154_/Y vdd gnd OAI21X1
XFILL_1__14318_ vdd gnd FILL
X_7105_ _7105_/A _7105_/Y vdd gnd INVX1
XFILL_0__9546_ vdd gnd FILL
X_8085_ _8085_/A _8085_/B _8085_/S _8085_/Y vdd gnd MUX2X1
XFILL_1__14249_ vdd gnd FILL
XFILL_0__9477_ vdd gnd FILL
XFILL_1__8270_ vdd gnd FILL
XFILL_1__7221_ vdd gnd FILL
XFILL_0__8428_ vdd gnd FILL
XFILL_1__7152_ vdd gnd FILL
XFILL_0__8359_ vdd gnd FILL
X_8987_ _8987_/A _8987_/B _8987_/C _8987_/Y vdd gnd OAI21X1
XFILL_1_BUFX2_insert209 vdd gnd FILL
X_7938_ _7938_/D _7938_/CLK _7938_/Q vdd gnd DFFPOSX1
XFILL_1__7083_ vdd gnd FILL
X_7869_ _7869_/A _7869_/B _7869_/C _7869_/Y vdd gnd OAI21X1
XFILL257550x150 vdd gnd FILL
X_9608_ _9608_/A _9608_/B _9608_/Y vdd gnd NAND2X1
X_11470_ _11470_/A _11470_/B _11470_/Y vdd gnd OR2X2
X_9539_ _9539_/A _9539_/B _9539_/Y vdd gnd NAND2X1
X_10421_ _10421_/A _10421_/B _10421_/Y vdd gnd NAND2X1
XFILL_1__9724_ vdd gnd FILL
X_13140_ _13140_/A _13140_/Y vdd gnd INVX1
X_10352_ _10352_/A _10352_/B _10352_/C _10352_/Y vdd gnd OAI21X1
XFILL_1__9655_ vdd gnd FILL
XFILL_1__8606_ vdd gnd FILL
X_13071_ _13071_/A _13071_/B _13071_/Y vdd gnd NAND2X1
X_10283_ _10283_/A _10283_/B _10283_/C _10283_/Y vdd gnd OAI21X1
XFILL_1__9586_ vdd gnd FILL
X_12022_ _12022_/A _12022_/B _12022_/Y vdd gnd NAND2X1
XFILL_1__8537_ vdd gnd FILL
XFILL_1__8468_ vdd gnd FILL
XFILL_2__9000_ vdd gnd FILL
X_13973_ _13973_/A _13973_/B _13973_/C _13973_/Y vdd gnd NAND3X1
XFILL_1__7419_ vdd gnd FILL
XFILL_1__8399_ vdd gnd FILL
X_12924_ _12924_/A _12924_/B _12924_/C _12924_/Y vdd gnd OAI21X1
XFILL_0__10660_ vdd gnd FILL
X_12855_ _12855_/A _12855_/B _12855_/C _12855_/Y vdd gnd AOI21X1
XFILL_2__11220_ vdd gnd FILL
XFILL_1__11950_ vdd gnd FILL
XFILL_0__10591_ vdd gnd FILL
X_11806_ _11806_/A _11806_/B _11806_/S _11806_/Y vdd gnd MUX2X1
XFILL_2__9902_ vdd gnd FILL
X_12786_ _12786_/A _12786_/B _12786_/C _12786_/Y vdd gnd OAI21X1
XFILL_0__12330_ vdd gnd FILL
XFILL_1__10901_ vdd gnd FILL
XFILL_2__11151_ vdd gnd FILL
XFILL_1__11881_ vdd gnd FILL
X_14525_ _14525_/D _14525_/CLK _14525_/Q vdd gnd DFFPOSX1
X_11737_ _11737_/A _11737_/Y vdd gnd INVX1
XFILL_1__13620_ vdd gnd FILL
XFILL_2__11082_ vdd gnd FILL
XFILL_0__12261_ vdd gnd FILL
XFILL_1__10832_ vdd gnd FILL
X_14456_ _14456_/A _14456_/B _14456_/C _14456_/Y vdd gnd OAI21X1
X_11668_ _11668_/D _11668_/CLK _11668_/Q vdd gnd DFFPOSX1
XFILL_0__14000_ vdd gnd FILL
XFILL_0__11212_ vdd gnd FILL
XFILL_1__13551_ vdd gnd FILL
XFILL_0__12192_ vdd gnd FILL
X_13407_ _13407_/A _13407_/B _13407_/C _13407_/Y vdd gnd OAI21X1
X_10619_ _10619_/A _10619_/B _10619_/Y vdd gnd NAND2X1
X_14387_ _14387_/A _14387_/B _14387_/Y vdd gnd NAND2X1
XFILL_2__14841_ vdd gnd FILL
XFILL_2__8715_ vdd gnd FILL
XFILL_1__12502_ vdd gnd FILL
X_11599_ _11599_/A _11599_/B _11599_/C _11599_/Y vdd gnd OAI21X1
XFILL_0__11143_ vdd gnd FILL
XFILL_0__7730_ vdd gnd FILL
X_13338_ _13338_/A _13338_/B _13338_/Y vdd gnd NAND2X1
XFILL_2__8646_ vdd gnd FILL
XFILL_2__14772_ vdd gnd FILL
XFILL_1__12433_ vdd gnd FILL
XFILL_0__11074_ vdd gnd FILL
XFILL_2__11984_ vdd gnd FILL
XFILL_0__7661_ vdd gnd FILL
X_13269_ _13269_/A _13269_/B _13269_/Y vdd gnd OR2X2
XFILL_2__13723_ vdd gnd FILL
XFILL_0__10025_ vdd gnd FILL
XFILL_2__8577_ vdd gnd FILL
XFILL_0__9400_ vdd gnd FILL
XFILL_1__12364_ vdd gnd FILL
XFILL_0__7592_ vdd gnd FILL
XFILL_1__14103_ vdd gnd FILL
XFILL_1__11315_ vdd gnd FILL
XFILL_0__14833_ vdd gnd FILL
XFILL_0__9331_ vdd gnd FILL
XFILL_1__12295_ vdd gnd FILL
XFILL256650x223350 vdd gnd FILL
XFILL257250x208950 vdd gnd FILL
XFILL_1__14034_ vdd gnd FILL
XFILL_1__11246_ vdd gnd FILL
XFILL_0__14764_ vdd gnd FILL
XFILL_0__9262_ vdd gnd FILL
XFILL_0__11976_ vdd gnd FILL
X_8910_ _8910_/D _8910_/CLK _8910_/Q vdd gnd DFFPOSX1
X_9890_ _9890_/A _9890_/B _9890_/Y vdd gnd NAND2X1
XFILL_1__11177_ vdd gnd FILL
XFILL_0__13715_ vdd gnd FILL
XFILL_0__8213_ vdd gnd FILL
XFILL_0__10927_ vdd gnd FILL
XFILL_0__14695_ vdd gnd FILL
XFILL_2__9129_ vdd gnd FILL
XFILL_0__9193_ vdd gnd FILL
X_8841_ _8841_/D _8841_/CLK _8841_/Q vdd gnd DFFPOSX1
XFILL_1__10128_ vdd gnd FILL
XFILL_0__13646_ vdd gnd FILL
XFILL_0__8144_ vdd gnd FILL
XFILL_0__10858_ vdd gnd FILL
X_8772_ _8772_/A _8772_/B _8772_/C _8772_/Y vdd gnd OAI21X1
XFILL_2__11418_ vdd gnd FILL
XFILL_1__10059_ vdd gnd FILL
XFILL_2__12398_ vdd gnd FILL
XFILL_0__13577_ vdd gnd FILL
XFILL_0__10789_ vdd gnd FILL
X_7723_ _7723_/A _7723_/Y vdd gnd INVX1
XFILL_0__8075_ vdd gnd FILL
XFILL_2__14137_ vdd gnd FILL
XFILL_2__11349_ vdd gnd FILL
XFILL_1__14867_ vdd gnd FILL
XFILL_0__12528_ vdd gnd FILL
X_7654_ _7654_/A _7654_/Y vdd gnd INVX1
XFILL_2__14068_ vdd gnd FILL
XFILL_1__13818_ vdd gnd FILL
XFILL_1__14798_ vdd gnd FILL
XFILL_0__12459_ vdd gnd FILL
XFILL_2__13019_ vdd gnd FILL
X_7585_ _7585_/A _7585_/B _7585_/C _7585_/Y vdd gnd AOI21X1
XFILL_1__13749_ vdd gnd FILL
X_9324_ _9324_/A _9324_/B _9324_/C _9324_/Y vdd gnd OAI21X1
XFILL_0__8977_ vdd gnd FILL
XFILL_1__7770_ vdd gnd FILL
XFILL_0__14129_ vdd gnd FILL
X_9255_ _9255_/A _9255_/B _9255_/Y vdd gnd NAND2X1
XFILL_1__9440_ vdd gnd FILL
X_8206_ _8206_/A _8206_/B _8206_/Y vdd gnd NAND2X1
XFILL_0__7859_ vdd gnd FILL
X_9186_ _9186_/A _9186_/B _9186_/C _9186_/Y vdd gnd NAND3X1
XFILL_1__9371_ vdd gnd FILL
X_8137_ _8137_/A _8137_/B _8137_/C _8137_/D _8137_/Y vdd gnd OAI22X1
XFILL_0__9529_ vdd gnd FILL
XFILL_1__8322_ vdd gnd FILL
X_8068_ _8068_/A _8068_/Y vdd gnd INVX1
XFILL_1__8253_ vdd gnd FILL
XFILL_1__7204_ vdd gnd FILL
X_10970_ _10970_/A _10970_/B _10970_/C _10970_/Y vdd gnd OAI21X1
XFILL_1__8184_ vdd gnd FILL
XFILL_1__7135_ vdd gnd FILL
X_12640_ _12640_/A _12640_/B _12640_/C _12640_/D _12640_/Y vdd gnd AOI22X1
X_12571_ _12571_/D _12571_/CLK _12571_/Q vdd gnd DFFPOSX1
X_14310_ _14310_/A _14310_/B _14310_/Y vdd gnd NOR2X1
X_11522_ _11522_/A _11522_/B _11522_/Y vdd gnd AND2X2
X_14241_ _14241_/A _14241_/B _14241_/Y vdd gnd NAND2X1
X_11453_ _11453_/A _11453_/Y vdd gnd INVX1
X_10404_ _10404_/A _10404_/B _10404_/Y vdd gnd NAND2X1
X_14172_ _14172_/D _14172_/CLK _14172_/Q vdd gnd DFFPOSX1
XFILL_1__9707_ vdd gnd FILL
X_11384_ _11384_/A _11384_/B _11384_/Y vdd gnd NOR2X1
XFILL257550x198150 vdd gnd FILL
XFILL_1__7899_ vdd gnd FILL
X_13123_ _13123_/A _13123_/B _13123_/Y vdd gnd NOR2X1
X_10335_ _10335_/A _10335_/B _10335_/Y vdd gnd NAND2X1
XFILL_2__8431_ vdd gnd FILL
XFILL_1__9638_ vdd gnd FILL
X_13054_ _13054_/A _13054_/B _13054_/Y vdd gnd OR2X2
X_10266_ _10266_/A _10266_/B _10266_/Y vdd gnd NAND2X1
XFILL_1__9569_ vdd gnd FILL
XFILL_2__8362_ vdd gnd FILL
X_12005_ _12005_/A _12005_/B _12005_/C _12005_/Y vdd gnd NAND3X1
X_10197_ _10197_/A _10197_/B _10197_/Y vdd gnd NAND2X1
XFILL_1__11100_ vdd gnd FILL
XFILL_2__10651_ vdd gnd FILL
XFILL_2__8293_ vdd gnd FILL
XFILL_1__12080_ vdd gnd FILL
XFILL_0__11830_ vdd gnd FILL
XFILL_1__11031_ vdd gnd FILL
XFILL_2__13370_ vdd gnd FILL
XFILL_2__10582_ vdd gnd FILL
XFILL_0__11761_ vdd gnd FILL
X_13956_ _13956_/A _13956_/B _13956_/C _13956_/Y vdd gnd NAND3X1
XFILL_0__11692_ vdd gnd FILL
XFILL_0__14480_ vdd gnd FILL
X_12907_ _12907_/A _12907_/B _12907_/C _12907_/D _12907_/Y vdd gnd AOI22X1
X_13887_ _13887_/A _13887_/B _13887_/C _13887_/Y vdd gnd NAND3X1
XFILL_0__10643_ vdd gnd FILL
XFILL_1__12982_ vdd gnd FILL
X_12838_ _12838_/A _12838_/B _12838_/C _12838_/Y vdd gnd NAND3X1
XFILL_2__11203_ vdd gnd FILL
XFILL_1__14721_ vdd gnd FILL
XFILL_1__11933_ vdd gnd FILL
XFILL_0__10574_ vdd gnd FILL
XFILL_0__13362_ vdd gnd FILL
X_12769_ _12769_/A _12769_/Y vdd gnd INVX2
XFILL_2__11134_ vdd gnd FILL
XFILL_1__14652_ vdd gnd FILL
XFILL_0__12313_ vdd gnd FILL
XFILL_1__11864_ vdd gnd FILL
XFILL_0__13293_ vdd gnd FILL
X_14508_ _14508_/D _14508_/CLK _14508_/Q vdd gnd DFFPOSX1
XFILL_0__9880_ vdd gnd FILL
XFILL_1__13603_ vdd gnd FILL
XFILL_0__12244_ vdd gnd FILL
XFILL_1__10815_ vdd gnd FILL
XFILL_2__11065_ vdd gnd FILL
XFILL_1__14583_ vdd gnd FILL
XFILL_0__8831_ vdd gnd FILL
XFILL_1__11795_ vdd gnd FILL
X_14439_ _14439_/A _14439_/B _14439_/Y vdd gnd AND2X2
X_7370_ _7370_/A _7370_/B _7370_/C _7370_/D _7370_/Y vdd gnd AOI22X1
XFILL_1__13534_ vdd gnd FILL
XFILL_0__12175_ vdd gnd FILL
XFILL_0__8762_ vdd gnd FILL
XFILL_2_CLKBUF1_insert41 vdd gnd FILL
XFILL_0__11126_ vdd gnd FILL
XFILL_1__10677_ vdd gnd FILL
XFILL_0__7713_ vdd gnd FILL
X_9040_ _9040_/A _9040_/B _9040_/S _9040_/Y vdd gnd MUX2X1
XFILL_2_CLKBUF1_insert63 vdd gnd FILL
XFILL_0__8693_ vdd gnd FILL
XFILL_2__14755_ vdd gnd FILL
XFILL_2__8629_ vdd gnd FILL
XFILL_1__12416_ vdd gnd FILL
XFILL_0__11057_ vdd gnd FILL
XFILL_2_CLKBUF1_insert96 vdd gnd FILL
XFILL_2__11967_ vdd gnd FILL
XFILL_1__13396_ vdd gnd FILL
XFILL_0__7644_ vdd gnd FILL
XFILL_2__13706_ vdd gnd FILL
XFILL_0__10008_ vdd gnd FILL
XFILL_2__14686_ vdd gnd FILL
XFILL_1__12347_ vdd gnd FILL
XFILL_2__11898_ vdd gnd FILL
XFILL_0__7575_ vdd gnd FILL
XFILL_2__13637_ vdd gnd FILL
XFILL_0__14816_ vdd gnd FILL
XFILL_0__9314_ vdd gnd FILL
XFILL_1__12278_ vdd gnd FILL
X_9942_ _9942_/A _9942_/Y vdd gnd INVX1
XFILL_0_BUFX2_insert12 vdd gnd FILL
XFILL_1__14017_ vdd gnd FILL
XFILL_1__11229_ vdd gnd FILL
XFILL_0_BUFX2_insert23 vdd gnd FILL
XFILL_2__13568_ vdd gnd FILL
XFILL_0__14747_ vdd gnd FILL
XFILL_0__9245_ vdd gnd FILL
XFILL_0__11959_ vdd gnd FILL
X_9873_ _9873_/A _9873_/B _9873_/C _9873_/Y vdd gnd OAI21X1
XFILL_0__14678_ vdd gnd FILL
XFILL_0__9176_ vdd gnd FILL
X_8824_ _8824_/A _8824_/B _8824_/Y vdd gnd NAND2X1
XFILL_0__13629_ vdd gnd FILL
XFILL_0__8127_ vdd gnd FILL
X_8755_ _8755_/A _8755_/B _8755_/C _8755_/Y vdd gnd OAI21X1
XFILL_1__14919_ vdd gnd FILL
X_7706_ _7706_/A _7706_/B _7706_/Y vdd gnd NAND2X1
XFILL_0__8058_ vdd gnd FILL
XFILL_1__8940_ vdd gnd FILL
X_8686_ _8686_/A _8686_/B _8686_/Y vdd gnd NAND2X1
X_7637_ _7637_/A _7637_/B _7637_/C _7637_/Y vdd gnd OAI21X1
XFILL_1__7822_ vdd gnd FILL
X_7568_ _7568_/A _7568_/B _7568_/Y vdd gnd NOR2X1
X_9307_ _9307_/A _9307_/B _9307_/Y vdd gnd NAND2X1
XFILL_1__7753_ vdd gnd FILL
X_7499_ _7499_/A _7499_/B _7499_/C _7499_/Y vdd gnd OAI21X1
X_9238_ _9238_/A _9238_/B _9238_/Y vdd gnd AND2X2
XFILL_1__7684_ vdd gnd FILL
X_10120_ _10120_/A _10120_/Y vdd gnd INVX1
XFILL_1__9423_ vdd gnd FILL
X_9169_ _9169_/A _9169_/Y vdd gnd INVX1
X_10051_ _10051_/A _10051_/B _10051_/C _10051_/Y vdd gnd OAI21X1
XFILL_1__9354_ vdd gnd FILL
XFILL_1__8305_ vdd gnd FILL
XFILL_1__9285_ vdd gnd FILL
X_13810_ _13810_/A _13810_/Y vdd gnd INVX1
X_14790_ _14790_/A _14790_/B _14790_/Y vdd gnd NAND2X1
XFILL_1__8236_ vdd gnd FILL
X_13741_ _13741_/A _13741_/B _13741_/C _13741_/Y vdd gnd AOI21X1
X_10953_ _10953_/A _10953_/B _10953_/C _10953_/Y vdd gnd AOI21X1
XFILL_1__8167_ vdd gnd FILL
X_13672_ _13672_/A _13672_/Y vdd gnd INVX1
XFILL_1__7118_ vdd gnd FILL
X_10884_ _10884_/A _10884_/B _10884_/S _10884_/Y vdd gnd MUX2X1
XFILL_1__8098_ vdd gnd FILL
X_12623_ _12623_/A _12623_/B _12623_/Y vdd gnd NOR2X1
X_12554_ _12554_/D _12554_/CLK _12554_/Q vdd gnd DFFPOSX1
XFILL_0__10290_ vdd gnd FILL
X_11505_ _11505_/A _11505_/B _11505_/C _11505_/Y vdd gnd OAI21X1
XFILL_2__9601_ vdd gnd FILL
X_12485_ _12485_/A _12485_/B _12485_/C _12485_/Y vdd gnd OAI21X1
XFILL_1__10600_ vdd gnd FILL
X_14224_ _14224_/A _14224_/B _14224_/C _14224_/Y vdd gnd OAI21X1
XFILL_1__11580_ vdd gnd FILL
X_11436_ _11436_/A _11436_/B _11436_/C _11436_/Y vdd gnd OAI21X1
XFILL_1__10531_ vdd gnd FILL
X_14155_ _14155_/A _14155_/B _14155_/Y vdd gnd NAND2X1
X_11367_ _11367_/A _11367_/B _11367_/Y vdd gnd AND2X2
XFILL_1__13250_ vdd gnd FILL
X_13106_ _13106_/A _13106_/B _13106_/Y vdd gnd AND2X2
XFILL_1__10462_ vdd gnd FILL
XFILL_0__13980_ vdd gnd FILL
X_10318_ _10318_/A _10318_/B _10318_/Y vdd gnd NAND2X1
X_14086_ _14086_/A _14086_/B _14086_/Y vdd gnd NOR2X1
X_11298_ _11298_/A _11298_/B _11298_/Y vdd gnd NOR2X1
XFILL_1__12201_ vdd gnd FILL
XFILL_1__13181_ vdd gnd FILL
XFILL_1__10393_ vdd gnd FILL
XFILL_0__12931_ vdd gnd FILL
X_13037_ _13037_/A _13037_/B _13037_/C _13037_/Y vdd gnd NAND3X1
X_10249_ _10249_/A _10249_/B _10249_/C _10249_/Y vdd gnd AOI21X1
XFILL_2__14471_ vdd gnd FILL
XFILL_1__12132_ vdd gnd FILL
XFILL_0__12862_ vdd gnd FILL
XFILL_0__7360_ vdd gnd FILL
XFILL_2__13422_ vdd gnd FILL
XFILL_0__14601_ vdd gnd FILL
XFILL_1__12063_ vdd gnd FILL
XFILL_0__11813_ vdd gnd FILL
XFILL_0__12793_ vdd gnd FILL
XFILL_2__7227_ vdd gnd FILL
XFILL_0__7291_ vdd gnd FILL
XFILL_1__11014_ vdd gnd FILL
XFILL_2__13353_ vdd gnd FILL
XFILL_0__9030_ vdd gnd FILL
XFILL_0__11744_ vdd gnd FILL
X_13939_ _13939_/A _13939_/B _13939_/Y vdd gnd OR2X2
XFILL_2__7158_ vdd gnd FILL
XFILL_2__13284_ vdd gnd FILL
XFILL_2__10496_ vdd gnd FILL
XFILL_0__14463_ vdd gnd FILL
XFILL_0__13414_ vdd gnd FILL
XFILL_1__12965_ vdd gnd FILL
XFILL_0__10626_ vdd gnd FILL
XFILL_0__14394_ vdd gnd FILL
XFILL_1_BUFX2_insert370 vdd gnd FILL
X_8540_ _8540_/A _8540_/Y vdd gnd INVX1
XFILL_1__14704_ vdd gnd FILL
XFILL_1_BUFX2_insert381 vdd gnd FILL
XFILL_1__11916_ vdd gnd FILL
XFILL_0__13345_ vdd gnd FILL
XFILL_0__10557_ vdd gnd FILL
XFILL_1__12896_ vdd gnd FILL
XFILL_0__9932_ vdd gnd FILL
X_8471_ _8471_/A _8471_/B _8471_/Y vdd gnd OR2X2
XFILL_2__11117_ vdd gnd FILL
XFILL_1__14635_ vdd gnd FILL
XFILL_1__11847_ vdd gnd FILL
XFILL_0__10488_ vdd gnd FILL
XFILL_0__13276_ vdd gnd FILL
X_7422_ _7422_/A _7422_/B _7422_/Y vdd gnd NAND2X1
XFILL_0__9863_ vdd gnd FILL
XFILL_2__11048_ vdd gnd FILL
XFILL_1__14566_ vdd gnd FILL
XFILL_0__12227_ vdd gnd FILL
XFILL_1__11778_ vdd gnd FILL
XFILL_0__8814_ vdd gnd FILL
X_7353_ _7353_/A _7353_/B _7353_/Y vdd gnd NOR2X1
XFILL_1__13517_ vdd gnd FILL
XFILL_1__14497_ vdd gnd FILL
XFILL_0__12158_ vdd gnd FILL
XFILL_0__8745_ vdd gnd FILL
X_7284_ _7284_/A _7284_/B _7284_/C _7284_/Y vdd gnd AOI21X1
XFILL_0__11109_ vdd gnd FILL
XFILL_0__12089_ vdd gnd FILL
X_9023_ _9023_/A _9023_/Y vdd gnd INVX1
XFILL_0__8676_ vdd gnd FILL
XFILL_1__13379_ vdd gnd FILL
XFILL_0__7627_ vdd gnd FILL
XFILL_0__7558_ vdd gnd FILL
XFILL_1__9070_ vdd gnd FILL
X_9925_ _9925_/A _9925_/B _9925_/C _9925_/Y vdd gnd OAI21X1
XFILL_0__7489_ vdd gnd FILL
XFILL_0__9228_ vdd gnd FILL
XFILL_1__8021_ vdd gnd FILL
X_9856_ _9856_/A _9856_/B _9856_/Y vdd gnd NOR2X1
XFILL_0__9159_ vdd gnd FILL
X_8807_ _8807_/A _8807_/B _8807_/C _8807_/Y vdd gnd OAI21X1
X_9787_ _9787_/D _9787_/CLK _9787_/Q vdd gnd DFFPOSX1
X_8738_ _8738_/A _8738_/B _8738_/Y vdd gnd AND2X2
XFILL_1__9972_ vdd gnd FILL
XFILL_1__8923_ vdd gnd FILL
X_8669_ _8669_/A _8669_/B _8669_/Y vdd gnd AND2X2
X_12270_ _12270_/A _12270_/B _12270_/Y vdd gnd NAND2X1
XFILL_1__7805_ vdd gnd FILL
XFILL_1__8785_ vdd gnd FILL
X_11221_ _11221_/A _11221_/B _11221_/Y vdd gnd OR2X2
XFILL_1__7736_ vdd gnd FILL
X_11152_ _11152_/A _11152_/B _11152_/C _11152_/Y vdd gnd OAI21X1
XFILL_1__7667_ vdd gnd FILL
X_10103_ _10103_/A _10103_/B _10103_/Y vdd gnd NOR2X1
X_11083_ _11083_/A _11083_/B _11083_/C _11083_/Y vdd gnd OAI21X1
XFILL_1__9406_ vdd gnd FILL
XFILL_1__7598_ vdd gnd FILL
X_14911_ _14911_/A _14911_/Y vdd gnd BUFX2
X_10034_ _10034_/A _10034_/B _10034_/Y vdd gnd NAND2X1
XFILL_1__9337_ vdd gnd FILL
X_14842_ _14842_/A _14842_/B _14842_/C _14842_/Y vdd gnd AOI21X1
XFILL_1__9268_ vdd gnd FILL
XFILL_1__8219_ vdd gnd FILL
X_14773_ _14773_/A _14773_/B _14773_/Y vdd gnd NOR2X1
X_11985_ _11985_/A _11985_/B _11985_/C _11985_/Y vdd gnd NAND3X1
XFILL_1__9199_ vdd gnd FILL
XFILL_0_BUFX2_insert4 vdd gnd FILL
X_10936_ _10936_/A _10936_/B _10936_/Y vdd gnd NAND2X1
X_13724_ _13724_/A _13724_/B _13724_/C _13724_/Y vdd gnd NAND3X1
XFILL_0__11460_ vdd gnd FILL
XFILL_2__12020_ vdd gnd FILL
X_13655_ _13655_/A _13655_/B _13655_/C _13655_/Y vdd gnd OAI21X1
X_10867_ _10867_/A _10867_/Y vdd gnd INVX8
XFILL_0__10411_ vdd gnd FILL
XFILL_1__12750_ vdd gnd FILL
XFILL_0_BUFX2_insert300 vdd gnd FILL
XFILL_0_BUFX2_insert311 vdd gnd FILL
XFILL_0__11391_ vdd gnd FILL
X_12606_ _12606_/D _12606_/CLK _12606_/Q vdd gnd DFFPOSX1
XFILL_0_BUFX2_insert322 vdd gnd FILL
X_13586_ _13586_/A _13586_/Y vdd gnd INVX1
XFILL_1__11701_ vdd gnd FILL
X_10798_ _10798_/A _10798_/B _10798_/C _10798_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert333 vdd gnd FILL
XFILL_0__13130_ vdd gnd FILL
XFILL_0_BUFX2_insert344 vdd gnd FILL
XFILL_0__10342_ vdd gnd FILL
XFILL_1__12681_ vdd gnd FILL
XFILL_0_BUFX2_insert355 vdd gnd FILL
X_12537_ _12537_/D _12537_/CLK _12537_/Q vdd gnd DFFPOSX1
XFILL_0_BUFX2_insert366 vdd gnd FILL
XFILL_1__14420_ vdd gnd FILL
XFILL_0_BUFX2_insert377 vdd gnd FILL
XFILL_0__13061_ vdd gnd FILL
XFILL_0__10273_ vdd gnd FILL
X_12468_ _12468_/A _12468_/B _12468_/C _12468_/Y vdd gnd OAI21X1
XFILL_2__12922_ vdd gnd FILL
XFILL_0__12012_ vdd gnd FILL
XFILL_1__14351_ vdd gnd FILL
XFILL_1__11563_ vdd gnd FILL
X_14207_ _14207_/D _14207_/CLK _14207_/Q vdd gnd DFFPOSX1
X_11419_ _11419_/A _11419_/Y vdd gnd INVX1
XFILL_2__9515_ vdd gnd FILL
X_12399_ _12399_/A _12399_/B _12399_/Y vdd gnd NAND2X1
XFILL_1__13302_ vdd gnd FILL
XFILL_1__10514_ vdd gnd FILL
XFILL_2__12853_ vdd gnd FILL
XFILL_1__14282_ vdd gnd FILL
XFILL_0__8530_ vdd gnd FILL
XFILL_1__11494_ vdd gnd FILL
X_14138_ _14138_/A _14138_/Y vdd gnd INVX1
XFILL_2__9446_ vdd gnd FILL
XFILL_1__13233_ vdd gnd FILL
XFILL_1__10445_ vdd gnd FILL
XFILL_0__13963_ vdd gnd FILL
XFILL_0__8461_ vdd gnd FILL
X_14069_ _14069_/A _14069_/Y vdd gnd INVX1
XFILL_1__13164_ vdd gnd FILL
XFILL_0__12914_ vdd gnd FILL
XFILL_1__10376_ vdd gnd FILL
XFILL_0__7412_ vdd gnd FILL
XFILL_0__13894_ vdd gnd FILL
XFILL_0__8392_ vdd gnd FILL
XFILL_2__14454_ vdd gnd FILL
XFILL_1__12115_ vdd gnd FILL
XFILL_1__13095_ vdd gnd FILL
XFILL_0__12845_ vdd gnd FILL
XFILL_0__7343_ vdd gnd FILL
XFILL_2__13405_ vdd gnd FILL
X_7971_ _7971_/D _7971_/CLK _7971_/Q vdd gnd DFFPOSX1
XFILL_1__12046_ vdd gnd FILL
XFILL_2__14385_ vdd gnd FILL
X_9710_ _9710_/A _9710_/B _9710_/Y vdd gnd NAND2X1
XFILL_0__12776_ vdd gnd FILL
XFILL_0__7274_ vdd gnd FILL
XFILL_2__13336_ vdd gnd FILL
XFILL_0__9013_ vdd gnd FILL
XFILL_0__11727_ vdd gnd FILL
X_9641_ _9641_/A _9641_/B _9641_/C _9641_/D _9641_/Y vdd gnd AOI22X1
XFILL_2__13267_ vdd gnd FILL
XFILL_0__14446_ vdd gnd FILL
XFILL_1__13997_ vdd gnd FILL
X_9572_ _9572_/A _9572_/Y vdd gnd INVX1
XFILL_1__12948_ vdd gnd FILL
XFILL_2__13198_ vdd gnd FILL
XFILL_0__10609_ vdd gnd FILL
XFILL_0__14377_ vdd gnd FILL
X_8523_ _8523_/A _8523_/Y vdd gnd INVX1
XFILL_0__11589_ vdd gnd FILL
XFILL_0__13328_ vdd gnd FILL
XFILL_1__12879_ vdd gnd FILL
XFILL_0__9915_ vdd gnd FILL
X_8454_ _8454_/A _8454_/B _8454_/Y vdd gnd NAND2X1
XFILL_1__14618_ vdd gnd FILL
XFILL_0__13259_ vdd gnd FILL
X_7405_ _7405_/A _7405_/B _7405_/Y vdd gnd NAND2X1
XFILL_0__9846_ vdd gnd FILL
X_8385_ _8385_/A _8385_/B _8385_/Y vdd gnd NAND2X1
X_7336_ _7336_/A _7336_/B _7336_/C _7336_/Y vdd gnd OAI21X1
XFILL_1__8570_ vdd gnd FILL
XFILL_1__7521_ vdd gnd FILL
XFILL_0__8728_ vdd gnd FILL
X_7267_ _7267_/A _7267_/B _7267_/C _7267_/Y vdd gnd OAI21X1
X_9006_ _9006_/A _9006_/B _9006_/Y vdd gnd NAND2X1
XFILL_1__7452_ vdd gnd FILL
XFILL_0__8659_ vdd gnd FILL
X_7198_ _7198_/A _7198_/B _7198_/C _7198_/Y vdd gnd NAND3X1
XFILL_1__7383_ vdd gnd FILL
XFILL_1__9122_ vdd gnd FILL
XFILL_1__9053_ vdd gnd FILL
X_9908_ _9908_/A _9908_/B _9908_/C _9908_/Y vdd gnd OAI21X1
XFILL_1__8004_ vdd gnd FILL
X_11770_ _11770_/A _11770_/B _11770_/Y vdd gnd NAND2X1
X_9839_ _9839_/D _9839_/CLK _9839_/Q vdd gnd DFFPOSX1
X_10721_ _10721_/D _10721_/CLK _10721_/Q vdd gnd DFFPOSX1
X_13440_ _13440_/D _13440_/CLK _13440_/Q vdd gnd DFFPOSX1
X_10652_ _10652_/A _10652_/B _10652_/Y vdd gnd NAND2X1
XFILL_1__9955_ vdd gnd FILL
X_13371_ _13371_/A _13371_/B _13371_/C _13371_/Y vdd gnd OAI21X1
X_10583_ _10583_/A _10583_/B _10583_/Y vdd gnd OR2X2
XFILL_1__9886_ vdd gnd FILL
X_12322_ _12322_/A _12322_/B _12322_/C _12322_/Y vdd gnd OAI21X1
XFILL_1__8837_ vdd gnd FILL
X_12253_ _12253_/A _12253_/B _12253_/C _12253_/Y vdd gnd AOI21X1
XFILL_1__8768_ vdd gnd FILL
X_11204_ _11204_/A _11204_/B _11204_/C _11204_/Y vdd gnd OAI21X1
XFILL_2__9300_ vdd gnd FILL
X_12184_ _12184_/A _12184_/B _12184_/C _12184_/Y vdd gnd AOI21X1
XFILL_1__7719_ vdd gnd FILL
XFILL_1__8699_ vdd gnd FILL
X_11135_ _11135_/A _11135_/B _11135_/Y vdd gnd NOR2X1
XFILL_2__9231_ vdd gnd FILL
XFILL_1__10230_ vdd gnd FILL
XFILL_0__10960_ vdd gnd FILL
X_11066_ _11066_/A _11066_/B _11066_/C _11066_/D _11066_/Y vdd gnd AOI22X1
XFILL_2__9162_ vdd gnd FILL
XFILL_2__11520_ vdd gnd FILL
XFILL_1__10161_ vdd gnd FILL
X_10017_ _10017_/A _10017_/B _10017_/C _10017_/Y vdd gnd OAI21X1
XFILL_0__10891_ vdd gnd FILL
XFILL_2__9093_ vdd gnd FILL
XFILL_2__11451_ vdd gnd FILL
XFILL_1__10092_ vdd gnd FILL
XFILL_0__12630_ vdd gnd FILL
X_14825_ _14825_/A _14825_/Y vdd gnd INVX1
XFILL_1__13920_ vdd gnd FILL
XFILL_2__11382_ vdd gnd FILL
X_14756_ _14756_/A _14756_/B _14756_/C _14756_/Y vdd gnd OAI21X1
XFILL_0__14300_ vdd gnd FILL
X_11968_ _11968_/A _11968_/Y vdd gnd INVX1
XFILL_1__13851_ vdd gnd FILL
XFILL_0__11512_ vdd gnd FILL
XFILL_0__12492_ vdd gnd FILL
X_13707_ _13707_/A _13707_/Y vdd gnd INVX1
X_10919_ _10919_/A _10919_/B _10919_/Y vdd gnd OR2X2
X_14687_ _14687_/A _14687_/B _14687_/C _14687_/Y vdd gnd AOI21X1
X_11899_ _11899_/A _11899_/B _11899_/C _11899_/Y vdd gnd OAI21X1
XFILL_1__12802_ vdd gnd FILL
XFILL_0__14231_ vdd gnd FILL
XFILL_2__9995_ vdd gnd FILL
XFILL_0__11443_ vdd gnd FILL
XFILL_1__13782_ vdd gnd FILL
XFILL_1__10994_ vdd gnd FILL
X_13638_ _13638_/A _13638_/B _13638_/Y vdd gnd NOR2X1
XFILL_2__12003_ vdd gnd FILL
XFILL_0_BUFX2_insert130 vdd gnd FILL
XFILL_1__12733_ vdd gnd FILL
XFILL_0_BUFX2_insert141 vdd gnd FILL
XFILL_0__11374_ vdd gnd FILL
XFILL_0_BUFX2_insert152 vdd gnd FILL
XFILL_0_BUFX2_insert163 vdd gnd FILL
X_13569_ _13569_/A _13569_/B _13569_/C _13569_/Y vdd gnd OAI21X1
XFILL_0__13113_ vdd gnd FILL
XFILL_0_BUFX2_insert174 vdd gnd FILL
XFILL_1__12664_ vdd gnd FILL
XFILL_0__10325_ vdd gnd FILL
XFILL_0_BUFX2_insert185 vdd gnd FILL
XFILL_0__9700_ vdd gnd FILL
XFILL_0__14093_ vdd gnd FILL
XFILL_0_BUFX2_insert196 vdd gnd FILL
XFILL_0__7892_ vdd gnd FILL
XFILL_1__14403_ vdd gnd FILL
XFILL_2__13954_ vdd gnd FILL
XFILL_0__10256_ vdd gnd FILL
XFILL_0__13044_ vdd gnd FILL
XFILL_0__9631_ vdd gnd FILL
X_8170_ _8170_/A _8170_/B _8170_/C _8170_/Y vdd gnd NAND3X1
XFILL_2__12905_ vdd gnd FILL
XFILL_1__14334_ vdd gnd FILL
XFILL_1__11546_ vdd gnd FILL
XFILL_2__13885_ vdd gnd FILL
XFILL_0__10187_ vdd gnd FILL
X_7121_ _7121_/A _7121_/B _7121_/C _7121_/D _7121_/Y vdd gnd AOI22X1
XFILL_0__9562_ vdd gnd FILL
XFILL_1__14265_ vdd gnd FILL
XFILL_2__12836_ vdd gnd FILL
XFILL_1__11477_ vdd gnd FILL
XFILL_0__8513_ vdd gnd FILL
XFILL_0__9493_ vdd gnd FILL
XFILL_1__13216_ vdd gnd FILL
XFILL_2__9429_ vdd gnd FILL
XFILL_1__10428_ vdd gnd FILL
XFILL_2__12767_ vdd gnd FILL
XFILL_0__13946_ vdd gnd FILL
XFILL_0__8444_ vdd gnd FILL
XFILL_1__13147_ vdd gnd FILL
XFILL_1__10359_ vdd gnd FILL
XFILL_2__12698_ vdd gnd FILL
XFILL_0__13877_ vdd gnd FILL
XFILL_0__8375_ vdd gnd FILL
XFILL_2__14437_ vdd gnd FILL
XFILL_1__13078_ vdd gnd FILL
XFILL_0__12828_ vdd gnd FILL
XFILL_0__7326_ vdd gnd FILL
X_7954_ _7954_/D _7954_/CLK _7954_/Q vdd gnd DFFPOSX1
XFILL_1__12029_ vdd gnd FILL
XFILL_2__14368_ vdd gnd FILL
XFILL_0__12759_ vdd gnd FILL
XFILL_0__7257_ vdd gnd FILL
X_7885_ _7885_/A _7885_/B _7885_/C _7885_/Y vdd gnd OAI21X1
XFILL_2__14299_ vdd gnd FILL
X_9624_ _9624_/A _9624_/Y vdd gnd INVX1
XFILL_0__7188_ vdd gnd FILL
XFILL_0__14429_ vdd gnd FILL
X_9555_ _9555_/A _9555_/B _9555_/C _9555_/Y vdd gnd OAI21X1
X_8506_ _8506_/A _8506_/B _8506_/Y vdd gnd NAND2X1
XFILL_1__9740_ vdd gnd FILL
XBUFX2_insert14 BUFX2_insert14/A BUFX2_insert14/Y vdd gnd BUFX2
X_9486_ _9486_/A _9486_/B _9486_/C _9486_/D _9486_/Y vdd gnd OAI22X1
XBUFX2_insert25 BUFX2_insert25/A BUFX2_insert25/Y vdd gnd BUFX2
X_8437_ _8437_/A _8437_/B _8437_/Y vdd gnd NOR2X1
XFILL_1__9671_ vdd gnd FILL
XFILL_1__8622_ vdd gnd FILL
X_8368_ _8368_/A _8368_/B _8368_/C _8368_/Y vdd gnd OAI21X1
XFILL256350x144150 vdd gnd FILL
X_7319_ _7319_/A _7319_/B _7319_/C _7319_/Y vdd gnd OAI21X1
XFILL_1__8553_ vdd gnd FILL
X_8299_ _8299_/A _8299_/B _8299_/C _8299_/Y vdd gnd OAI21X1
XFILL_1__7504_ vdd gnd FILL
XFILL_1__8484_ vdd gnd FILL
XFILL_1__7435_ vdd gnd FILL
XFILL_2_BUFX2_insert203 vdd gnd FILL
X_12940_ _12940_/A _12940_/Y vdd gnd INVX1
XFILL_2_BUFX2_insert225 vdd gnd FILL
XFILL_1__7366_ vdd gnd FILL
XFILL_1__9105_ vdd gnd FILL
XFILL_2_BUFX2_insert258 vdd gnd FILL
X_12871_ _12871_/A _12871_/B _12871_/C _12871_/Y vdd gnd NAND3X1
XFILL_1__7297_ vdd gnd FILL
X_14610_ _14610_/A _14610_/B _14610_/C _14610_/Y vdd gnd OAI21X1
XFILL_1__9036_ vdd gnd FILL
X_11822_ _11822_/A _11822_/B _11822_/C _11822_/Y vdd gnd AOI21X1
X_11753_ _11753_/A _11753_/Y vdd gnd INVX8
X_14541_ _14541_/D _14541_/CLK _14541_/Q vdd gnd DFFPOSX1
X_10704_ _10704_/D _10704_/CLK _10704_/Q vdd gnd DFFPOSX1
XBUFX2_insert202 BUFX2_insert202/A BUFX2_insert202/Y vdd gnd BUFX2
XBUFX2_insert213 BUFX2_insert213/A BUFX2_insert213/Y vdd gnd BUFX2
X_14472_ _14472_/A _14472_/B _14472_/Y vdd gnd NAND2X1
X_11684_ _11684_/D _11684_/CLK _11684_/Q vdd gnd DFFPOSX1
XBUFX2_insert224 BUFX2_insert224/A BUFX2_insert224/Y vdd gnd BUFX2
XBUFX2_insert235 BUFX2_insert235/A BUFX2_insert235/Y vdd gnd BUFX2
XBUFX2_insert246 BUFX2_insert246/A BUFX2_insert246/Y vdd gnd BUFX2
X_10635_ _10635_/A _10635_/B _10635_/C _10635_/Y vdd gnd OAI21X1
XBUFX2_insert257 BUFX2_insert257/A BUFX2_insert257/Y vdd gnd BUFX2
X_13423_ _13423_/A _13423_/B _13423_/C _13423_/Y vdd gnd OAI21X1
XBUFX2_insert268 BUFX2_insert268/A BUFX2_insert268/Y vdd gnd BUFX2
XBUFX2_insert279 BUFX2_insert279/A BUFX2_insert279/Y vdd gnd BUFX2
XFILL_1__9938_ vdd gnd FILL
X_13354_ _13354_/A _13354_/B _13354_/C _13354_/Y vdd gnd OAI21X1
X_10566_ _10566_/A _10566_/B _10566_/Y vdd gnd NAND2X1
XFILL_0__10110_ vdd gnd FILL
XFILL_1__9869_ vdd gnd FILL
X_12305_ _12305_/A _12305_/B _12305_/C _12305_/Y vdd gnd OAI21X1
XFILL_0__11090_ vdd gnd FILL
X_13285_ _13285_/A _13285_/B _13285_/Y vdd gnd NAND2X1
XFILL_2__7613_ vdd gnd FILL
X_10497_ _10497_/A _10497_/B _10497_/Y vdd gnd NOR2X1
XFILL_1__11400_ vdd gnd FILL
XFILL_0__10041_ vdd gnd FILL
XFILL_2__10951_ vdd gnd FILL
XFILL_2__8593_ vdd gnd FILL
XFILL_1__12380_ vdd gnd FILL
X_12236_ _12236_/A _12236_/Y vdd gnd INVX1
XFILL_2__7544_ vdd gnd FILL
XFILL_1__11331_ vdd gnd FILL
XFILL_2__13670_ vdd gnd FILL
X_12167_ _12167_/A _12167_/B _12167_/Y vdd gnd OR2X2
XFILL_2__12621_ vdd gnd FILL
XFILL_1__14050_ vdd gnd FILL
XFILL_0__13800_ vdd gnd FILL
XFILL_1__11262_ vdd gnd FILL
XFILL_0__14780_ vdd gnd FILL
X_11118_ _11118_/A _11118_/B _11118_/Y vdd gnd NAND2X1
XFILL_0__11992_ vdd gnd FILL
XFILL_2__9214_ vdd gnd FILL
X_12098_ _12098_/A _12098_/Y vdd gnd INVX1
XFILL_1__13001_ vdd gnd FILL
XFILL_1__10213_ vdd gnd FILL
XFILL_0__13731_ vdd gnd FILL
XFILL_1__11193_ vdd gnd FILL
XFILL_0__10943_ vdd gnd FILL
X_11049_ _11049_/A _11049_/B _11049_/Y vdd gnd NOR2X1
XFILL_2__11503_ vdd gnd FILL
XFILL_2__9145_ vdd gnd FILL
XFILL_1__10144_ vdd gnd FILL
XFILL_0__13662_ vdd gnd FILL
XFILL_0__8160_ vdd gnd FILL
XFILL_0__10874_ vdd gnd FILL
XFILL_2__9076_ vdd gnd FILL
XFILL_2__11434_ vdd gnd FILL
XFILL_0__7111_ vdd gnd FILL
XFILL_1__10075_ vdd gnd FILL
XFILL_0__13593_ vdd gnd FILL
X_14808_ _14808_/A _14808_/B _14808_/C _14808_/Y vdd gnd AOI21X1
XFILL_0__8091_ vdd gnd FILL
XFILL_2__11365_ vdd gnd FILL
XFILL_1__13903_ vdd gnd FILL
X_14739_ _14739_/A _14739_/B _14739_/C _14739_/Y vdd gnd AOI21X1
X_7670_ _7670_/A _7670_/B _7670_/Y vdd gnd NAND2X1
XFILL_1__13834_ vdd gnd FILL
XFILL_2__11296_ vdd gnd FILL
XFILL_0__12475_ vdd gnd FILL
XFILL256950x93750 vdd gnd FILL
XFILL_2__9978_ vdd gnd FILL
XFILL_0__11426_ vdd gnd FILL
XFILL_1__13765_ vdd gnd FILL
XFILL_1__10977_ vdd gnd FILL
X_9340_ _9340_/A _9340_/B _9340_/Y vdd gnd NAND2X1
XFILL_0__8993_ vdd gnd FILL
XFILL_1__12716_ vdd gnd FILL
XFILL_0__14145_ vdd gnd FILL
XFILL_0__11357_ vdd gnd FILL
XFILL_1__13696_ vdd gnd FILL
X_9271_ _9271_/A _9271_/B _9271_/Y vdd gnd NAND2X1
XFILL_0__10308_ vdd gnd FILL
XFILL_1__12647_ vdd gnd FILL
XFILL_0__14076_ vdd gnd FILL
X_8222_ _8222_/A _8222_/B _8222_/C _8222_/Y vdd gnd OAI21X1
XFILL_0__11288_ vdd gnd FILL
XFILL_0__7875_ vdd gnd FILL
XFILL_2__13937_ vdd gnd FILL
XFILL_0__13027_ vdd gnd FILL
XFILL_0__10239_ vdd gnd FILL
XFILL_0__9614_ vdd gnd FILL
X_8153_ _8153_/A _8153_/B _8153_/C _8153_/Y vdd gnd OAI21X1
XFILL_1__14317_ vdd gnd FILL
XFILL_1__11529_ vdd gnd FILL
XFILL_2__13868_ vdd gnd FILL
X_7104_ _7104_/A _7104_/B _7104_/Y vdd gnd NAND2X1
XFILL_0__9545_ vdd gnd FILL
X_8084_ _8084_/A _8084_/B _8084_/S _8084_/Y vdd gnd MUX2X1
XFILL_1__14248_ vdd gnd FILL
XFILL_2__12819_ vdd gnd FILL
XFILL_2__13799_ vdd gnd FILL
XFILL_0__9476_ vdd gnd FILL
XFILL_0__13929_ vdd gnd FILL
XFILL_1__7220_ vdd gnd FILL
XFILL_0__8427_ vdd gnd FILL
XFILL_1__7151_ vdd gnd FILL
XFILL_0__8358_ vdd gnd FILL
X_8986_ _8986_/A _8986_/B _8986_/Y vdd gnd NAND2X1
XFILL_0__7309_ vdd gnd FILL
X_7937_ _7937_/D _7937_/CLK _7937_/Q vdd gnd DFFPOSX1
XFILL_1__7082_ vdd gnd FILL
XFILL_0__8289_ vdd gnd FILL
X_7868_ _7868_/A _7868_/Y vdd gnd INVX1
X_9607_ _9607_/A _9607_/B _9607_/Y vdd gnd NAND2X1
X_7799_ _7799_/A _7799_/B _7799_/C _7799_/Y vdd gnd AOI21X1
X_9538_ _9538_/A _9538_/B _9538_/Y vdd gnd NAND2X1
X_10420_ _10420_/A _10420_/B _10420_/Y vdd gnd NAND2X1
XFILL_1__9723_ vdd gnd FILL
X_9469_ _9469_/A _9469_/B _9469_/C _9469_/Y vdd gnd AOI21X1
X_10351_ _10351_/A _10351_/Y vdd gnd INVX1
XFILL_1__9654_ vdd gnd FILL
X_13070_ _13070_/A _13070_/B _13070_/C _13070_/Y vdd gnd OAI21X1
X_10282_ _10282_/A _10282_/B _10282_/Y vdd gnd NAND2X1
XFILL_1__8605_ vdd gnd FILL
XFILL_1__9585_ vdd gnd FILL
X_12021_ _12021_/A _12021_/B _12021_/C _12021_/Y vdd gnd OAI21X1
XFILL_1__8536_ vdd gnd FILL
XFILL_2__7260_ vdd gnd FILL
XFILL_1__8467_ vdd gnd FILL
X_13972_ _13972_/A _13972_/Y vdd gnd INVX1
XFILL_1__7418_ vdd gnd FILL
XFILL_2__7191_ vdd gnd FILL
XFILL_1__8398_ vdd gnd FILL
X_12923_ _12923_/A _12923_/B _12923_/C _12923_/Y vdd gnd NAND3X1
XFILL_1__7349_ vdd gnd FILL
X_12854_ _12854_/A _12854_/B _12854_/Y vdd gnd NAND2X1
XFILL_0__10590_ vdd gnd FILL
X_11805_ _11805_/A _11805_/B _11805_/S _11805_/Y vdd gnd MUX2X1
XFILL_1__9019_ vdd gnd FILL
XFILL_1__10900_ vdd gnd FILL
X_12785_ _12785_/A _12785_/Y vdd gnd INVX1
XFILL_1__11880_ vdd gnd FILL
X_14524_ _14524_/D _14524_/CLK _14524_/Q vdd gnd DFFPOSX1
XFILL_2__10101_ vdd gnd FILL
X_11736_ _11736_/A _11736_/B _11736_/C _11736_/Y vdd gnd AOI21X1
XFILL_1__10831_ vdd gnd FILL
XFILL_0__12260_ vdd gnd FILL
X_14455_ _14455_/A _14455_/B _14455_/Y vdd gnd NAND2X1
XFILL_2__10032_ vdd gnd FILL
X_11667_ _11667_/D _11667_/CLK _11667_/Q vdd gnd DFFPOSX1
XFILL_0__11211_ vdd gnd FILL
XFILL_2__9763_ vdd gnd FILL
XFILL_1__13550_ vdd gnd FILL
XFILL_0__12191_ vdd gnd FILL
X_13406_ _13406_/A _13406_/Y vdd gnd INVX1
X_10618_ _10618_/A _10618_/B _10618_/Y vdd gnd NAND2X1
X_14386_ _14386_/A _14386_/B _14386_/Y vdd gnd NAND2X1
XFILL_1__12501_ vdd gnd FILL
X_11598_ _11598_/A _11598_/B _11598_/Y vdd gnd NAND2X1
XFILL_0__11142_ vdd gnd FILL
X_10549_ _10549_/A _10549_/B _10549_/Y vdd gnd NOR2X1
X_13337_ _13337_/A _13337_/Y vdd gnd INVX1
XFILL256350x21750 vdd gnd FILL
XFILL_1__12432_ vdd gnd FILL
XFILL_0__11073_ vdd gnd FILL
XFILL_0__7660_ vdd gnd FILL
X_13268_ _13268_/A _13268_/B _13268_/C _13268_/Y vdd gnd OAI21X1
XFILL_0__10024_ vdd gnd FILL
XFILL_1__12363_ vdd gnd FILL
XFILL_2__10934_ vdd gnd FILL
X_12219_ _12219_/A _12219_/Y vdd gnd INVX1
X_13199_ _13199_/A _13199_/B _13199_/Y vdd gnd OR2X2
XFILL_0__7591_ vdd gnd FILL
XFILL_1__14102_ vdd gnd FILL
XFILL_2__7527_ vdd gnd FILL
XFILL_1__11314_ vdd gnd FILL
XFILL_0__14832_ vdd gnd FILL
XFILL_2__13653_ vdd gnd FILL
XFILL_2__10865_ vdd gnd FILL
XFILL_1__12294_ vdd gnd FILL
XFILL_0__9330_ vdd gnd FILL
XFILL_1__14033_ vdd gnd FILL
XFILL_2__13584_ vdd gnd FILL
XFILL_2__7458_ vdd gnd FILL
XFILL_1__11245_ vdd gnd FILL
XFILL_0__14763_ vdd gnd FILL
XFILL_2__10796_ vdd gnd FILL
XFILL_0__9261_ vdd gnd FILL
XFILL_0__11975_ vdd gnd FILL
XFILL_2__7389_ vdd gnd FILL
XFILL_0__13714_ vdd gnd FILL
XFILL_0__8212_ vdd gnd FILL
XFILL_0__10926_ vdd gnd FILL
XFILL_1__11176_ vdd gnd FILL
XFILL_0__14694_ vdd gnd FILL
XFILL_0__9192_ vdd gnd FILL
X_8840_ _8840_/D _8840_/CLK _8840_/Q vdd gnd DFFPOSX1
XFILL_1__10127_ vdd gnd FILL
XFILL_0__13645_ vdd gnd FILL
XFILL_0__8143_ vdd gnd FILL
XFILL_0__10857_ vdd gnd FILL
X_8771_ _8771_/A _8771_/B _8771_/Y vdd gnd NAND2X1
XFILL_1__10058_ vdd gnd FILL
XFILL_0__13576_ vdd gnd FILL
X_7722_ _7722_/A _7722_/B _7722_/Y vdd gnd NAND2X1
XFILL_0__8074_ vdd gnd FILL
XFILL_0__10788_ vdd gnd FILL
XFILL_0__12527_ vdd gnd FILL
XFILL_1__14866_ vdd gnd FILL
X_7653_ _7653_/A _7653_/B _7653_/C _7653_/Y vdd gnd OAI21X1
XFILL_1__13817_ vdd gnd FILL
XFILL_2__11279_ vdd gnd FILL
XFILL_0__12458_ vdd gnd FILL
XFILL_1__14797_ vdd gnd FILL
X_7584_ _7584_/A _7584_/B _7584_/Y vdd gnd NAND2X1
XFILL_0__11409_ vdd gnd FILL
XFILL_1__13748_ vdd gnd FILL
X_9323_ _9323_/A _9323_/B _9323_/S _9323_/Y vdd gnd MUX2X1
XFILL_0__12389_ vdd gnd FILL
XFILL_0__8976_ vdd gnd FILL
XFILL_0__14128_ vdd gnd FILL
XFILL_1__13679_ vdd gnd FILL
X_9254_ _9254_/A _9254_/B _9254_/C _9254_/Y vdd gnd NAND3X1
XFILL_0__14059_ vdd gnd FILL
X_8205_ _8205_/A _8205_/B _8205_/C _8205_/Y vdd gnd NAND3X1
XFILL_0__7858_ vdd gnd FILL
X_9185_ _9185_/A _9185_/B _9185_/Y vdd gnd NAND2X1
X_8136_ _8136_/A _8136_/B _8136_/Y vdd gnd NAND2X1
XFILL_1__9370_ vdd gnd FILL
XFILL_0__7789_ vdd gnd FILL
XFILL_0__9528_ vdd gnd FILL
XFILL_1__8321_ vdd gnd FILL
X_8067_ _8067_/A _8067_/B _8067_/C _8067_/Y vdd gnd OAI21X1
XFILL_1__8252_ vdd gnd FILL
XFILL_0__9459_ vdd gnd FILL
XFILL_1__7203_ vdd gnd FILL
XFILL_1__8183_ vdd gnd FILL
XFILL_1__7134_ vdd gnd FILL
X_8969_ _8969_/A _8969_/B _8969_/C _8969_/D _8969_/Y vdd gnd AOI22X1
XFILL_0_CLKBUF1_insert100 vdd gnd FILL
X_12570_ _12570_/D _12570_/CLK _12570_/Q vdd gnd DFFPOSX1
X_11521_ _11521_/A _11521_/B _11521_/Y vdd gnd NAND2X1
X_14240_ _14240_/A _14240_/Y vdd gnd INVX1
X_11452_ _11452_/A _11452_/B _11452_/Y vdd gnd NAND2X1
X_10403_ _10403_/A _10403_/B _10403_/C _10403_/Y vdd gnd NAND3X1
X_14171_ _14171_/D _14171_/CLK _14171_/Q vdd gnd DFFPOSX1
XFILL_1__9706_ vdd gnd FILL
X_11383_ _11383_/A _11383_/Y vdd gnd INVX1
XFILL_1__7898_ vdd gnd FILL
X_13122_ _13122_/A _13122_/B _13122_/C _13122_/Y vdd gnd AOI21X1
X_10334_ _10334_/A _10334_/B _10334_/C _10334_/Y vdd gnd OAI21X1
XFILL_1__9637_ vdd gnd FILL
X_13053_ _13053_/A _13053_/B _13053_/Y vdd gnd NAND2X1
X_10265_ _10265_/A _10265_/B _10265_/Y vdd gnd NAND2X1
XFILL_1__9568_ vdd gnd FILL
X_12004_ _12004_/A _12004_/B _12004_/C _12004_/Y vdd gnd OAI21X1
XFILL_2__7312_ vdd gnd FILL
X_10196_ _10196_/A _10196_/Y vdd gnd INVX1
XFILL_1__8519_ vdd gnd FILL
XFILL_1__9499_ vdd gnd FILL
XFILL_2__7243_ vdd gnd FILL
XFILL_1__11030_ vdd gnd FILL
XFILL_0__11760_ vdd gnd FILL
X_13955_ _13955_/A _13955_/B _13955_/C _13955_/Y vdd gnd OAI21X1
XFILL_2__12320_ vdd gnd FILL
XFILL_2__7174_ vdd gnd FILL
X_12906_ _12906_/A _12906_/B _12906_/C _12906_/Y vdd gnd OAI21X1
X_13886_ _13886_/A _13886_/B _13886_/C _13886_/Y vdd gnd OAI21X1
XFILL_2__12251_ vdd gnd FILL
XFILL_0__10642_ vdd gnd FILL
XFILL_1__12981_ vdd gnd FILL
X_12837_ _12837_/A _12837_/Y vdd gnd INVX1
XFILL_1__14720_ vdd gnd FILL
XFILL_1__11932_ vdd gnd FILL
XFILL_2__12182_ vdd gnd FILL
XFILL_0__13361_ vdd gnd FILL
XFILL_0__10573_ vdd gnd FILL
X_12768_ _12768_/A _12768_/Y vdd gnd INVX1
XFILL_0__12312_ vdd gnd FILL
XFILL_1__14651_ vdd gnd FILL
XFILL_1__11863_ vdd gnd FILL
X_14507_ _14507_/D _14507_/CLK _14507_/Q vdd gnd DFFPOSX1
XFILL_0__13292_ vdd gnd FILL
X_11719_ _11719_/A _11719_/Y vdd gnd INVX1
XFILL_1__10814_ vdd gnd FILL
X_12699_ _12699_/A _12699_/B _12699_/S _12699_/Y vdd gnd MUX2X1
XFILL_1__13602_ vdd gnd FILL
XFILL_1__14582_ vdd gnd FILL
XFILL_0__12243_ vdd gnd FILL
XFILL_1__11794_ vdd gnd FILL
XFILL_0__8830_ vdd gnd FILL
X_14438_ _14438_/A _14438_/B _14438_/Y vdd gnd NOR2X1
XFILL_2__10015_ vdd gnd FILL
XFILL_2__9746_ vdd gnd FILL
XFILL_1__13533_ vdd gnd FILL
XFILL_0__12174_ vdd gnd FILL
XFILL_0__8761_ vdd gnd FILL
X_14369_ _14369_/A _14369_/B _14369_/Y vdd gnd NOR2X1
XFILL_2__9677_ vdd gnd FILL
XFILL_0__11125_ vdd gnd FILL
XFILL_1__10676_ vdd gnd FILL
XFILL_0__7712_ vdd gnd FILL
XFILL_2_CLKBUF1_insert53 vdd gnd FILL
XFILL_0__8692_ vdd gnd FILL
XFILL_1__12415_ vdd gnd FILL
XFILL_2_CLKBUF1_insert75 vdd gnd FILL
XFILL_0__11056_ vdd gnd FILL
XFILL_2_CLKBUF1_insert86 vdd gnd FILL
XFILL_1__13395_ vdd gnd FILL
XFILL_0__7643_ vdd gnd FILL
XFILL_0__10007_ vdd gnd FILL
XFILL_1__12346_ vdd gnd FILL
XFILL_2__10917_ vdd gnd FILL
XFILL_0__7574_ vdd gnd FILL
XFILL_0__14815_ vdd gnd FILL
XFILL_1__12277_ vdd gnd FILL
XFILL_2__10848_ vdd gnd FILL
XFILL_0__9313_ vdd gnd FILL
X_9941_ _9941_/A _9941_/B _9941_/C _9941_/D _9941_/Y vdd gnd OAI22X1
XFILL_1__14016_ vdd gnd FILL
XFILL_1__11228_ vdd gnd FILL
XFILL_0_BUFX2_insert13 vdd gnd FILL
XFILL_0__14746_ vdd gnd FILL
XFILL_0_BUFX2_insert24 vdd gnd FILL
XFILL_2__10779_ vdd gnd FILL
XFILL_0__11958_ vdd gnd FILL
XFILL_0__9244_ vdd gnd FILL
X_9872_ _9872_/A _9872_/B _9872_/Y vdd gnd NAND2X1
XFILL_2__12518_ vdd gnd FILL
XFILL_0_CLKBUF1_insert90 vdd gnd FILL
XFILL_0__10909_ vdd gnd FILL
XFILL_1__11159_ vdd gnd FILL
XFILL_0__14677_ vdd gnd FILL
XFILL_0__9175_ vdd gnd FILL
XFILL_0__11889_ vdd gnd FILL
X_8823_ _8823_/A _8823_/B _8823_/C _8823_/Y vdd gnd OAI21X1
XFILL_0__13628_ vdd gnd FILL
XFILL_0__8126_ vdd gnd FILL
X_8754_ _8754_/A _8754_/B _8754_/C _8754_/Y vdd gnd OAI21X1
XFILL_1__14918_ vdd gnd FILL
XFILL_0__13559_ vdd gnd FILL
X_7705_ _7705_/A _7705_/B _7705_/Y vdd gnd NAND2X1
XFILL_0__8057_ vdd gnd FILL
X_8685_ _8685_/A _8685_/B _8685_/C _8685_/D _8685_/Y vdd gnd OAI22X1
XFILL_1__14849_ vdd gnd FILL
X_7636_ _7636_/A _7636_/B _7636_/Y vdd gnd OR2X2
XFILL_1__7821_ vdd gnd FILL
X_7567_ _7567_/A _7567_/B _7567_/Y vdd gnd NAND2X1
X_9306_ _9306_/A _9306_/B _9306_/Y vdd gnd NOR2X1
XFILL_0__8959_ vdd gnd FILL
XFILL_1__7752_ vdd gnd FILL
X_7498_ _7498_/A _7498_/B _7498_/C _7498_/Y vdd gnd AOI21X1
X_9237_ _9237_/A _9237_/B _9237_/Y vdd gnd AND2X2
XFILL_1__7683_ vdd gnd FILL
XFILL_1__9422_ vdd gnd FILL
X_9168_ _9168_/A _9168_/B _9168_/C _9168_/D _9168_/Y vdd gnd AOI22X1
X_10050_ _10050_/A _10050_/B _10050_/C _10050_/D _10050_/Y vdd gnd AOI22X1
X_8119_ _8119_/A _8119_/B _8119_/C _8119_/Y vdd gnd OAI21X1
XFILL_1__9353_ vdd gnd FILL
X_9099_ _9099_/A _9099_/B _9099_/C _9099_/Y vdd gnd AOI21X1
XFILL_1__8304_ vdd gnd FILL
XFILL_1__9284_ vdd gnd FILL
XFILL_1__8235_ vdd gnd FILL
X_13740_ _13740_/A _13740_/B _13740_/C _13740_/Y vdd gnd OAI21X1
X_10952_ _10952_/A _10952_/B _10952_/C _10952_/D _10952_/Y vdd gnd AOI22X1
XFILL_1__8166_ vdd gnd FILL
X_13671_ _13671_/A _13671_/B _13671_/C _13671_/Y vdd gnd AOI21X1
XFILL_1__7117_ vdd gnd FILL
XFILL_1__8097_ vdd gnd FILL
X_10883_ _10883_/A _10883_/B _10883_/C _10883_/Y vdd gnd NAND3X1
X_12622_ _12622_/A _12622_/B _12622_/Y vdd gnd AND2X2
X_12553_ _12553_/D _12553_/CLK _12553_/Q vdd gnd DFFPOSX1
XFILL_2__7861_ vdd gnd FILL
X_11504_ _11504_/A _11504_/B _11504_/Y vdd gnd NAND2X1
X_12484_ _12484_/A _12484_/B _12484_/Y vdd gnd NAND2X1
XFILL_1__8999_ vdd gnd FILL
X_14223_ _14223_/A _14223_/B _14223_/Y vdd gnd NAND2X1
X_11435_ _11435_/A _11435_/B _11435_/C _11435_/Y vdd gnd OAI21X1
XFILL_2__9531_ vdd gnd FILL
XFILL_1__10530_ vdd gnd FILL
X_11366_ _11366_/A _11366_/B _11366_/Y vdd gnd NAND2X1
X_14154_ _14154_/A _14154_/B _14154_/C _14154_/Y vdd gnd OAI21X1
XFILL_2__9462_ vdd gnd FILL
XFILL_1__10461_ vdd gnd FILL
X_13105_ _13105_/A _13105_/B _13105_/Y vdd gnd NOR2X1
X_10317_ _10317_/A _10317_/B _10317_/C _10317_/Y vdd gnd NAND3X1
XFILL_1__12200_ vdd gnd FILL
X_14085_ _14085_/A _14085_/B _14085_/Y vdd gnd AND2X2
X_11297_ _11297_/A _11297_/B _11297_/Y vdd gnd NAND2X1
XFILL_0__12930_ vdd gnd FILL
XFILL_1__13180_ vdd gnd FILL
XFILL_2__9393_ vdd gnd FILL
XFILL_1__10392_ vdd gnd FILL
X_10248_ _10248_/A _10248_/B _10248_/C _10248_/Y vdd gnd OAI21X1
X_13036_ _13036_/A _13036_/B _13036_/C _13036_/Y vdd gnd OAI21X1
XFILL_1__12131_ vdd gnd FILL
XFILL_0__12861_ vdd gnd FILL
X_10179_ _10179_/A _10179_/B _10179_/Y vdd gnd NAND2X1
XFILL_0__14600_ vdd gnd FILL
XFILL_1__12062_ vdd gnd FILL
XFILL_0__11812_ vdd gnd FILL
XFILL_0__12792_ vdd gnd FILL
XFILL_0__7290_ vdd gnd FILL
XFILL_1__11013_ vdd gnd FILL
XFILL_0__11743_ vdd gnd FILL
X_13938_ _13938_/A _13938_/B _13938_/Y vdd gnd NAND2X1
XFILL_2__12303_ vdd gnd FILL
XFILL_0__14462_ vdd gnd FILL
XFILL_2__12234_ vdd gnd FILL
X_13869_ _13869_/A _13869_/B _13869_/C _13869_/Y vdd gnd OAI21X1
XFILL_2__7088_ vdd gnd FILL
XFILL_0__13413_ vdd gnd FILL
XFILL_0__10625_ vdd gnd FILL
XFILL_1__12964_ vdd gnd FILL
XFILL_0__14393_ vdd gnd FILL
XFILL_1_BUFX2_insert360 vdd gnd FILL
XFILL_1_BUFX2_insert371 vdd gnd FILL
XFILL_1__14703_ vdd gnd FILL
XFILL_1_BUFX2_insert382 vdd gnd FILL
XFILL_2__12165_ vdd gnd FILL
XFILL_1__11915_ vdd gnd FILL
XFILL_0__13344_ vdd gnd FILL
XFILL_0__10556_ vdd gnd FILL
XFILL_1__12895_ vdd gnd FILL
XFILL_0__9931_ vdd gnd FILL
X_8470_ _8470_/A _8470_/B _8470_/Y vdd gnd NAND2X1
XFILL_1__14634_ vdd gnd FILL
XFILL_1__11846_ vdd gnd FILL
XFILL_2__12096_ vdd gnd FILL
XFILL_0__13275_ vdd gnd FILL
X_7421_ _7421_/A _7421_/Y vdd gnd INVX1
XFILL_0__10487_ vdd gnd FILL
XFILL_0__9862_ vdd gnd FILL
XFILL_0__12226_ vdd gnd FILL
XFILL_1__14565_ vdd gnd FILL
XFILL_1__11777_ vdd gnd FILL
XFILL_0__8813_ vdd gnd FILL
X_7352_ _7352_/A _7352_/B _7352_/C _7352_/Y vdd gnd OAI21X1
XFILL_2__9729_ vdd gnd FILL
XFILL_1__13516_ vdd gnd FILL
XFILL_0__12157_ vdd gnd FILL
XFILL_1__14496_ vdd gnd FILL
XFILL_0__8744_ vdd gnd FILL
X_7283_ _7283_/A _7283_/Y vdd gnd INVX1
XFILL_0__11108_ vdd gnd FILL
XFILL_1__10659_ vdd gnd FILL
X_9022_ _9022_/A _9022_/B _9022_/C _9022_/Y vdd gnd OAI21X1
XFILL_0__12088_ vdd gnd FILL
XFILL_2__12998_ vdd gnd FILL
XFILL_0__8675_ vdd gnd FILL
XFILL_0__11039_ vdd gnd FILL
XFILL_1__13378_ vdd gnd FILL
XFILL_0__7626_ vdd gnd FILL
XFILL_1__12329_ vdd gnd FILL
XFILL_0__7557_ vdd gnd FILL
X_9924_ _9924_/A _9924_/B _9924_/Y vdd gnd NAND2X1
XFILL_0__7488_ vdd gnd FILL
XFILL_0__14729_ vdd gnd FILL
XFILL_0__9227_ vdd gnd FILL
XFILL_1__8020_ vdd gnd FILL
X_9855_ _9855_/A _9855_/B _9855_/C _9855_/Y vdd gnd OAI21X1
XFILL_0__9158_ vdd gnd FILL
X_8806_ _8806_/A _8806_/B _8806_/C _8806_/Y vdd gnd OAI21X1
X_9786_ _9786_/D _9786_/CLK _9786_/Q vdd gnd DFFPOSX1
XFILL_0__8109_ vdd gnd FILL
XFILL_0__9089_ vdd gnd FILL
XFILL_1__9971_ vdd gnd FILL
X_8737_ _8737_/A _8737_/B _8737_/Y vdd gnd NAND2X1
XFILL_1__8922_ vdd gnd FILL
X_8668_ _8668_/A _8668_/B _8668_/C _8668_/Y vdd gnd AOI21X1
X_7619_ _7619_/A _7619_/B _7619_/C _7619_/Y vdd gnd OAI21X1
X_8599_ _8599_/A _8599_/B _8599_/Y vdd gnd NAND2X1
XFILL_1__7804_ vdd gnd FILL
XFILL_1__8784_ vdd gnd FILL
X_11220_ _11220_/A _11220_/B _11220_/Y vdd gnd NAND2X1
XFILL_1__7735_ vdd gnd FILL
X_11151_ _11151_/A _11151_/B _11151_/C _11151_/Y vdd gnd OAI21X1
XFILL_1__7666_ vdd gnd FILL
X_10102_ _10102_/A _10102_/Y vdd gnd INVX1
X_11082_ _11082_/A _11082_/B _11082_/C _11082_/Y vdd gnd NAND3X1
XFILL_1__9405_ vdd gnd FILL
XFILL_1__7597_ vdd gnd FILL
X_10033_ _10033_/A _10033_/B _10033_/C _10033_/Y vdd gnd OAI21X1
X_14910_ _14910_/A _14910_/Y vdd gnd BUFX2
XFILL_1__9336_ vdd gnd FILL
X_14841_ _14841_/A _14841_/Y vdd gnd INVX1
XFILL_1__9267_ vdd gnd FILL
XFILL_2__8060_ vdd gnd FILL
X_14772_ _14772_/A _14772_/Y vdd gnd INVX1
XFILL_1__8218_ vdd gnd FILL
X_11984_ _11984_/A _11984_/B _11984_/C _11984_/Y vdd gnd OAI21X1
XFILL_1__9198_ vdd gnd FILL
XFILL257550x75750 vdd gnd FILL
XFILL_0_BUFX2_insert5 vdd gnd FILL
X_13723_ _13723_/A _13723_/B _13723_/C _13723_/Y vdd gnd NAND3X1
X_10935_ _10935_/A _10935_/B _10935_/C _10935_/Y vdd gnd OAI21X1
XFILL_1__8149_ vdd gnd FILL
XFILL_2__10280_ vdd gnd FILL
X_13654_ _13654_/A _13654_/B _13654_/Y vdd gnd NAND2X1
X_10866_ _10866_/A _10866_/Y vdd gnd INVX1
XFILL_0__10410_ vdd gnd FILL
XFILL_2__8962_ vdd gnd FILL
X_12605_ _12605_/D _12605_/CLK _12605_/Q vdd gnd DFFPOSX1
XFILL_0__11390_ vdd gnd FILL
XFILL_0_BUFX2_insert301 vdd gnd FILL
XFILL_0_BUFX2_insert312 vdd gnd FILL
X_13585_ _13585_/A _13585_/Y vdd gnd INVX8
XFILL_0_BUFX2_insert323 vdd gnd FILL
XFILL_2__7913_ vdd gnd FILL
XFILL_1__11700_ vdd gnd FILL
XFILL_0_BUFX2_insert334 vdd gnd FILL
X_10797_ _10797_/A _10797_/B _10797_/C _10797_/Y vdd gnd OAI21X1
XFILL_0__10341_ vdd gnd FILL
XFILL_1__12680_ vdd gnd FILL
XFILL_0_BUFX2_insert345 vdd gnd FILL
XFILL_0_BUFX2_insert356 vdd gnd FILL
X_12536_ _12536_/D _12536_/CLK _12536_/Q vdd gnd DFFPOSX1
XFILL_0_BUFX2_insert367 vdd gnd FILL
XFILL_2__7844_ vdd gnd FILL
XFILL_0_BUFX2_insert378 vdd gnd FILL
XFILL_2__13970_ vdd gnd FILL
XFILL_0__13060_ vdd gnd FILL
XFILL_0__10272_ vdd gnd FILL
X_12467_ _12467_/A _12467_/B _12467_/Y vdd gnd NAND2X1
XFILL_0__12011_ vdd gnd FILL
XFILL_1__14350_ vdd gnd FILL
XFILL_2__7775_ vdd gnd FILL
XFILL_1__11562_ vdd gnd FILL
X_14206_ _14206_/D _14206_/CLK _14206_/Q vdd gnd DFFPOSX1
X_11418_ _11418_/A _11418_/B _11418_/Y vdd gnd NAND2X1
XFILL_1__13301_ vdd gnd FILL
XFILL_1__10513_ vdd gnd FILL
X_12398_ _12398_/A _12398_/B _12398_/Y vdd gnd NAND2X1
XFILL_1__14281_ vdd gnd FILL
XFILL_1__11493_ vdd gnd FILL
X_14137_ _14137_/A _14137_/B _14137_/C _14137_/Y vdd gnd OAI21X1
X_11349_ _11349_/A _11349_/B _11349_/C _11349_/Y vdd gnd OAI21X1
XFILL_2__11803_ vdd gnd FILL
XFILL_1__13232_ vdd gnd FILL
XFILL_1__10444_ vdd gnd FILL
XFILL_0__13962_ vdd gnd FILL
XFILL_2__12783_ vdd gnd FILL
XFILL_0__8460_ vdd gnd FILL
X_14068_ _14068_/A _14068_/Y vdd gnd INVX1
XFILL_1__13163_ vdd gnd FILL
XFILL_0__12913_ vdd gnd FILL
XFILL_2__9376_ vdd gnd FILL
XFILL_2__11734_ vdd gnd FILL
XFILL_1__10375_ vdd gnd FILL
XFILL_0__13893_ vdd gnd FILL
XFILL_0__7411_ vdd gnd FILL
X_13019_ _13019_/A _13019_/B _13019_/Y vdd gnd OR2X2
XFILL_2__8327_ vdd gnd FILL
XFILL_1__12114_ vdd gnd FILL
XFILL_0__8391_ vdd gnd FILL
XFILL_0__12844_ vdd gnd FILL
XFILL_1__13094_ vdd gnd FILL
XFILL_0__7342_ vdd gnd FILL
X_7970_ _7970_/D _7970_/CLK _7970_/Q vdd gnd DFFPOSX1
XFILL_2__10616_ vdd gnd FILL
XFILL_1__12045_ vdd gnd FILL
XFILL_2__11596_ vdd gnd FILL
XFILL_0__12775_ vdd gnd FILL
XFILL_0__7273_ vdd gnd FILL
XFILL_0__11726_ vdd gnd FILL
XFILL_0__9012_ vdd gnd FILL
X_9640_ _9640_/A _9640_/B _9640_/C _9640_/Y vdd gnd AOI21X1
XFILL_0__14445_ vdd gnd FILL
XFILL_1__13996_ vdd gnd FILL
X_9571_ _9571_/A _9571_/Y vdd gnd INVX1
XFILL_2__12217_ vdd gnd FILL
XFILL_0__10608_ vdd gnd FILL
XFILL_1__12947_ vdd gnd FILL
XFILL_0__14376_ vdd gnd FILL
XFILL_1_BUFX2_insert190 vdd gnd FILL
X_8522_ _8522_/A _8522_/B _8522_/C _8522_/Y vdd gnd OAI21X1
XFILL_0__11588_ vdd gnd FILL
XFILL_2__12148_ vdd gnd FILL
XFILL_0__13327_ vdd gnd FILL
XFILL_0__10539_ vdd gnd FILL
XFILL_0__9914_ vdd gnd FILL
XFILL_1__12878_ vdd gnd FILL
X_8453_ _8453_/A _8453_/B _8453_/C _8453_/Y vdd gnd AOI21X1
XFILL_2__12079_ vdd gnd FILL
XFILL_1__14617_ vdd gnd FILL
XFILL_1__11829_ vdd gnd FILL
XFILL_0__13258_ vdd gnd FILL
X_7404_ _7404_/A _7404_/B _7404_/Y vdd gnd AND2X2
XFILL_0__9845_ vdd gnd FILL
X_8384_ _8384_/A _8384_/B _8384_/C _8384_/Y vdd gnd OAI21X1
XFILL_0__12209_ vdd gnd FILL
XFILL_0__13189_ vdd gnd FILL
X_7335_ _7335_/A _7335_/Y vdd gnd INVX1
XFILL_1__14479_ vdd gnd FILL
XFILL_1__7520_ vdd gnd FILL
XFILL_0__8727_ vdd gnd FILL
X_7266_ _7266_/A _7266_/Y vdd gnd INVX2
X_9005_ _9005_/A _9005_/Y vdd gnd INVX8
XFILL_1__7451_ vdd gnd FILL
XFILL_0__8658_ vdd gnd FILL
X_7197_ _7197_/A _7197_/Y vdd gnd INVX1
XFILL_0__7609_ vdd gnd FILL
XFILL_1__7382_ vdd gnd FILL
XFILL_0__8589_ vdd gnd FILL
XFILL_1__9121_ vdd gnd FILL
X_9907_ _9907_/A _9907_/B _9907_/Y vdd gnd NAND2X1
XFILL_1__9052_ vdd gnd FILL
XFILL_1__8003_ vdd gnd FILL
X_9838_ _9838_/D _9838_/CLK _9838_/Q vdd gnd DFFPOSX1
X_10720_ _10720_/D _10720_/CLK _10720_/Q vdd gnd DFFPOSX1
X_9769_ _9769_/D _9769_/CLK _9769_/Q vdd gnd DFFPOSX1
X_10651_ _10651_/A _10651_/B _10651_/C _10651_/Y vdd gnd OAI21X1
XFILL_1__9954_ vdd gnd FILL
X_10582_ _10582_/A _10582_/B _10582_/C _10582_/Y vdd gnd AOI21X1
X_13370_ _13370_/A _13370_/B _13370_/C _13370_/Y vdd gnd OAI21X1
XFILL_1__9885_ vdd gnd FILL
X_12321_ _12321_/A _12321_/B _12321_/Y vdd gnd OR2X2
XFILL_1__8836_ vdd gnd FILL
X_12252_ _12252_/A _12252_/B _12252_/Y vdd gnd NAND2X1
XFILL_2__7560_ vdd gnd FILL
XFILL_1__8767_ vdd gnd FILL
XFILL257550x50550 vdd gnd FILL
X_11203_ _11203_/A _11203_/B _11203_/C _11203_/Y vdd gnd OAI21X1
X_12183_ _12183_/A _12183_/B _12183_/Y vdd gnd NAND2X1
XFILL_1__7718_ vdd gnd FILL
XFILL_2__7491_ vdd gnd FILL
XFILL_1__8698_ vdd gnd FILL
X_11134_ _11134_/A _11134_/B _11134_/Y vdd gnd NAND2X1
XFILL_1__7649_ vdd gnd FILL
X_11065_ _11065_/A _11065_/B _11065_/C _11065_/Y vdd gnd OAI21X1
XFILL_1__10160_ vdd gnd FILL
X_10016_ _10016_/A _10016_/B _10016_/C _10016_/D _10016_/Y vdd gnd AOI22X1
XFILL_0__10890_ vdd gnd FILL
XFILL_1__9319_ vdd gnd FILL
XFILL_2__8112_ vdd gnd FILL
XFILL_1__10091_ vdd gnd FILL
X_14824_ _14824_/A _14824_/B _14824_/Y vdd gnd NAND2X1
XFILL_2__10401_ vdd gnd FILL
XFILL_2__8043_ vdd gnd FILL
X_14755_ _14755_/A _14755_/B _14755_/C _14755_/Y vdd gnd AOI21X1
XFILL_2__10332_ vdd gnd FILL
X_11967_ _11967_/A _11967_/B _11967_/C _11967_/Y vdd gnd OAI21X1
XFILL_0__11511_ vdd gnd FILL
XFILL_1__13850_ vdd gnd FILL
XFILL_0__12491_ vdd gnd FILL
X_13706_ _13706_/A _13706_/B _13706_/C _13706_/Y vdd gnd AOI21X1
X_10918_ _10918_/A _10918_/Y vdd gnd INVX1
X_14686_ _14686_/A _14686_/Y vdd gnd INVX1
XFILL_2__10263_ vdd gnd FILL
XFILL_0__14230_ vdd gnd FILL
X_11898_ _11898_/A _11898_/B _11898_/C _11898_/D _11898_/Y vdd gnd AOI22X1
XFILL_1__12801_ vdd gnd FILL
XFILL_0__11442_ vdd gnd FILL
XFILL_1__10993_ vdd gnd FILL
XFILL_1__13781_ vdd gnd FILL
X_13637_ _13637_/A _13637_/B _13637_/Y vdd gnd OR2X2
X_10849_ _10849_/A _10849_/B _10849_/C _10849_/Y vdd gnd OAI21X1
XFILL_2__8945_ vdd gnd FILL
XFILL_2__10194_ vdd gnd FILL
XFILL_0_BUFX2_insert120 vdd gnd FILL
XFILL_1__12732_ vdd gnd FILL
XFILL_0__11373_ vdd gnd FILL
XFILL_0_BUFX2_insert131 vdd gnd FILL
XFILL_0_BUFX2_insert142 vdd gnd FILL
XFILL_0_BUFX2_insert153 vdd gnd FILL
X_13568_ _13568_/A _13568_/Y vdd gnd INVX2
XFILL_0__13112_ vdd gnd FILL
XFILL_1__12663_ vdd gnd FILL
XFILL_0__10324_ vdd gnd FILL
XFILL_0_BUFX2_insert164 vdd gnd FILL
XFILL_0_BUFX2_insert175 vdd gnd FILL
XFILL_0__14092_ vdd gnd FILL
XFILL_0_BUFX2_insert186 vdd gnd FILL
X_12519_ _12519_/A _12519_/B _12519_/C _12519_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert197 vdd gnd FILL
X_13499_ _13499_/D _13499_/CLK _13499_/Q vdd gnd DFFPOSX1
XFILL_0__7891_ vdd gnd FILL
XFILL_2__7827_ vdd gnd FILL
XFILL_1__14402_ vdd gnd FILL
XFILL_0__13043_ vdd gnd FILL
XFILL_0__10255_ vdd gnd FILL
XFILL_0__9630_ vdd gnd FILL
XFILL_2__7758_ vdd gnd FILL
XFILL_1__14333_ vdd gnd FILL
XFILL_1__11545_ vdd gnd FILL
X_7120_ _7120_/A _7120_/B _7120_/C _7120_/Y vdd gnd OAI21X1
XFILL_0__10186_ vdd gnd FILL
XFILL_0__9561_ vdd gnd FILL
XFILL_2__7689_ vdd gnd FILL
XFILL_1__14264_ vdd gnd FILL
XFILL_1__11476_ vdd gnd FILL
XFILL_0__8512_ vdd gnd FILL
XFILL_0__9492_ vdd gnd FILL
XFILL_1__13215_ vdd gnd FILL
XFILL_1__10427_ vdd gnd FILL
XFILL_0__13945_ vdd gnd FILL
XFILL_0__8443_ vdd gnd FILL
XFILL_1__13146_ vdd gnd FILL
XFILL_2__11717_ vdd gnd FILL
XFILL_1__10358_ vdd gnd FILL
XFILL_0__13876_ vdd gnd FILL
XFILL_0__8374_ vdd gnd FILL
XFILL_1__13077_ vdd gnd FILL
XFILL_1__10289_ vdd gnd FILL
XFILL_0__12827_ vdd gnd FILL
XFILL_0__7325_ vdd gnd FILL
X_7953_ _7953_/D _7953_/CLK _7953_/Q vdd gnd DFFPOSX1
XFILL_1__12028_ vdd gnd FILL
XFILL_0__12758_ vdd gnd FILL
XFILL_0__7256_ vdd gnd FILL
X_7884_ _7884_/A _7884_/B _7884_/C _7884_/Y vdd gnd OAI21X1
XFILL_0__11709_ vdd gnd FILL
XFILL_0__12689_ vdd gnd FILL
XFILL_0__7187_ vdd gnd FILL
X_9623_ _9623_/A _9623_/B _9623_/Y vdd gnd NAND2X1
XFILL_0__14428_ vdd gnd FILL
XFILL_1__13979_ vdd gnd FILL
X_9554_ _9554_/A _9554_/B _9554_/Y vdd gnd NAND2X1
XFILL_0__14359_ vdd gnd FILL
X_8505_ _8505_/A _8505_/B _8505_/Y vdd gnd NAND2X1
XBUFX2_insert15 BUFX2_insert15/A BUFX2_insert15/Y vdd gnd BUFX2
X_9485_ _9485_/A _9485_/B _9485_/C _9485_/Y vdd gnd OAI21X1
XBUFX2_insert26 BUFX2_insert26/A BUFX2_insert26/Y vdd gnd BUFX2
XFILL_1__9670_ vdd gnd FILL
X_8436_ _8436_/A _8436_/B _8436_/S _8436_/Y vdd gnd MUX2X1
XFILL_1__8621_ vdd gnd FILL
X_8367_ _8367_/A _8367_/B _8367_/Y vdd gnd NAND2X1
X_7318_ _7318_/A _7318_/B _7318_/C _7318_/Y vdd gnd AOI21X1
XFILL_0__9759_ vdd gnd FILL
XFILL_1__8552_ vdd gnd FILL
X_8298_ _8298_/A _8298_/B _8298_/C _8298_/Y vdd gnd NAND3X1
XFILL_1__7503_ vdd gnd FILL
X_7249_ _7249_/A _7249_/B _7249_/C _7249_/Y vdd gnd OAI21X1
XFILL_1__8483_ vdd gnd FILL
XFILL_1__7434_ vdd gnd FILL
XFILL_2_BUFX2_insert215 vdd gnd FILL
XFILL_1__7365_ vdd gnd FILL
XFILL_2_BUFX2_insert237 vdd gnd FILL
XFILL_1__9104_ vdd gnd FILL
X_12870_ _12870_/A _12870_/B _12870_/C _12870_/Y vdd gnd OAI21X1
XFILL_1__7296_ vdd gnd FILL
X_11821_ _11821_/A _11821_/B _11821_/Y vdd gnd OR2X2
XFILL_1__9035_ vdd gnd FILL
X_14540_ _14540_/D _14540_/CLK _14540_/Q vdd gnd DFFPOSX1
X_11752_ _11752_/A _11752_/Y vdd gnd INVX8
XFILL256950x198150 vdd gnd FILL
X_10703_ _10703_/D _10703_/CLK _10703_/Q vdd gnd DFFPOSX1
X_14471_ _14471_/A _14471_/B _14471_/C _14471_/Y vdd gnd OAI21X1
XBUFX2_insert203 BUFX2_insert203/A BUFX2_insert203/Y vdd gnd BUFX2
XBUFX2_insert214 BUFX2_insert214/A BUFX2_insert214/Y vdd gnd BUFX2
X_11683_ _11683_/D _11683_/CLK _11683_/Q vdd gnd DFFPOSX1
XBUFX2_insert225 BUFX2_insert225/A BUFX2_insert225/Y vdd gnd BUFX2
XBUFX2_insert236 BUFX2_insert236/A BUFX2_insert236/Y vdd gnd BUFX2
XBUFX2_insert247 BUFX2_insert247/A BUFX2_insert247/Y vdd gnd BUFX2
X_13422_ _13422_/A _13422_/B _13422_/C _13422_/Y vdd gnd OAI21X1
X_10634_ _10634_/A _10634_/B _10634_/Y vdd gnd NAND2X1
XFILL_1__9937_ vdd gnd FILL
XBUFX2_insert258 BUFX2_insert258/A BUFX2_insert258/Y vdd gnd BUFX2
XBUFX2_insert269 BUFX2_insert269/A BUFX2_insert269/Y vdd gnd BUFX2
X_13353_ _13353_/A _13353_/B _13353_/C _13353_/Y vdd gnd OAI21X1
X_10565_ _10565_/A _10565_/B _10565_/C _10565_/D _10565_/Y vdd gnd AOI22X1
XFILL_1__9868_ vdd gnd FILL
X_12304_ _12304_/A _12304_/B _12304_/C _12304_/Y vdd gnd OAI21X1
XFILL_1__8819_ vdd gnd FILL
X_13284_ _13284_/A _13284_/B _13284_/Y vdd gnd NAND2X1
X_10496_ _10496_/A _10496_/Y vdd gnd INVX1
XFILL_0__10040_ vdd gnd FILL
X_12235_ _12235_/A _12235_/B _12235_/Y vdd gnd NOR2X1
XFILL_1__11330_ vdd gnd FILL
XFILL_2__10881_ vdd gnd FILL
X_12166_ _12166_/A _12166_/B _12166_/Y vdd gnd NAND2X1
XFILL_2__7474_ vdd gnd FILL
XFILL_1__11261_ vdd gnd FILL
XFILL_0__11991_ vdd gnd FILL
X_11117_ _11117_/A _11117_/Y vdd gnd INVX1
XFILL_1__13000_ vdd gnd FILL
XFILL_1__10212_ vdd gnd FILL
X_12097_ _12097_/A _12097_/B _12097_/C _12097_/Y vdd gnd AOI21X1
XFILL_0__10942_ vdd gnd FILL
XFILL_0__13730_ vdd gnd FILL
XFILL_1__11192_ vdd gnd FILL
X_11048_ _11048_/A _11048_/B _11048_/C _11048_/Y vdd gnd OAI21X1
XFILL_1__10143_ vdd gnd FILL
XFILL_0__13661_ vdd gnd FILL
XFILL_2__12482_ vdd gnd FILL
XFILL_0__10873_ vdd gnd FILL
XFILL_1__10074_ vdd gnd FILL
XFILL_0__13592_ vdd gnd FILL
X_14807_ _14807_/A _14807_/B _14807_/C _14807_/Y vdd gnd OAI21X1
XFILL_0__7110_ vdd gnd FILL
XFILL_0__8090_ vdd gnd FILL
XFILL_2__8026_ vdd gnd FILL
X_12999_ _12999_/A _12999_/B _12999_/C _12999_/Y vdd gnd OAI21X1
XFILL_1__13902_ vdd gnd FILL
X_14738_ _14738_/A _14738_/Y vdd gnd INVX1
XFILL_2__13103_ vdd gnd FILL
XFILL_2__10315_ vdd gnd FILL
XFILL_1__13833_ vdd gnd FILL
XFILL_0__12474_ vdd gnd FILL
X_14669_ _14669_/A _14669_/B _14669_/Y vdd gnd NAND2X1
XFILL_2__13034_ vdd gnd FILL
XFILL_2__10246_ vdd gnd FILL
XFILL_0__11425_ vdd gnd FILL
XFILL_1__13764_ vdd gnd FILL
XFILL_1__10976_ vdd gnd FILL
XFILL_0__8992_ vdd gnd FILL
XFILL_2__8928_ vdd gnd FILL
XFILL_2__10177_ vdd gnd FILL
XFILL_1__12715_ vdd gnd FILL
XFILL_0__14144_ vdd gnd FILL
XFILL_0__11356_ vdd gnd FILL
XFILL_1__13695_ vdd gnd FILL
X_9270_ _9270_/A _9270_/B _9270_/Y vdd gnd NAND2X1
XFILL_0__10307_ vdd gnd FILL
XFILL_0__14075_ vdd gnd FILL
XFILL_1__12646_ vdd gnd FILL
X_8221_ _8221_/A _8221_/B _8221_/C _8221_/Y vdd gnd OAI21X1
XFILL_0__11287_ vdd gnd FILL
XFILL_0__7874_ vdd gnd FILL
XFILL_0__13026_ vdd gnd FILL
XFILL_0__10238_ vdd gnd FILL
XFILL_0__9613_ vdd gnd FILL
X_8152_ _8152_/A _8152_/Y vdd gnd INVX2
XFILL_1__14316_ vdd gnd FILL
XFILL_1__11528_ vdd gnd FILL
XFILL_0__10169_ vdd gnd FILL
X_7103_ _7103_/A _7103_/B _7103_/C _7103_/D _7103_/Y vdd gnd AOI22X1
XFILL_0__9544_ vdd gnd FILL
X_8083_ _8083_/A _8083_/B _8083_/Y vdd gnd NOR2X1
XFILL257550x248550 vdd gnd FILL
XFILL_1__14247_ vdd gnd FILL
XFILL_1__11459_ vdd gnd FILL
XFILL_0__9475_ vdd gnd FILL
XFILL_0__13928_ vdd gnd FILL
XFILL_0__8426_ vdd gnd FILL
XFILL_1__13129_ vdd gnd FILL
XFILL_0__13859_ vdd gnd FILL
XFILL_1__7150_ vdd gnd FILL
XFILL_0__8357_ vdd gnd FILL
X_8985_ _8985_/A _8985_/Y vdd gnd INVX1
XFILL_0__7308_ vdd gnd FILL
XFILL_1__7081_ vdd gnd FILL
X_7936_ _7936_/D _7936_/CLK _7936_/Q vdd gnd DFFPOSX1
XFILL_0__8288_ vdd gnd FILL
XFILL_0__7239_ vdd gnd FILL
X_7867_ _7867_/A _7867_/B _7867_/C _7867_/Y vdd gnd OAI21X1
X_9606_ _9606_/A _9606_/B _9606_/Y vdd gnd NOR2X1
X_7798_ _7798_/A _7798_/Y vdd gnd INVX1
X_9537_ _9537_/A _9537_/B _9537_/Y vdd gnd NAND2X1
XFILL_1__9722_ vdd gnd FILL
X_9468_ _9468_/A _9468_/B _9468_/Y vdd gnd NOR2X1
X_10350_ _10350_/A _10350_/B _10350_/C _10350_/Y vdd gnd NOR3X1
XFILL_1__9653_ vdd gnd FILL
X_8419_ _8419_/A _8419_/B _8419_/C _8419_/Y vdd gnd AOI21X1
X_9399_ _9399_/A _9399_/Y vdd gnd INVX1
X_10281_ _10281_/A _10281_/Y vdd gnd INVX1
XFILL_1__8604_ vdd gnd FILL
XFILL_1__9584_ vdd gnd FILL
X_12020_ _12020_/A _12020_/B _12020_/Y vdd gnd NAND2X1
XFILL_1__8535_ vdd gnd FILL
XFILL257550x158550 vdd gnd FILL
XFILL_1__8466_ vdd gnd FILL
X_13971_ _13971_/A _13971_/B _13971_/C _13971_/Y vdd gnd OAI21X1
XFILL_1__7417_ vdd gnd FILL
XFILL_1__8397_ vdd gnd FILL
X_12922_ _12922_/A _12922_/B _12922_/C _12922_/Y vdd gnd NAND3X1
XFILL_1__7348_ vdd gnd FILL
X_12853_ _12853_/A _12853_/B _12853_/C _12853_/Y vdd gnd OAI21X1
XFILL_1__7279_ vdd gnd FILL
X_11804_ _11804_/A _11804_/B _11804_/C _11804_/Y vdd gnd OAI21X1
XFILL_1__9018_ vdd gnd FILL
XFILL_2__9900_ vdd gnd FILL
X_12784_ _12784_/A _12784_/Y vdd gnd INVX1
XFILL257250x72150 vdd gnd FILL
X_14523_ _14523_/D _14523_/CLK _14523_/Q vdd gnd DFFPOSX1
X_11735_ _11735_/A _11735_/B _11735_/C _11735_/Y vdd gnd OAI21X1
XFILL_1__10830_ vdd gnd FILL
X_14454_ _14454_/A _14454_/B _14454_/C _14454_/Y vdd gnd OAI21X1
X_11666_ _11666_/D _11666_/CLK _11666_/Q vdd gnd DFFPOSX1
XFILL_0__11210_ vdd gnd FILL
XFILL_0__12190_ vdd gnd FILL
X_13405_ _13405_/A _13405_/B _13405_/C _13405_/Y vdd gnd OAI21X1
X_10617_ _10617_/A _10617_/B _10617_/C _10617_/Y vdd gnd OAI21X1
X_14385_ _14385_/A _14385_/Y vdd gnd INVX1
XFILL_2__8713_ vdd gnd FILL
XFILL_1__12500_ vdd gnd FILL
X_11597_ _11597_/A _11597_/B _11597_/C _11597_/Y vdd gnd OAI21X1
XFILL_2__9693_ vdd gnd FILL
XFILL_0__11141_ vdd gnd FILL
X_13336_ _13336_/A _13336_/B _13336_/C _13336_/Y vdd gnd AOI21X1
X_10548_ _10548_/A _10548_/Y vdd gnd INVX1
XFILL_2__8644_ vdd gnd FILL
XFILL_2__14770_ vdd gnd FILL
XFILL_1__12431_ vdd gnd FILL
XFILL_0__11072_ vdd gnd FILL
X_13267_ _13267_/A _13267_/B _13267_/C _13267_/Y vdd gnd OAI21X1
X_10479_ _10479_/A _10479_/B _10479_/C _10479_/Y vdd gnd OAI21X1
XFILL_0__10023_ vdd gnd FILL
XFILL_1__12362_ vdd gnd FILL
X_12218_ _12218_/A _12218_/B _12218_/C _12218_/Y vdd gnd OAI21X1
X_13198_ _13198_/A _13198_/Y vdd gnd INVX1
XFILL_0__7590_ vdd gnd FILL
XFILL_1__11313_ vdd gnd FILL
XFILL_1__14101_ vdd gnd FILL
XFILL_0__14831_ vdd gnd FILL
XFILL_1__12293_ vdd gnd FILL
X_12149_ _12149_/A _12149_/B _12149_/C _12149_/Y vdd gnd AOI21X1
XFILL_1__14032_ vdd gnd FILL
XFILL_1__11244_ vdd gnd FILL
XFILL_0__14762_ vdd gnd FILL
XFILL_0__11974_ vdd gnd FILL
XFILL_0__9260_ vdd gnd FILL
XFILL_2__12534_ vdd gnd FILL
XFILL_0__13713_ vdd gnd FILL
XFILL_0__10925_ vdd gnd FILL
XFILL_1__11175_ vdd gnd FILL
XFILL_0__8211_ vdd gnd FILL
XFILL_0__14693_ vdd gnd FILL
XFILL_0__9191_ vdd gnd FILL
XFILL_1__10126_ vdd gnd FILL
XFILL_2__12465_ vdd gnd FILL
XFILL_0__13644_ vdd gnd FILL
XFILL_0__10856_ vdd gnd FILL
XFILL_0__8142_ vdd gnd FILL
X_8770_ _8770_/A _8770_/B _8770_/Y vdd gnd NAND2X1
XFILL_1__10057_ vdd gnd FILL
XFILL_2__12396_ vdd gnd FILL
XFILL_0__13575_ vdd gnd FILL
XFILL_0__10787_ vdd gnd FILL
X_7721_ _7721_/A _7721_/B _7721_/Y vdd gnd NOR2X1
XFILL_0__8073_ vdd gnd FILL
XFILL_2__14135_ vdd gnd FILL
XFILL_0__12526_ vdd gnd FILL
XFILL_1__14865_ vdd gnd FILL
X_7652_ _7652_/A _7652_/B _7652_/C _7652_/Y vdd gnd OAI21X1
XFILL_2__14066_ vdd gnd FILL
XFILL_1__13816_ vdd gnd FILL
XFILL257550x223350 vdd gnd FILL
XFILL_0__12457_ vdd gnd FILL
XFILL_1__14796_ vdd gnd FILL
X_7583_ _7583_/A _7583_/B _7583_/C _7583_/Y vdd gnd NAND3X1
XFILL_2__13017_ vdd gnd FILL
XFILL_2__10229_ vdd gnd FILL
XFILL_0__11408_ vdd gnd FILL
XFILL_1__13747_ vdd gnd FILL
XFILL_1__10959_ vdd gnd FILL
XFILL_0__12388_ vdd gnd FILL
X_9322_ _9322_/A _9322_/B _9322_/S _9322_/Y vdd gnd MUX2X1
XFILL_0__8975_ vdd gnd FILL
XFILL_0__11339_ vdd gnd FILL
XFILL_0__14127_ vdd gnd FILL
XFILL_1__13678_ vdd gnd FILL
X_9253_ _9253_/A _9253_/B _9253_/Y vdd gnd NAND2X1
XFILL_0__14058_ vdd gnd FILL
XFILL_1__12629_ vdd gnd FILL
X_8204_ _8204_/A _8204_/Y vdd gnd INVX1
XFILL_0__7857_ vdd gnd FILL
X_9184_ _9184_/A _9184_/B _9184_/C _9184_/Y vdd gnd OAI21X1
XFILL_0__13009_ vdd gnd FILL
X_8135_ _8135_/A _8135_/B _8135_/S _8135_/Y vdd gnd MUX2X1
XFILL_0__7788_ vdd gnd FILL
XFILL_0__9527_ vdd gnd FILL
XFILL_1__8320_ vdd gnd FILL
X_8066_ _8066_/A _8066_/B _8066_/Y vdd gnd NAND2X1
XFILL_0__9458_ vdd gnd FILL
XFILL_1__8251_ vdd gnd FILL
XFILL_1__7202_ vdd gnd FILL
XFILL_0__8409_ vdd gnd FILL
XFILL_0__9389_ vdd gnd FILL
XFILL_1__8182_ vdd gnd FILL
XFILL_1__7133_ vdd gnd FILL
X_8968_ _8968_/A _8968_/B _8968_/C _8968_/Y vdd gnd OAI21X1
X_7919_ _7919_/D _7919_/CLK _7919_/Q vdd gnd DFFPOSX1
X_8899_ _8899_/D _8899_/CLK _8899_/Q vdd gnd DFFPOSX1
XFILL_0_CLKBUF1_insert101 vdd gnd FILL
XFILL257550x133350 vdd gnd FILL
X_11520_ _11520_/A _11520_/B _11520_/Y vdd gnd NAND2X1
X_11451_ _11451_/A _11451_/B _11451_/Y vdd gnd NAND2X1
X_10402_ _10402_/A _10402_/B _10402_/C _10402_/Y vdd gnd AOI21X1
XFILL_1__9705_ vdd gnd FILL
X_14170_ _14170_/D _14170_/CLK _14170_/Q vdd gnd DFFPOSX1
X_11382_ _11382_/A _11382_/B _11382_/C _11382_/Y vdd gnd OAI21X1
XFILL_1__7897_ vdd gnd FILL
X_13121_ _13121_/A _13121_/B _13121_/Y vdd gnd NAND2X1
X_10333_ _10333_/A _10333_/B _10333_/C _10333_/Y vdd gnd NAND3X1
XFILL_1__9636_ vdd gnd FILL
X_13052_ _13052_/A _13052_/B _13052_/Y vdd gnd NAND2X1
X_10264_ _10264_/A _10264_/B _10264_/Y vdd gnd NAND2X1
XFILL_1__9567_ vdd gnd FILL
XFILL_2__8360_ vdd gnd FILL
X_12003_ _12003_/A _12003_/Y vdd gnd INVX1
X_10195_ _10195_/A _10195_/B _10195_/Y vdd gnd NAND2X1
XFILL_1__8518_ vdd gnd FILL
XFILL_1__9498_ vdd gnd FILL
XFILL_2__8291_ vdd gnd FILL
XFILL_1__8449_ vdd gnd FILL
XFILL_2__10580_ vdd gnd FILL
X_13954_ _13954_/A _13954_/B _13954_/Y vdd gnd NOR2X1
X_12905_ _12905_/A _12905_/B _12905_/C _12905_/Y vdd gnd AOI21X1
X_13885_ _13885_/A _13885_/B _13885_/C _13885_/Y vdd gnd OAI21X1
XFILL_0__10641_ vdd gnd FILL
XFILL_1__12980_ vdd gnd FILL
X_12836_ _12836_/A _12836_/Y vdd gnd INVX1
XFILL_2__11201_ vdd gnd FILL
XFILL_1__11931_ vdd gnd FILL
XFILL_0__13360_ vdd gnd FILL
XFILL_0__10572_ vdd gnd FILL
X_12767_ _12767_/A _12767_/B _12767_/C _12767_/Y vdd gnd OAI21X1
XFILL_0__12311_ vdd gnd FILL
XFILL_2__11132_ vdd gnd FILL
XFILL_1__14650_ vdd gnd FILL
X_14506_ _14506_/D _14506_/CLK _14506_/Q vdd gnd DFFPOSX1
XFILL_1__11862_ vdd gnd FILL
XFILL_0__13291_ vdd gnd FILL
X_11718_ _11718_/A _11718_/B _11718_/C _11718_/Y vdd gnd AOI21X1
XFILL_1__13601_ vdd gnd FILL
X_12698_ _12698_/A _12698_/B _12698_/S _12698_/Y vdd gnd MUX2X1
XFILL_2__11063_ vdd gnd FILL
XFILL_0__12242_ vdd gnd FILL
XFILL_1__10813_ vdd gnd FILL
XFILL_1__14581_ vdd gnd FILL
XFILL_1__11793_ vdd gnd FILL
X_14437_ _14437_/A _14437_/B _14437_/Y vdd gnd NAND2X1
X_11649_ _11649_/D _11649_/CLK _11649_/Q vdd gnd DFFPOSX1
XFILL_1__13532_ vdd gnd FILL
XFILL_0__12173_ vdd gnd FILL
XFILL_0__8760_ vdd gnd FILL
X_14368_ _14368_/A _14368_/Y vdd gnd INVX1
XFILL_2__14822_ vdd gnd FILL
XFILL_0__11124_ vdd gnd FILL
XFILL_1__10675_ vdd gnd FILL
XFILL_2_CLKBUF1_insert32 vdd gnd FILL
XFILL_0__7711_ vdd gnd FILL
X_13319_ _13319_/A _13319_/B _13319_/C _13319_/Y vdd gnd AOI21X1
X_14299_ _14299_/A _14299_/B _14299_/Y vdd gnd NAND2X1
XFILL_0__8691_ vdd gnd FILL
XFILL_2__8627_ vdd gnd FILL
XFILL_2_CLKBUF1_insert65 vdd gnd FILL
XFILL_2__14753_ vdd gnd FILL
XFILL_1__12414_ vdd gnd FILL
XFILL_0__11055_ vdd gnd FILL
XFILL_2__11965_ vdd gnd FILL
XFILL_1__13394_ vdd gnd FILL
XFILL_0__7642_ vdd gnd FILL
XFILL_2_CLKBUF1_insert98 vdd gnd FILL
XFILL_0__10006_ vdd gnd FILL
XFILL_2__8558_ vdd gnd FILL
XFILL_2__14684_ vdd gnd FILL
XFILL_1__12345_ vdd gnd FILL
XFILL_2__11896_ vdd gnd FILL
XFILL_0__7573_ vdd gnd FILL
XFILL_0__14814_ vdd gnd FILL
XFILL_2__8489_ vdd gnd FILL
XFILL_0__9312_ vdd gnd FILL
XFILL_1__12276_ vdd gnd FILL
X_9940_ _9940_/A _9940_/B _9940_/C _9940_/Y vdd gnd NAND3X1
XFILL_1__14015_ vdd gnd FILL
XFILL_1__11227_ vdd gnd FILL
XFILL_0__14745_ vdd gnd FILL
XFILL_0_BUFX2_insert14 vdd gnd FILL
XFILL_0__9243_ vdd gnd FILL
XFILL_0__11957_ vdd gnd FILL
XFILL_0_BUFX2_insert25 vdd gnd FILL
XFILL_0_CLKBUF1_insert80 vdd gnd FILL
X_9871_ _9871_/A _9871_/Y vdd gnd INVX1
XFILL_0_CLKBUF1_insert91 vdd gnd FILL
XFILL_1__11158_ vdd gnd FILL
XFILL_0__10908_ vdd gnd FILL
XFILL_0__14676_ vdd gnd FILL
XFILL_0__9174_ vdd gnd FILL
XFILL_0__11888_ vdd gnd FILL
X_8822_ _8822_/A _8822_/B _8822_/C _8822_/Y vdd gnd OAI21X1
XFILL_1__10109_ vdd gnd FILL
XFILL_2__12448_ vdd gnd FILL
XFILL_0__13627_ vdd gnd FILL
XFILL_1__11089_ vdd gnd FILL
XFILL_0__8125_ vdd gnd FILL
XFILL_0__10839_ vdd gnd FILL
X_8753_ _8753_/A _8753_/B _8753_/Y vdd gnd NAND2X1
XFILL_1__14917_ vdd gnd FILL
XFILL_2__12379_ vdd gnd FILL
XFILL_0__13558_ vdd gnd FILL
X_7704_ _7704_/A _7704_/B _7704_/Y vdd gnd NOR2X1
XFILL_0__8056_ vdd gnd FILL
XFILL_2__14118_ vdd gnd FILL
X_8684_ _8684_/A _8684_/B _8684_/Y vdd gnd NAND2X1
XFILL_1__14848_ vdd gnd FILL
XFILL_0__12509_ vdd gnd FILL
X_7635_ _7635_/A _7635_/Y vdd gnd INVX1
XFILL_2__14049_ vdd gnd FILL
XFILL_1__14779_ vdd gnd FILL
XFILL_1__7820_ vdd gnd FILL
X_7566_ _7566_/A _7566_/B _7566_/C _7566_/Y vdd gnd NAND3X1
X_9305_ _9305_/A _9305_/B _9305_/Y vdd gnd NAND2X1
XFILL_0__8958_ vdd gnd FILL
XFILL_1__7751_ vdd gnd FILL
X_7497_ _7497_/A _7497_/B _7497_/C _7497_/Y vdd gnd NAND3X1
XFILL_0__7909_ vdd gnd FILL
X_9236_ _9236_/A _9236_/B _9236_/C _9236_/Y vdd gnd NAND3X1
XFILL_1__7682_ vdd gnd FILL
XFILL_1__9421_ vdd gnd FILL
X_9167_ _9167_/A _9167_/B _9167_/C _9167_/Y vdd gnd OAI21X1
XFILL_1__9352_ vdd gnd FILL
X_8118_ _8118_/A _8118_/B _8118_/S _8118_/Y vdd gnd MUX2X1
X_9098_ _9098_/A _9098_/B _9098_/C _9098_/Y vdd gnd NAND3X1
XFILL_1__8303_ vdd gnd FILL
XFILL_1__9283_ vdd gnd FILL
X_8049_ _8049_/A _8049_/B _8049_/C _8049_/Y vdd gnd OAI21X1
XFILL_1__8234_ vdd gnd FILL
X_10951_ _10951_/A _10951_/B _10951_/C _10951_/Y vdd gnd OAI21X1
XFILL_1__8165_ vdd gnd FILL
XFILL_1__7116_ vdd gnd FILL
X_13670_ _13670_/A _13670_/B _13670_/C _13670_/D _13670_/Y vdd gnd AOI22X1
X_10882_ _10882_/A _10882_/B _10882_/S _10882_/Y vdd gnd MUX2X1
XFILL_1__8096_ vdd gnd FILL
X_12621_ _12621_/A _12621_/Y vdd gnd INVX2
X_12552_ _12552_/D _12552_/CLK _12552_/Q vdd gnd DFFPOSX1
X_11503_ _11503_/A _11503_/B _11503_/Y vdd gnd NAND2X1
X_12483_ _12483_/A _12483_/B _12483_/C _12483_/Y vdd gnd OAI21X1
XFILL_1__8998_ vdd gnd FILL
XFILL_2__7791_ vdd gnd FILL
X_14222_ _14222_/A _14222_/Y vdd gnd INVX1
X_11434_ _11434_/A _11434_/B _11434_/C _11434_/Y vdd gnd AOI21X1
X_14153_ _14153_/A _14153_/B _14153_/Y vdd gnd NAND2X1
X_11365_ _11365_/A _11365_/B _11365_/C _11365_/Y vdd gnd OAI21X1
XFILL_1__10460_ vdd gnd FILL
X_13104_ _13104_/A _13104_/B _13104_/Y vdd gnd NAND2X1
X_10316_ _10316_/A _10316_/B _10316_/C _10316_/Y vdd gnd OAI21X1
XFILL_2__8412_ vdd gnd FILL
X_14084_ _14084_/A _14084_/B _14084_/Y vdd gnd NAND2X1
XFILL_1__9619_ vdd gnd FILL
X_11296_ _11296_/A _11296_/Y vdd gnd INVX1
XFILL_2__11750_ vdd gnd FILL
XFILL_1__10391_ vdd gnd FILL
X_13035_ _13035_/A _13035_/B _13035_/C _13035_/Y vdd gnd AOI21X1
X_10247_ _10247_/A _10247_/B _10247_/S _10247_/Y vdd gnd MUX2X1
XFILL_2__8343_ vdd gnd FILL
XFILL_1__12130_ vdd gnd FILL
XFILL_0__12860_ vdd gnd FILL
X_10178_ _10178_/A _10178_/B _10178_/C _10178_/Y vdd gnd NAND3X1
XFILL_2__13420_ vdd gnd FILL
XFILL_2__10632_ vdd gnd FILL
XFILL_2__8274_ vdd gnd FILL
XFILL_1__12061_ vdd gnd FILL
XFILL_0__11811_ vdd gnd FILL
XFILL_0__12791_ vdd gnd FILL
XFILL_1__11012_ vdd gnd FILL
XFILL_2__13351_ vdd gnd FILL
XFILL_2__10563_ vdd gnd FILL
XFILL_0__11742_ vdd gnd FILL
X_13937_ _13937_/A _13937_/B _13937_/C _13937_/Y vdd gnd NAND3X1
XFILL_2__13282_ vdd gnd FILL
XFILL_2__10494_ vdd gnd FILL
XFILL_0__14461_ vdd gnd FILL
X_13868_ _13868_/A _13868_/B _13868_/C _13868_/Y vdd gnd OAI21X1
XFILL_0__10624_ vdd gnd FILL
XFILL_0__13412_ vdd gnd FILL
XFILL_1__12963_ vdd gnd FILL
XFILL_0__14392_ vdd gnd FILL
XFILL_1_BUFX2_insert350 vdd gnd FILL
X_12819_ _12819_/A _12819_/B _12819_/Y vdd gnd NAND2X1
XFILL_1__14702_ vdd gnd FILL
XFILL_1_BUFX2_insert361 vdd gnd FILL
X_13799_ _13799_/A _13799_/B _13799_/C _13799_/Y vdd gnd NAND3X1
XFILL_1_BUFX2_insert372 vdd gnd FILL
XFILL_1__11914_ vdd gnd FILL
XFILL_0__10555_ vdd gnd FILL
XFILL_1_BUFX2_insert383 vdd gnd FILL
XFILL_0__13343_ vdd gnd FILL
XFILL_0__9930_ vdd gnd FILL
XFILL_1__12894_ vdd gnd FILL
XFILL256350x219750 vdd gnd FILL
XFILL_2__11115_ vdd gnd FILL
XFILL_1__14633_ vdd gnd FILL
XFILL_1__11845_ vdd gnd FILL
XFILL_0__13274_ vdd gnd FILL
XFILL_0__10486_ vdd gnd FILL
X_7420_ _7420_/A _7420_/B _7420_/Y vdd gnd NAND2X1
XFILL_0__9861_ vdd gnd FILL
XFILL_0__12225_ vdd gnd FILL
XFILL_2__11046_ vdd gnd FILL
XFILL_1__14564_ vdd gnd FILL
XFILL_1__11776_ vdd gnd FILL
XFILL_0__8812_ vdd gnd FILL
X_7351_ _7351_/A _7351_/Y vdd gnd INVX1
XFILL_1__13515_ vdd gnd FILL
XFILL_0__12156_ vdd gnd FILL
XFILL_1__14495_ vdd gnd FILL
XFILL_0__8743_ vdd gnd FILL
X_7282_ _7282_/A _7282_/B _7282_/Y vdd gnd NAND2X1
XFILL_2__14805_ vdd gnd FILL
XFILL_0__11107_ vdd gnd FILL
XFILL_1__10658_ vdd gnd FILL
XFILL_0__12087_ vdd gnd FILL
X_9021_ _9021_/A _9021_/B _9021_/Y vdd gnd NAND2X1
XFILL_0__8674_ vdd gnd FILL
XFILL_2__14736_ vdd gnd FILL
XFILL_0__11038_ vdd gnd FILL
XFILL_2__11948_ vdd gnd FILL
XFILL_1__13377_ vdd gnd FILL
XFILL_0__7625_ vdd gnd FILL
XFILL_1__10589_ vdd gnd FILL
XFILL_2__14667_ vdd gnd FILL
XFILL_1__12328_ vdd gnd FILL
XFILL_2__11879_ vdd gnd FILL
XFILL_0__7556_ vdd gnd FILL
XFILL_2__13618_ vdd gnd FILL
XFILL_2__14598_ vdd gnd FILL
XFILL_1__12259_ vdd gnd FILL
X_9923_ _9923_/A _9923_/Y vdd gnd INVX1
XFILL_0__12989_ vdd gnd FILL
XFILL_0__7487_ vdd gnd FILL
XFILL_2__13549_ vdd gnd FILL
XFILL_0__14728_ vdd gnd FILL
XFILL_0__9226_ vdd gnd FILL
X_9854_ _9854_/A _9854_/B _9854_/C _9854_/D _9854_/Y vdd gnd AOI22X1
XFILL_0__14659_ vdd gnd FILL
XFILL_0__9157_ vdd gnd FILL
X_8805_ _8805_/A _8805_/B _8805_/C _8805_/Y vdd gnd OAI21X1
X_9785_ _9785_/D _9785_/CLK _9785_/Q vdd gnd DFFPOSX1
XFILL_0__8108_ vdd gnd FILL
XFILL_0__9088_ vdd gnd FILL
XFILL_1__9970_ vdd gnd FILL
X_8736_ _8736_/A _8736_/B _8736_/Y vdd gnd NAND2X1
XFILL_1__8921_ vdd gnd FILL
XFILL_0__8039_ vdd gnd FILL
X_8667_ _8667_/A _8667_/B _8667_/Y vdd gnd NAND2X1
X_7618_ _7618_/A _7618_/B _7618_/C _7618_/D _7618_/Y vdd gnd AOI22X1
X_8598_ _8598_/A _8598_/B _8598_/C _8598_/D _8598_/Y vdd gnd AOI22X1
XFILL_1__7803_ vdd gnd FILL
X_7549_ _7549_/A _7549_/B _7549_/Y vdd gnd NAND2X1
XFILL_1__8783_ vdd gnd FILL
XFILL_1__7734_ vdd gnd FILL
X_11150_ _11150_/A _11150_/B _11150_/C _11150_/Y vdd gnd OAI21X1
X_9219_ _9219_/A _9219_/B _9219_/Y vdd gnd NAND2X1
XFILL_1__7665_ vdd gnd FILL
X_10101_ _10101_/A _10101_/B _10101_/C _10101_/Y vdd gnd NAND3X1
XFILL_1__9404_ vdd gnd FILL
X_11081_ _11081_/A _11081_/B _11081_/C _11081_/Y vdd gnd NAND3X1
XFILL_1__7596_ vdd gnd FILL
X_10032_ _10032_/A _10032_/B _10032_/Y vdd gnd NAND2X1
XFILL_1__9335_ vdd gnd FILL
X_14840_ _14840_/A _14840_/B _14840_/C _14840_/Y vdd gnd AOI21X1
XFILL_1__9266_ vdd gnd FILL
X_14771_ _14771_/A _14771_/B _14771_/Y vdd gnd NAND2X1
XFILL_1__8217_ vdd gnd FILL
X_11983_ _11983_/A _11983_/B _11983_/C _11983_/Y vdd gnd NAND3X1
XFILL_1__9197_ vdd gnd FILL
X_13722_ _13722_/A _13722_/B _13722_/Y vdd gnd NAND2X1
X_10934_ _10934_/A _10934_/B _10934_/Y vdd gnd NAND2X1
XFILL_0_BUFX2_insert6 vdd gnd FILL
XFILL_1__8148_ vdd gnd FILL
X_13653_ _13653_/A _13653_/B _13653_/C _13653_/Y vdd gnd OAI21X1
X_10865_ _10865_/A _10865_/B _10865_/C _10865_/D _10865_/Y vdd gnd OAI22X1
XFILL_1__8079_ vdd gnd FILL
X_12604_ _12604_/D _12604_/CLK _12604_/Q vdd gnd DFFPOSX1
XFILL_0_BUFX2_insert302 vdd gnd FILL
X_13584_ _13584_/A _13584_/Y vdd gnd INVX1
XFILL_0_BUFX2_insert313 vdd gnd FILL
X_10796_ _10796_/A _10796_/B _10796_/Y vdd gnd NAND2X1
XFILL_0__10340_ vdd gnd FILL
XFILL_0_BUFX2_insert324 vdd gnd FILL
XFILL_0_BUFX2_insert335 vdd gnd FILL
X_12535_ _12535_/A _12535_/B _12535_/C _12535_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert346 vdd gnd FILL
XFILL_0_BUFX2_insert357 vdd gnd FILL
XFILL_0_BUFX2_insert368 vdd gnd FILL
XFILL_0__10271_ vdd gnd FILL
XFILL_0_BUFX2_insert379 vdd gnd FILL
X_12466_ _12466_/A _12466_/B _12466_/Y vdd gnd NAND2X1
XFILL_0__12010_ vdd gnd FILL
X_14205_ _14205_/D _14205_/CLK _14205_/Q vdd gnd DFFPOSX1
XFILL_1__11561_ vdd gnd FILL
X_11417_ _11417_/A _11417_/B _11417_/Y vdd gnd NOR2X1
X_12397_ _12397_/A _12397_/B _12397_/Y vdd gnd NOR2X1
XFILL_1__13300_ vdd gnd FILL
XFILL_1__10512_ vdd gnd FILL
XFILL_1__14280_ vdd gnd FILL
XFILL_1__11492_ vdd gnd FILL
X_14136_ _14136_/A _14136_/B _14136_/C _14136_/Y vdd gnd OAI21X1
X_11348_ _11348_/A _11348_/B _11348_/C _11348_/Y vdd gnd OAI21X1
XFILL_1__13231_ vdd gnd FILL
XFILL_1__10443_ vdd gnd FILL
XFILL_0__13961_ vdd gnd FILL
X_14067_ _14067_/A _14067_/B _14067_/C _14067_/Y vdd gnd OAI21X1
X_11279_ _11279_/A _11279_/B _11279_/C _11279_/Y vdd gnd NAND3X1
XFILL_1__13162_ vdd gnd FILL
XFILL_1__10374_ vdd gnd FILL
XFILL_0__12912_ vdd gnd FILL
XFILL_0__7410_ vdd gnd FILL
X_13018_ _13018_/A _13018_/B _13018_/Y vdd gnd NAND2X1
XFILL_0__13892_ vdd gnd FILL
XFILL_0__8390_ vdd gnd FILL
XFILL_1__12113_ vdd gnd FILL
XFILL_2__14452_ vdd gnd FILL
XFILL_0__12843_ vdd gnd FILL
XFILL_1__13093_ vdd gnd FILL
XFILL_0__7341_ vdd gnd FILL
XFILL_2__13403_ vdd gnd FILL
XFILL_2__8257_ vdd gnd FILL
XFILL_1__12044_ vdd gnd FILL
XFILL_0__12774_ vdd gnd FILL
XFILL_2__7208_ vdd gnd FILL
XFILL_0__7272_ vdd gnd FILL
XFILL_2__13334_ vdd gnd FILL
XFILL_2__10546_ vdd gnd FILL
XFILL_2__8188_ vdd gnd FILL
XFILL_0__9011_ vdd gnd FILL
XFILL_0__11725_ vdd gnd FILL
XFILL_2__13265_ vdd gnd FILL
XFILL_2__10477_ vdd gnd FILL
XFILL_0__14444_ vdd gnd FILL
XFILL_1__13995_ vdd gnd FILL
X_9570_ _9570_/A _9570_/B _9570_/Y vdd gnd NAND2X1
XFILL_2__13196_ vdd gnd FILL
XFILL_1__12946_ vdd gnd FILL
XFILL_0__10607_ vdd gnd FILL
XFILL_0__14375_ vdd gnd FILL
XFILL_0__11587_ vdd gnd FILL
XFILL_1_BUFX2_insert180 vdd gnd FILL
X_8521_ _8521_/A _8521_/B _8521_/Y vdd gnd NAND2X1
XFILL_1_BUFX2_insert191 vdd gnd FILL
XFILL_0__10538_ vdd gnd FILL
XFILL_0__13326_ vdd gnd FILL
XFILL_1__12877_ vdd gnd FILL
XFILL_0__9913_ vdd gnd FILL
X_8452_ _8452_/A _8452_/B _8452_/C _8452_/D _8452_/Y vdd gnd AOI22X1
XFILL_1__14616_ vdd gnd FILL
XFILL_1__11828_ vdd gnd FILL
XFILL_0__10469_ vdd gnd FILL
XFILL_0__13257_ vdd gnd FILL
X_7403_ _7403_/A _7403_/Y vdd gnd INVX1
XFILL_0__9844_ vdd gnd FILL
XFILL_2__11029_ vdd gnd FILL
X_8383_ _8383_/A _8383_/B _8383_/Y vdd gnd NAND2X1
XFILL_0__12208_ vdd gnd FILL
XFILL_0__13188_ vdd gnd FILL
XFILL_1__11759_ vdd gnd FILL
X_7334_ _7334_/A _7334_/B _7334_/C _7334_/Y vdd gnd NAND3X1
XFILL_0__12139_ vdd gnd FILL
XFILL_1__14478_ vdd gnd FILL
XFILL_0__8726_ vdd gnd FILL
X_7265_ _7265_/A _7265_/B _7265_/C _7265_/Y vdd gnd OAI21X1
X_9004_ _9004_/A _9004_/B _9004_/C _9004_/Y vdd gnd OAI21X1
XFILL_1__7450_ vdd gnd FILL
XFILL_0__8657_ vdd gnd FILL
X_7196_ _7196_/A _7196_/B _7196_/C _7196_/Y vdd gnd AOI21X1
XFILL_0__7608_ vdd gnd FILL
XFILL_1__7381_ vdd gnd FILL
XFILL_0__8588_ vdd gnd FILL
XFILL_1__9120_ vdd gnd FILL
XFILL_0__7539_ vdd gnd FILL
XFILL_1__9051_ vdd gnd FILL
X_9906_ _9906_/A _9906_/Y vdd gnd INVX1
XFILL_0__9209_ vdd gnd FILL
XFILL_1__8002_ vdd gnd FILL
X_9837_ _9837_/D _9837_/CLK _9837_/Q vdd gnd DFFPOSX1
X_9768_ _9768_/D _9768_/CLK _9768_/Q vdd gnd DFFPOSX1
X_10650_ _10650_/A _10650_/B _10650_/Y vdd gnd NAND2X1
X_8719_ _8719_/A _8719_/B _8719_/Y vdd gnd NOR2X1
XFILL_1__9953_ vdd gnd FILL
X_9699_ _9699_/A _9699_/B _9699_/Y vdd gnd AND2X2
X_10581_ _10581_/A _10581_/B _10581_/C _10581_/Y vdd gnd OAI21X1
XFILL_1__9884_ vdd gnd FILL
X_12320_ _12320_/A _12320_/B _12320_/Y vdd gnd OR2X2
XFILL_1__8835_ vdd gnd FILL
X_12251_ _12251_/A _12251_/B _12251_/C _12251_/Y vdd gnd NAND3X1
XFILL257250x169350 vdd gnd FILL
XFILL_1__8766_ vdd gnd FILL
X_11202_ _11202_/A _11202_/B _11202_/C _11202_/Y vdd gnd OAI21X1
XFILL_1__7717_ vdd gnd FILL
X_12182_ _12182_/A _12182_/B _12182_/C _12182_/Y vdd gnd OAI21X1
XFILL_1__8697_ vdd gnd FILL
X_11133_ _11133_/A _11133_/B _11133_/C _11133_/Y vdd gnd OAI21X1
XFILL_1__7648_ vdd gnd FILL
X_11064_ _11064_/A _11064_/B _11064_/C _11064_/Y vdd gnd AOI21X1
XFILL_2__9160_ vdd gnd FILL
XFILL_1__7579_ vdd gnd FILL
X_10015_ _10015_/A _10015_/B _10015_/Y vdd gnd NOR2X1
XFILL_1__9318_ vdd gnd FILL
XFILL_2__9091_ vdd gnd FILL
XFILL_1__10090_ vdd gnd FILL
X_14823_ _14823_/A _14823_/B _14823_/Y vdd gnd NOR2X1
XFILL_1__9249_ vdd gnd FILL
X_14754_ _14754_/A _14754_/B _14754_/Y vdd gnd OR2X2
X_11966_ _11966_/A _11966_/B _11966_/C _11966_/Y vdd gnd OAI21X1
XFILL_0__11510_ vdd gnd FILL
XFILL_0__12490_ vdd gnd FILL
X_10917_ _10917_/A _10917_/B _10917_/C _10917_/Y vdd gnd NAND3X1
X_13705_ _13705_/A _13705_/B _13705_/C _13705_/Y vdd gnd NAND3X1
X_14685_ _14685_/A _14685_/B _14685_/Y vdd gnd NOR2X1
X_11897_ _11897_/A _11897_/B _11897_/C _11897_/Y vdd gnd OAI21X1
XFILL_1__12800_ vdd gnd FILL
XFILL_2__13050_ vdd gnd FILL
XFILL_0__11441_ vdd gnd FILL
XFILL_2__9993_ vdd gnd FILL
XFILL_1__13780_ vdd gnd FILL
X_13636_ _13636_/A _13636_/Y vdd gnd INVX1
XFILL_1__10992_ vdd gnd FILL
X_10848_ _10848_/A _10848_/B _10848_/Y vdd gnd NAND2X1
XFILL_0_BUFX2_insert110 vdd gnd FILL
XFILL_1__12731_ vdd gnd FILL
XFILL_0_BUFX2_insert121 vdd gnd FILL
XFILL_0__11372_ vdd gnd FILL
X_13567_ _13567_/A _13567_/B _13567_/C _13567_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert132 vdd gnd FILL
XFILL_0_BUFX2_insert143 vdd gnd FILL
X_10779_ _10779_/A _10779_/B _10779_/C _10779_/Y vdd gnd OAI21X1
XFILL_0__10323_ vdd gnd FILL
XFILL_0_BUFX2_insert154 vdd gnd FILL
XFILL_0__13111_ vdd gnd FILL
XFILL_1__12662_ vdd gnd FILL
XFILL_0_BUFX2_insert165 vdd gnd FILL
XFILL_0__14091_ vdd gnd FILL
XFILL_0_BUFX2_insert176 vdd gnd FILL
X_12518_ _12518_/A _12518_/B _12518_/C _12518_/Y vdd gnd OAI21X1
X_13498_ _13498_/D _13498_/CLK _13498_/Q vdd gnd DFFPOSX1
XFILL_0__7890_ vdd gnd FILL
XFILL_0_BUFX2_insert187 vdd gnd FILL
XFILL_1__14401_ vdd gnd FILL
XFILL_0__13042_ vdd gnd FILL
XFILL_0_BUFX2_insert198 vdd gnd FILL
XFILL_0__10254_ vdd gnd FILL
X_12449_ _12449_/A _12449_/B _12449_/Y vdd gnd NAND2X1
XFILL_2__12903_ vdd gnd FILL
XFILL_1__14332_ vdd gnd FILL
XFILL_1__11544_ vdd gnd FILL
XFILL_0__10185_ vdd gnd FILL
XFILL_0__9560_ vdd gnd FILL
XFILL_1_CLKBUF1_insert390 vdd gnd FILL
XFILL_2__12834_ vdd gnd FILL
XFILL_1__14263_ vdd gnd FILL
XFILL_0__8511_ vdd gnd FILL
XFILL_1__11475_ vdd gnd FILL
X_14119_ _14119_/A _14119_/B _14119_/Y vdd gnd NAND2X1
XFILL_0__9491_ vdd gnd FILL
XFILL_1__13214_ vdd gnd FILL
XFILL_2__9427_ vdd gnd FILL
XFILL_1__10426_ vdd gnd FILL
XFILL_0__13944_ vdd gnd FILL
XFILL_0__8442_ vdd gnd FILL
XFILL_1__13145_ vdd gnd FILL
XFILL_1__10357_ vdd gnd FILL
XFILL_0__13875_ vdd gnd FILL
XFILL_0__8373_ vdd gnd FILL
XFILL_2__14435_ vdd gnd FILL
XFILL_1__13076_ vdd gnd FILL
XFILL_1__10288_ vdd gnd FILL
XFILL_0__12826_ vdd gnd FILL
XFILL_0__7324_ vdd gnd FILL
X_7952_ _7952_/D _7952_/CLK _7952_/Q vdd gnd DFFPOSX1
XFILL_1__12027_ vdd gnd FILL
XFILL_2__14366_ vdd gnd FILL
XFILL257250x234150 vdd gnd FILL
XFILL_0__12757_ vdd gnd FILL
XFILL_0__7255_ vdd gnd FILL
XFILL_2__13317_ vdd gnd FILL
X_7883_ _7883_/A _7883_/B _7883_/C _7883_/Y vdd gnd OAI21X1
XFILL_2__14297_ vdd gnd FILL
XFILL_0__11708_ vdd gnd FILL
X_9622_ _9622_/A _9622_/B _9622_/Y vdd gnd OR2X2
XFILL_0__12688_ vdd gnd FILL
XFILL_0__7186_ vdd gnd FILL
XFILL_2__13248_ vdd gnd FILL
XFILL_0__14427_ vdd gnd FILL
XFILL_1__13978_ vdd gnd FILL
X_9553_ _9553_/A _9553_/B _9553_/Y vdd gnd NAND2X1
XFILL_1__12929_ vdd gnd FILL
XFILL_2__13179_ vdd gnd FILL
XFILL_0__14358_ vdd gnd FILL
X_8504_ _8504_/A _8504_/B _8504_/C _8504_/Y vdd gnd OAI21X1
X_9484_ _9484_/A _9484_/B _9484_/Y vdd gnd OR2X2
XBUFX2_insert16 BUFX2_insert16/A BUFX2_insert16/Y vdd gnd BUFX2
XFILL_0__13309_ vdd gnd FILL
XBUFX2_insert27 BUFX2_insert27/A BUFX2_insert27/Y vdd gnd BUFX2
XFILL_0__14289_ vdd gnd FILL
X_8435_ _8435_/A _8435_/B _8435_/C _8435_/Y vdd gnd OAI21X1
XFILL_1__8620_ vdd gnd FILL
X_8366_ _8366_/A _8366_/B _8366_/C _8366_/Y vdd gnd NAND3X1
X_7317_ _7317_/A _7317_/B _7317_/Y vdd gnd NAND2X1
XFILL_1__8551_ vdd gnd FILL
XFILL_0__9758_ vdd gnd FILL
X_8297_ _8297_/A _8297_/B _8297_/Y vdd gnd AND2X2
XFILL_1__7502_ vdd gnd FILL
XFILL_0__8709_ vdd gnd FILL
X_7248_ _7248_/A _7248_/Y vdd gnd INVX1
XFILL_0__9689_ vdd gnd FILL
XFILL_1__8482_ vdd gnd FILL
XFILL_1__7433_ vdd gnd FILL
X_7179_ _7179_/A _7179_/Y vdd gnd INVX1
XFILL_1__7364_ vdd gnd FILL
XFILL_2_BUFX2_insert227 vdd gnd FILL
XFILL_1__9103_ vdd gnd FILL
XFILL_2_BUFX2_insert249 vdd gnd FILL
XFILL_1__7295_ vdd gnd FILL
X_11820_ _11820_/A _11820_/B _11820_/C _11820_/Y vdd gnd OAI21X1
XFILL_1__9034_ vdd gnd FILL
XFILL257250x144150 vdd gnd FILL
X_11751_ _11751_/A _11751_/Y vdd gnd INVX1
X_10702_ _10702_/D _10702_/CLK _10702_/Q vdd gnd DFFPOSX1
X_14470_ _14470_/A _14470_/B _14470_/Y vdd gnd NAND2X1
XBUFX2_insert204 BUFX2_insert204/A BUFX2_insert204/Y vdd gnd BUFX2
X_11682_ _11682_/D _11682_/CLK _11682_/Q vdd gnd DFFPOSX1
XBUFX2_insert215 BUFX2_insert215/A BUFX2_insert215/Y vdd gnd BUFX2
X_13421_ _13421_/A _13421_/B _13421_/C _13421_/Y vdd gnd OAI21X1
XBUFX2_insert226 BUFX2_insert226/A BUFX2_insert226/Y vdd gnd BUFX2
XBUFX2_insert237 BUFX2_insert237/A BUFX2_insert237/Y vdd gnd BUFX2
X_10633_ _10633_/A _10633_/B _10633_/C _10633_/Y vdd gnd OAI21X1
XBUFX2_insert248 BUFX2_insert248/A BUFX2_insert248/Y vdd gnd BUFX2
XFILL_1__9936_ vdd gnd FILL
XBUFX2_insert259 BUFX2_insert259/A BUFX2_insert259/Y vdd gnd BUFX2
X_13352_ _13352_/A _13352_/B _13352_/Y vdd gnd OR2X2
X_10564_ _10564_/A _10564_/B _10564_/C _10564_/Y vdd gnd AOI21X1
XFILL_2__8660_ vdd gnd FILL
XFILL_1__9867_ vdd gnd FILL
X_12303_ _12303_/A _12303_/B _12303_/C _12303_/Y vdd gnd OAI21X1
X_13283_ _13283_/A _13283_/B _13283_/Y vdd gnd NOR2X1
X_10495_ _10495_/A _10495_/Y vdd gnd INVX1
XFILL_1__8818_ vdd gnd FILL
XFILL_2__8591_ vdd gnd FILL
X_12234_ _12234_/A _12234_/B _12234_/C _12234_/Y vdd gnd OAI21X1
XFILL_1__8749_ vdd gnd FILL
X_12165_ _12165_/A _12165_/B _12165_/C _12165_/Y vdd gnd NAND3X1
XFILL_1__11260_ vdd gnd FILL
X_11116_ _11116_/A _11116_/B _11116_/Y vdd gnd NAND2X1
XFILL_2__9212_ vdd gnd FILL
XFILL_0__11990_ vdd gnd FILL
X_12096_ _12096_/A _12096_/B _12096_/C _12096_/Y vdd gnd OAI21X1
XFILL_1__10211_ vdd gnd FILL
XFILL_1__11191_ vdd gnd FILL
XFILL_0__10941_ vdd gnd FILL
X_11047_ _11047_/A _11047_/Y vdd gnd INVX1
XFILL_2__9143_ vdd gnd FILL
XFILL_2__11501_ vdd gnd FILL
XFILL_1__10142_ vdd gnd FILL
XFILL_0__13660_ vdd gnd FILL
XFILL_0__10872_ vdd gnd FILL
XFILL_2__14220_ vdd gnd FILL
XFILL_2__9074_ vdd gnd FILL
XFILL_2__11432_ vdd gnd FILL
XFILL_1__10073_ vdd gnd FILL
XFILL_0__13591_ vdd gnd FILL
X_14806_ _14806_/A _14806_/B _14806_/Y vdd gnd NAND2X1
XFILL_1__13901_ vdd gnd FILL
XFILL_2__14151_ vdd gnd FILL
X_12998_ _12998_/A _12998_/B _12998_/Y vdd gnd NAND2X1
XFILL_2__11363_ vdd gnd FILL
X_14737_ _14737_/A _14737_/B _14737_/C _14737_/Y vdd gnd NAND3X1
X_11949_ _11949_/A _11949_/B _11949_/C _11949_/Y vdd gnd NAND3X1
XFILL_1__13832_ vdd gnd FILL
XFILL_2__14082_ vdd gnd FILL
XFILL_2__11294_ vdd gnd FILL
XFILL_0__12473_ vdd gnd FILL
X_14668_ _14668_/A _14668_/B _14668_/C _14668_/Y vdd gnd OAI21X1
XFILL_2__9976_ vdd gnd FILL
XFILL_0__11424_ vdd gnd FILL
XFILL_1__13763_ vdd gnd FILL
XFILL_1__10975_ vdd gnd FILL
X_13619_ _13619_/A _13619_/B _13619_/Y vdd gnd NAND2X1
XFILL_0__8991_ vdd gnd FILL
X_14599_ _14599_/A _14599_/B _14599_/Y vdd gnd NOR2X1
XFILL_1__12714_ vdd gnd FILL
XFILL_0__14143_ vdd gnd FILL
XFILL_0__11355_ vdd gnd FILL
XFILL_1__13694_ vdd gnd FILL
XFILL_0__10306_ vdd gnd FILL
XFILL_1__12645_ vdd gnd FILL
XFILL_0__11286_ vdd gnd FILL
XFILL_0__14074_ vdd gnd FILL
X_8220_ _8220_/A _8220_/B _8220_/C _8220_/Y vdd gnd OAI21X1
XFILL_0__7873_ vdd gnd FILL
XFILL_2__13935_ vdd gnd FILL
XFILL_0__10237_ vdd gnd FILL
XFILL_0__13025_ vdd gnd FILL
XFILL_2__8789_ vdd gnd FILL
XFILL_0__9612_ vdd gnd FILL
X_8151_ _8151_/A _8151_/B _8151_/C _8151_/Y vdd gnd AOI21X1
XFILL_1__14315_ vdd gnd FILL
XFILL_1__11527_ vdd gnd FILL
XFILL_2__13866_ vdd gnd FILL
XFILL_0__10168_ vdd gnd FILL
X_7102_ _7102_/A _7102_/B _7102_/C _7102_/Y vdd gnd OAI21X1
XFILL_0__9543_ vdd gnd FILL
X_8082_ _8082_/A _8082_/B _8082_/Y vdd gnd NAND2X1
XFILL_1__14246_ vdd gnd FILL
XFILL_2__12817_ vdd gnd FILL
XFILL_1__11458_ vdd gnd FILL
XFILL_0__10099_ vdd gnd FILL
XFILL_0__9474_ vdd gnd FILL
XFILL_1__10409_ vdd gnd FILL
XFILL_2__12748_ vdd gnd FILL
XFILL_0__13927_ vdd gnd FILL
XFILL_0__8425_ vdd gnd FILL
XFILL_1__11389_ vdd gnd FILL
XFILL_1__13128_ vdd gnd FILL
XFILL_2__12679_ vdd gnd FILL
XFILL_0__13858_ vdd gnd FILL
XFILL_0__8356_ vdd gnd FILL
X_8984_ _8984_/A _8984_/B _8984_/C _8984_/Y vdd gnd OAI21X1
XFILL_2__14418_ vdd gnd FILL
XFILL_0__12809_ vdd gnd FILL
XFILL_1__13059_ vdd gnd FILL
XFILL_0__7307_ vdd gnd FILL
XFILL_0__13789_ vdd gnd FILL
XFILL_1__7080_ vdd gnd FILL
X_7935_ _7935_/D _7935_/CLK _7935_/Q vdd gnd DFFPOSX1
XFILL_0__8287_ vdd gnd FILL
XFILL_2__14349_ vdd gnd FILL
XFILL_0__7238_ vdd gnd FILL
X_7866_ _7866_/A _7866_/B _7866_/Y vdd gnd NAND2X1
X_9605_ _9605_/A _9605_/Y vdd gnd INVX1
XFILL_0__7169_ vdd gnd FILL
X_7797_ _7797_/A _7797_/B _7797_/C _7797_/Y vdd gnd NAND3X1
X_9536_ _9536_/A _9536_/B _9536_/Y vdd gnd NOR2X1
XFILL_1__9721_ vdd gnd FILL
X_9467_ _9467_/A _9467_/B _9467_/C _9467_/Y vdd gnd OAI21X1
X_8418_ _8418_/A _8418_/B _8418_/Y vdd gnd NAND2X1
XFILL_1__9652_ vdd gnd FILL
X_9398_ _9398_/A _9398_/B _9398_/C _9398_/D _9398_/Y vdd gnd AOI22X1
X_10280_ _10280_/A _10280_/B _10280_/C _10280_/Y vdd gnd OAI21X1
XFILL_1__8603_ vdd gnd FILL
XFILL_1__9583_ vdd gnd FILL
X_8349_ _8349_/A _8349_/B _8349_/Y vdd gnd NAND2X1
XFILL_1__8534_ vdd gnd FILL
XFILL_1__8465_ vdd gnd FILL
XFILL_1__7416_ vdd gnd FILL
X_13970_ _13970_/A _13970_/B _13970_/Y vdd gnd NAND2X1
XFILL_1__8396_ vdd gnd FILL
X_12921_ _12921_/A _12921_/B _12921_/C _12921_/Y vdd gnd OAI21X1
XFILL_1__7347_ vdd gnd FILL
X_12852_ _12852_/A _12852_/B _12852_/Y vdd gnd NOR2X1
XFILL_1__7278_ vdd gnd FILL
XFILL_1__9017_ vdd gnd FILL
X_11803_ _11803_/A _11803_/B _11803_/Y vdd gnd NAND2X1
X_12783_ _12783_/A _12783_/B _12783_/C _12783_/Y vdd gnd NAND3X1
X_14522_ _14522_/D _14522_/CLK _14522_/Q vdd gnd DFFPOSX1
X_11734_ _11734_/A _11734_/Y vdd gnd INVX1
X_14453_ _14453_/A _14453_/B _14453_/Y vdd gnd NAND2X1
X_11665_ _11665_/D _11665_/CLK _11665_/Q vdd gnd DFFPOSX1
X_10616_ _10616_/A _10616_/B _10616_/C _10616_/Y vdd gnd OAI21X1
X_13404_ _13404_/A _13404_/B _13404_/Y vdd gnd NAND2X1
X_14384_ _14384_/A _14384_/B _14384_/C _14384_/Y vdd gnd NAND3X1
XFILL_1__9919_ vdd gnd FILL
X_11596_ _11596_/A _11596_/B _11596_/Y vdd gnd NAND2X1
XFILL_0__11140_ vdd gnd FILL
X_13335_ _13335_/A _13335_/Y vdd gnd INVX1
X_10547_ _10547_/A _10547_/B _10547_/Y vdd gnd NAND2X1
XFILL_1__12430_ vdd gnd FILL
XFILL_0__11071_ vdd gnd FILL
XFILL_2__11981_ vdd gnd FILL
X_13266_ _13266_/A _13266_/B _13266_/C _13266_/Y vdd gnd AOI21X1
X_10478_ _10478_/A _10478_/B _10478_/Y vdd gnd NAND2X1
XFILL_0__10022_ vdd gnd FILL
XFILL_2__8574_ vdd gnd FILL
XFILL_2__13720_ vdd gnd FILL
XFILL_1__12361_ vdd gnd FILL
X_12217_ _12217_/A _12217_/B _12217_/Y vdd gnd NAND2X1
X_13197_ _13197_/A _13197_/B _13197_/C _13197_/Y vdd gnd OAI21X1
XFILL_1__14100_ vdd gnd FILL
XFILL_1__11312_ vdd gnd FILL
XFILL_2__13651_ vdd gnd FILL
XFILL_0__14830_ vdd gnd FILL
XFILL_1__12292_ vdd gnd FILL
X_12148_ _12148_/A _12148_/B _12148_/C _12148_/D _12148_/Y vdd gnd AOI22X1
XFILL_1__14031_ vdd gnd FILL
XFILL_1__11243_ vdd gnd FILL
XFILL_2__13582_ vdd gnd FILL
XFILL_0__14761_ vdd gnd FILL
XFILL_0__11973_ vdd gnd FILL
X_12079_ _12079_/A _12079_/B _12079_/Y vdd gnd NAND2X1
XFILL_0__13712_ vdd gnd FILL
XFILL_0__10924_ vdd gnd FILL
XFILL_0__8210_ vdd gnd FILL
XFILL_1__11174_ vdd gnd FILL
XFILL_0__14692_ vdd gnd FILL
XFILL_0__9190_ vdd gnd FILL
XFILL_2__9126_ vdd gnd FILL
XFILL_1__10125_ vdd gnd FILL
XFILL_0__13643_ vdd gnd FILL
XFILL_0__8141_ vdd gnd FILL
XFILL_0__10855_ vdd gnd FILL
XFILL_2__9057_ vdd gnd FILL
XFILL_2__11415_ vdd gnd FILL
XFILL_1__10056_ vdd gnd FILL
XFILL_0__13574_ vdd gnd FILL
XFILL256650x75750 vdd gnd FILL
X_7720_ _7720_/A _7720_/B _7720_/C _7720_/D _7720_/Y vdd gnd OAI22X1
XFILL_0__8072_ vdd gnd FILL
XFILL_0__10786_ vdd gnd FILL
XFILL_2__11346_ vdd gnd FILL
XFILL_1__14864_ vdd gnd FILL
XFILL_0__12525_ vdd gnd FILL
X_7651_ _7651_/A _7651_/B _7651_/Y vdd gnd AND2X2
XFILL_1__13815_ vdd gnd FILL
XFILL_2__11277_ vdd gnd FILL
XFILL_1__14795_ vdd gnd FILL
XFILL_0__12456_ vdd gnd FILL
X_7582_ _7582_/A _7582_/B _7582_/Y vdd gnd NAND2X1
XFILL_2__9959_ vdd gnd FILL
XFILL_0__11407_ vdd gnd FILL
XFILL_1__13746_ vdd gnd FILL
XFILL_1__10958_ vdd gnd FILL
X_9321_ _9321_/A _9321_/B _9321_/C _9321_/Y vdd gnd NAND3X1
XFILL_0__12387_ vdd gnd FILL
XFILL_0__8974_ vdd gnd FILL
XFILL_0__14126_ vdd gnd FILL
XFILL_0__11338_ vdd gnd FILL
XFILL_1__13677_ vdd gnd FILL
XFILL_1__10889_ vdd gnd FILL
X_9252_ _9252_/A _9252_/B _9252_/Y vdd gnd AND2X2
XFILL_1__12628_ vdd gnd FILL
XFILL_0__14057_ vdd gnd FILL
X_8203_ _8203_/A _8203_/B _8203_/C _8203_/Y vdd gnd OAI21X1
XFILL_0__11269_ vdd gnd FILL
XFILL_0__7856_ vdd gnd FILL
X_9183_ _9183_/A _9183_/Y vdd gnd INVX1
XFILL_2__13918_ vdd gnd FILL
XFILL_0__13008_ vdd gnd FILL
X_8134_ _8134_/A _8134_/B _8134_/S _8134_/Y vdd gnd MUX2X1
XFILL_0__7787_ vdd gnd FILL
XFILL_2__13849_ vdd gnd FILL
XFILL_0__9526_ vdd gnd FILL
X_8065_ _8065_/A _8065_/Y vdd gnd INVX1
XFILL_1__14229_ vdd gnd FILL
XFILL_1__8250_ vdd gnd FILL
XFILL_0__9457_ vdd gnd FILL
XFILL_1__7201_ vdd gnd FILL
XFILL_0__8408_ vdd gnd FILL
XFILL_0__9388_ vdd gnd FILL
XFILL_1__8181_ vdd gnd FILL
XFILL_1__7132_ vdd gnd FILL
XFILL_0__8339_ vdd gnd FILL
X_8967_ _8967_/A _8967_/B _8967_/C _8967_/Y vdd gnd OAI21X1
X_7918_ _7918_/D _7918_/CLK _7918_/Q vdd gnd DFFPOSX1
X_8898_ _8898_/D _8898_/CLK _8898_/Q vdd gnd DFFPOSX1
XFILL_0_CLKBUF1_insert102 vdd gnd FILL
X_7849_ _7849_/A _7849_/B _7849_/Y vdd gnd NAND2X1
X_11450_ _11450_/A _11450_/B _11450_/Y vdd gnd OR2X2
X_9519_ _9519_/A _9519_/B _9519_/Y vdd gnd AND2X2
X_10401_ _10401_/A _10401_/B _10401_/Y vdd gnd NAND2X1
XFILL_1__9704_ vdd gnd FILL
X_11381_ _11381_/A _11381_/B _11381_/C _11381_/Y vdd gnd OAI21X1
X_13120_ _13120_/A _13120_/B _13120_/C _13120_/Y vdd gnd NAND3X1
XFILL_1__7896_ vdd gnd FILL
X_10332_ _10332_/A _10332_/B _10332_/Y vdd gnd NOR2X1
XFILL_1__9635_ vdd gnd FILL
X_13051_ _13051_/A _13051_/B _13051_/Y vdd gnd NAND2X1
X_10263_ _10263_/A _10263_/B _10263_/C _10263_/Y vdd gnd OAI21X1
XFILL_1__9566_ vdd gnd FILL
X_12002_ _12002_/A _12002_/B _12002_/C _12002_/Y vdd gnd NAND3X1
XFILL_2__7310_ vdd gnd FILL
X_10194_ _10194_/A _10194_/B _10194_/Y vdd gnd NAND2X1
XFILL_1__8517_ vdd gnd FILL
XFILL_1__9497_ vdd gnd FILL
XFILL_2__7241_ vdd gnd FILL
XFILL_1__8448_ vdd gnd FILL
X_13953_ _13953_/A _13953_/B _13953_/Y vdd gnd OR2X2
XFILL_2__7172_ vdd gnd FILL
XFILL_1__8379_ vdd gnd FILL
X_12904_ _12904_/A _12904_/Y vdd gnd INVX1
X_13884_ _13884_/A _13884_/B _13884_/Y vdd gnd NAND2X1
XFILL_0__10640_ vdd gnd FILL
X_12835_ _12835_/A _12835_/B _12835_/C _12835_/Y vdd gnd OAI21X1
XFILL_1__11930_ vdd gnd FILL
XFILL_0__10571_ vdd gnd FILL
X_12766_ _12766_/A _12766_/B _12766_/C _12766_/Y vdd gnd OAI21X1
XFILL_0__12310_ vdd gnd FILL
XFILL_1__11861_ vdd gnd FILL
X_14505_ _14505_/D _14505_/CLK _14505_/Q vdd gnd DFFPOSX1
XFILL_0__13290_ vdd gnd FILL
X_11717_ _11717_/A _11717_/B _11717_/C _11717_/Y vdd gnd OAI21X1
XFILL_1__13600_ vdd gnd FILL
X_12697_ _12697_/A _12697_/B _12697_/S _12697_/Y vdd gnd MUX2X1
XFILL_1__10812_ vdd gnd FILL
XFILL_1__14580_ vdd gnd FILL
XFILL_0__12241_ vdd gnd FILL
XFILL_1__11792_ vdd gnd FILL
X_14436_ _14436_/A _14436_/Y vdd gnd INVX1
X_11648_ _11648_/D _11648_/CLK _11648_/Q vdd gnd DFFPOSX1
XFILL_2__10013_ vdd gnd FILL
XFILL_1__13531_ vdd gnd FILL
XFILL_0__12172_ vdd gnd FILL
X_14367_ _14367_/A _14367_/B _14367_/C _14367_/Y vdd gnd OAI21X1
X_11579_ _11579_/A _11579_/B _11579_/C _11579_/Y vdd gnd OAI21X1
XFILL_0__11123_ vdd gnd FILL
XFILL_1__10674_ vdd gnd FILL
XFILL_0__7710_ vdd gnd FILL
X_13318_ _13318_/A _13318_/Y vdd gnd INVX1
XFILL_2_CLKBUF1_insert44 vdd gnd FILL
X_14298_ _14298_/A _14298_/B _14298_/Y vdd gnd NAND2X1
XFILL_0__8690_ vdd gnd FILL
XFILL_1__12413_ vdd gnd FILL
XFILL_2_CLKBUF1_insert55 vdd gnd FILL
XFILL_0__11054_ vdd gnd FILL
XFILL_1__13393_ vdd gnd FILL
XFILL_0__7641_ vdd gnd FILL
XFILL_2_CLKBUF1_insert77 vdd gnd FILL
X_13249_ _13249_/A _13249_/B _13249_/Y vdd gnd NAND2X1
XFILL_0__10005_ vdd gnd FILL
XFILL_2__10915_ vdd gnd FILL
XFILL_2__13703_ vdd gnd FILL
XFILL_1__12344_ vdd gnd FILL
XFILL_0__7572_ vdd gnd FILL
XFILL_2__7508_ vdd gnd FILL
XFILL_2__13634_ vdd gnd FILL
XFILL_0__14813_ vdd gnd FILL
XFILL_2__10846_ vdd gnd FILL
XFILL_1__12275_ vdd gnd FILL
XFILL_0__9311_ vdd gnd FILL
XFILL_1__14014_ vdd gnd FILL
XFILL_2__7439_ vdd gnd FILL
XFILL_2__13565_ vdd gnd FILL
XFILL_1__11226_ vdd gnd FILL
XFILL_0__14744_ vdd gnd FILL
XFILL_2__10777_ vdd gnd FILL
XFILL_0__9242_ vdd gnd FILL
XFILL_0_BUFX2_insert15 vdd gnd FILL
XFILL_0__11956_ vdd gnd FILL
XFILL_0_CLKBUF1_insert70 vdd gnd FILL
X_9870_ _9870_/A _9870_/B _9870_/C _9870_/Y vdd gnd AOI21X1
XFILL_0_BUFX2_insert26 vdd gnd FILL
XFILL_0_CLKBUF1_insert81 vdd gnd FILL
XFILL_0__10907_ vdd gnd FILL
XFILL_1__11157_ vdd gnd FILL
XFILL_0__14675_ vdd gnd FILL
XFILL_0_CLKBUF1_insert92 vdd gnd FILL
XFILL_0__9173_ vdd gnd FILL
XFILL_0__11887_ vdd gnd FILL
X_8821_ _8821_/A _8821_/Y vdd gnd INVX1
XFILL_1__10108_ vdd gnd FILL
XFILL_0__13626_ vdd gnd FILL
XFILL_1__11088_ vdd gnd FILL
XFILL_0__8124_ vdd gnd FILL
XFILL_0__10838_ vdd gnd FILL
X_8752_ _8752_/A _8752_/B _8752_/C _8752_/Y vdd gnd OAI21X1
XFILL_1__10039_ vdd gnd FILL
XFILL_1__14916_ vdd gnd FILL
XFILL_0__13557_ vdd gnd FILL
X_7703_ _7703_/A _7703_/B _7703_/Y vdd gnd NAND2X1
XFILL_0__8055_ vdd gnd FILL
XFILL_0__10769_ vdd gnd FILL
X_8683_ _8683_/A _8683_/B _8683_/Y vdd gnd NAND2X1
XFILL_2__11329_ vdd gnd FILL
XFILL_0__12508_ vdd gnd FILL
XFILL_1__14847_ vdd gnd FILL
X_7634_ _7634_/A _7634_/B _7634_/C _7634_/Y vdd gnd OAI21X1
XFILL_1__14778_ vdd gnd FILL
XFILL_0__12439_ vdd gnd FILL
X_7565_ _7565_/A _7565_/Y vdd gnd INVX1
XFILL_1__13729_ vdd gnd FILL
X_9304_ _9304_/A _9304_/B _9304_/C _9304_/Y vdd gnd OAI21X1
XFILL_1__7750_ vdd gnd FILL
XFILL_0__8957_ vdd gnd FILL
X_7496_ _7496_/A _7496_/Y vdd gnd INVX1
XFILL_0__14109_ vdd gnd FILL
X_9235_ _9235_/A _9235_/B _9235_/C _9235_/Y vdd gnd OAI21X1
XFILL_0__7908_ vdd gnd FILL
XFILL_1__7681_ vdd gnd FILL
XFILL_1__9420_ vdd gnd FILL
XFILL_0__7839_ vdd gnd FILL
X_9166_ _9166_/A _9166_/B _9166_/C _9166_/Y vdd gnd AOI21X1
X_8117_ _8117_/A _8117_/B _8117_/S _8117_/Y vdd gnd MUX2X1
XFILL_1__9351_ vdd gnd FILL
X_9097_ _9097_/A _9097_/B _9097_/C _9097_/Y vdd gnd OAI21X1
XFILL_0__9509_ vdd gnd FILL
XFILL_1__8302_ vdd gnd FILL
XFILL_1__9282_ vdd gnd FILL
X_8048_ _8048_/A _8048_/B _8048_/Y vdd gnd NOR2X1
XFILL_1__8233_ vdd gnd FILL
X_10950_ _10950_/A _10950_/B _10950_/C _10950_/Y vdd gnd AOI21X1
XFILL_1__8164_ vdd gnd FILL
X_9999_ _9999_/A _9999_/B _9999_/C _9999_/Y vdd gnd AOI21X1
XFILL_1__7115_ vdd gnd FILL
X_10881_ _10881_/A _10881_/B _10881_/S _10881_/Y vdd gnd MUX2X1
XFILL_1__8095_ vdd gnd FILL
X_12620_ _12620_/A _12620_/B _12620_/Y vdd gnd NOR2X1
X_12551_ _12551_/D _12551_/CLK _12551_/Q vdd gnd DFFPOSX1
X_11502_ _11502_/A _11502_/B _11502_/Y vdd gnd NOR2X1
X_12482_ _12482_/A _12482_/B _12482_/Y vdd gnd NAND2X1
XFILL_1__8997_ vdd gnd FILL
X_14221_ _14221_/A _14221_/B _14221_/C _14221_/Y vdd gnd OAI21X1
X_11433_ _11433_/A _11433_/Y vdd gnd INVX1
X_14152_ _14152_/A _14152_/B _14152_/C _14152_/Y vdd gnd OAI21X1
X_11364_ _11364_/A _11364_/B _11364_/Y vdd gnd NOR2X1
XFILL_2__9460_ vdd gnd FILL
XFILL_1__7879_ vdd gnd FILL
X_13103_ _13103_/A _13103_/B _13103_/C _13103_/Y vdd gnd NAND3X1
X_10315_ _10315_/A _10315_/B _10315_/Y vdd gnd OR2X2
X_14083_ _14083_/A _14083_/B _14083_/C _14083_/Y vdd gnd OAI21X1
XFILL_1__9618_ vdd gnd FILL
X_11295_ _11295_/A _11295_/Y vdd gnd INVX1
XFILL_2__9391_ vdd gnd FILL
X_13034_ _13034_/A _13034_/B _13034_/C _13034_/Y vdd gnd NAND3X1
XFILL_1__10390_ vdd gnd FILL
X_10246_ _10246_/A _10246_/B _10246_/S _10246_/Y vdd gnd MUX2X1
XFILL_1__9549_ vdd gnd FILL
X_10177_ _10177_/A _10177_/B _10177_/Y vdd gnd NAND2X1
XFILL_1__12060_ vdd gnd FILL
XFILL_0__11810_ vdd gnd FILL
XFILL_0__12790_ vdd gnd FILL
XFILL_2__7224_ vdd gnd FILL
XFILL_1__11011_ vdd gnd FILL
XFILL_0__11741_ vdd gnd FILL
X_13936_ _13936_/A _13936_/Y vdd gnd INVX1
XFILL_2__12301_ vdd gnd FILL
XFILL_2__7155_ vdd gnd FILL
XFILL_0__14460_ vdd gnd FILL
X_13867_ _13867_/A _13867_/B _13867_/Y vdd gnd NAND2X1
XFILL_2__12232_ vdd gnd FILL
XFILL_2__7086_ vdd gnd FILL
XFILL_0__13411_ vdd gnd FILL
XFILL_1__12962_ vdd gnd FILL
XFILL_0__10623_ vdd gnd FILL
XFILL_0__14391_ vdd gnd FILL
XFILL_1_BUFX2_insert340 vdd gnd FILL
X_12818_ _12818_/A _12818_/B _12818_/C _12818_/Y vdd gnd NAND3X1
XFILL_1_BUFX2_insert351 vdd gnd FILL
XFILL_1__14701_ vdd gnd FILL
XFILL_1_BUFX2_insert362 vdd gnd FILL
XFILL_1__11913_ vdd gnd FILL
XFILL_2__12163_ vdd gnd FILL
X_13798_ _13798_/A _13798_/B _13798_/C _13798_/Y vdd gnd OAI21X1
XFILL_1_BUFX2_insert373 vdd gnd FILL
XFILL_0__13342_ vdd gnd FILL
XFILL_0__10554_ vdd gnd FILL
XFILL_1__12893_ vdd gnd FILL
X_12749_ _12749_/A _12749_/B _12749_/Y vdd gnd NAND2X1
XFILL_1__14632_ vdd gnd FILL
XFILL_1__11844_ vdd gnd FILL
XFILL_0__13273_ vdd gnd FILL
XFILL_0__10485_ vdd gnd FILL
XFILL_0__9860_ vdd gnd FILL
XFILL_1__14563_ vdd gnd FILL
XFILL_0__12224_ vdd gnd FILL
XFILL_1__11775_ vdd gnd FILL
X_14419_ _14419_/A _14419_/B _14419_/C _14419_/Y vdd gnd OAI21X1
XFILL_0__8811_ vdd gnd FILL
X_7350_ _7350_/A _7350_/B _7350_/C _7350_/Y vdd gnd OAI21X1
XFILL_2__9727_ vdd gnd FILL
XFILL_1__13514_ vdd gnd FILL
XFILL_1__14494_ vdd gnd FILL
XFILL_0__12155_ vdd gnd FILL
XFILL_0__8742_ vdd gnd FILL
X_7281_ _7281_/A _7281_/B _7281_/C _7281_/Y vdd gnd NAND3X1
XFILL_0__11106_ vdd gnd FILL
XFILL_2__9658_ vdd gnd FILL
XFILL_1__10657_ vdd gnd FILL
X_9020_ _9020_/A _9020_/Y vdd gnd INVX1
XFILL_0__12086_ vdd gnd FILL
XFILL_2__12996_ vdd gnd FILL
XFILL_0__8673_ vdd gnd FILL
XFILL_0__11037_ vdd gnd FILL
XFILL_2__9589_ vdd gnd FILL
XFILL_1__13376_ vdd gnd FILL
XFILL_1__10588_ vdd gnd FILL
XFILL_0__7624_ vdd gnd FILL
XFILL_1__12327_ vdd gnd FILL
XFILL_0__7555_ vdd gnd FILL
XFILL_2__10829_ vdd gnd FILL
XFILL_1__12258_ vdd gnd FILL
XFILL_0__12988_ vdd gnd FILL
XFILL_0__7486_ vdd gnd FILL
X_9922_ _9922_/A _9922_/B _9922_/Y vdd gnd NAND2X1
XFILL_1__11209_ vdd gnd FILL
XFILL_0__14727_ vdd gnd FILL
XFILL_0__11939_ vdd gnd FILL
XFILL_1__12189_ vdd gnd FILL
XFILL_0__9225_ vdd gnd FILL
X_9853_ _9853_/A _9853_/B _9853_/Y vdd gnd AND2X2
XFILL_0__14658_ vdd gnd FILL
XFILL_0__9156_ vdd gnd FILL
X_8804_ _8804_/A _8804_/B _8804_/Y vdd gnd NAND2X1
X_9784_ _9784_/D _9784_/CLK _9784_/Q vdd gnd DFFPOSX1
XFILL_0__13609_ vdd gnd FILL
XFILL_0__8107_ vdd gnd FILL
XFILL_0__14589_ vdd gnd FILL
XFILL_0__9087_ vdd gnd FILL
X_8735_ _8735_/A _8735_/B _8735_/Y vdd gnd OR2X2
XFILL_0__8038_ vdd gnd FILL
XFILL_1__8920_ vdd gnd FILL
X_8666_ _8666_/A _8666_/B _8666_/Y vdd gnd NAND2X1
X_7617_ _7617_/A _7617_/B _7617_/C _7617_/Y vdd gnd AOI21X1
X_8597_ _8597_/A _8597_/B _8597_/Y vdd gnd NOR2X1
XFILL_1__7802_ vdd gnd FILL
X_7548_ _7548_/A _7548_/B _7548_/Y vdd gnd NAND2X1
XFILL_0__9989_ vdd gnd FILL
XFILL_1__8782_ vdd gnd FILL
XFILL_1__7733_ vdd gnd FILL
X_7479_ _7479_/A _7479_/B _7479_/C _7479_/Y vdd gnd NAND3X1
X_9218_ _9218_/A _9218_/B _9218_/C _9218_/D _9218_/Y vdd gnd AOI22X1
XFILL_1__7664_ vdd gnd FILL
X_10100_ _10100_/A _10100_/Y vdd gnd INVX1
X_11080_ _11080_/A _11080_/B _11080_/C _11080_/Y vdd gnd OAI21X1
XFILL_1__9403_ vdd gnd FILL
X_9149_ _9149_/A _9149_/B _9149_/C _9149_/Y vdd gnd NAND3X1
XFILL_1__7595_ vdd gnd FILL
X_10031_ _10031_/A _10031_/Y vdd gnd INVX1
XFILL257550x10950 vdd gnd FILL
XFILL_1__9334_ vdd gnd FILL
XFILL_1__9265_ vdd gnd FILL
X_14770_ _14770_/A _14770_/B _14770_/Y vdd gnd NAND2X1
XFILL_1__8216_ vdd gnd FILL
XFILL_1__9196_ vdd gnd FILL
X_11982_ _11982_/A _11982_/B _11982_/C _11982_/Y vdd gnd NAND3X1
X_13721_ _13721_/A _13721_/B _13721_/C _13721_/Y vdd gnd OAI21X1
XFILL_1__8147_ vdd gnd FILL
X_10933_ _10933_/A _10933_/Y vdd gnd INVX1
XFILL_0_BUFX2_insert7 vdd gnd FILL
X_13652_ _13652_/A _13652_/B _13652_/Y vdd gnd NAND2X1
X_10864_ _10864_/A _10864_/B _10864_/C _10864_/Y vdd gnd NAND3X1
XFILL_1__8078_ vdd gnd FILL
X_12603_ _12603_/D _12603_/CLK _12603_/Q vdd gnd DFFPOSX1
XFILL_2__7911_ vdd gnd FILL
XFILL_0_BUFX2_insert303 vdd gnd FILL
X_10795_ _10795_/A _10795_/Y vdd gnd INVX1
X_13583_ _13583_/A _13583_/B _13583_/C _13583_/D _13583_/Y vdd gnd OAI22X1
XFILL_0_BUFX2_insert314 vdd gnd FILL
XFILL_0_BUFX2_insert325 vdd gnd FILL
XFILL_0_BUFX2_insert336 vdd gnd FILL
X_12534_ _12534_/A _12534_/B _12534_/Y vdd gnd NAND2X1
XFILL_0_BUFX2_insert347 vdd gnd FILL
XFILL_0_BUFX2_insert358 vdd gnd FILL
XFILL_0_BUFX2_insert369 vdd gnd FILL
XFILL_0__10270_ vdd gnd FILL
X_12465_ _12465_/A _12465_/B _12465_/C _12465_/Y vdd gnd OAI21X1
XFILL_1__11560_ vdd gnd FILL
X_14204_ _14204_/D _14204_/CLK _14204_/Q vdd gnd DFFPOSX1
X_11416_ _11416_/A _11416_/B _11416_/C _11416_/D _11416_/Y vdd gnd OAI22X1
XFILL_2__9512_ vdd gnd FILL
X_12396_ _12396_/A _12396_/Y vdd gnd INVX1
XFILL_1__10511_ vdd gnd FILL
XFILL_2__12850_ vdd gnd FILL
XFILL_1__11491_ vdd gnd FILL
X_11347_ _11347_/A _11347_/B _11347_/Y vdd gnd AND2X2
X_14135_ _14135_/A _14135_/Y vdd gnd INVX1
XFILL_2__9443_ vdd gnd FILL
XFILL_1__13230_ vdd gnd FILL
XFILL_1__10442_ vdd gnd FILL
XFILL_2__12781_ vdd gnd FILL
XFILL_0__13960_ vdd gnd FILL
X_14066_ _14066_/A _14066_/B _14066_/C _14066_/Y vdd gnd OAI21X1
X_11278_ _11278_/A _11278_/B _11278_/Y vdd gnd NAND2X1
XFILL_1__13161_ vdd gnd FILL
XFILL_2__9374_ vdd gnd FILL
XFILL_0__12911_ vdd gnd FILL
XFILL_1__10373_ vdd gnd FILL
XFILL_0__13891_ vdd gnd FILL
X_10229_ _10229_/A _10229_/B _10229_/Y vdd gnd NAND2X1
X_13017_ _13017_/A _13017_/B _13017_/Y vdd gnd AND2X2
XFILL_1__12112_ vdd gnd FILL
XFILL_0__12842_ vdd gnd FILL
XFILL_1__13092_ vdd gnd FILL
XFILL_0__7340_ vdd gnd FILL
XFILL_2__14382_ vdd gnd FILL
XFILL_1__12043_ vdd gnd FILL
XFILL_2__11594_ vdd gnd FILL
XFILL_0__12773_ vdd gnd FILL
XFILL_0__7271_ vdd gnd FILL
XFILL_0__9010_ vdd gnd FILL
XFILL_0__11724_ vdd gnd FILL
X_13919_ _13919_/A _13919_/B _13919_/Y vdd gnd NOR2X1
XFILL_2__7138_ vdd gnd FILL
X_14899_ _14899_/D _14899_/CLK _14899_/Q vdd gnd DFFPOSX1
XFILL_0__14443_ vdd gnd FILL
XFILL_1__13994_ vdd gnd FILL
XFILL_2__12215_ vdd gnd FILL
XFILL_0__10606_ vdd gnd FILL
XFILL_1__12945_ vdd gnd FILL
XFILL_0__14374_ vdd gnd FILL
XFILL_1_BUFX2_insert170 vdd gnd FILL
X_8520_ _8520_/A _8520_/B _8520_/C _8520_/Y vdd gnd OAI21X1
XFILL_0__11586_ vdd gnd FILL
XFILL_1_BUFX2_insert181 vdd gnd FILL
XFILL_2__12146_ vdd gnd FILL
XFILL_1_BUFX2_insert192 vdd gnd FILL
XFILL_0__13325_ vdd gnd FILL
XFILL_0__10537_ vdd gnd FILL
XFILL_1__12876_ vdd gnd FILL
XFILL_0__9912_ vdd gnd FILL
X_8451_ _8451_/A _8451_/B _8451_/Y vdd gnd NAND2X1
XFILL_1__14615_ vdd gnd FILL
XFILL_1__11827_ vdd gnd FILL
XFILL_2__12077_ vdd gnd FILL
XFILL_0__13256_ vdd gnd FILL
XFILL256950x248550 vdd gnd FILL
X_7402_ _7402_/A _7402_/B _7402_/Y vdd gnd NAND2X1
XFILL_0__10468_ vdd gnd FILL
X_8382_ _8382_/A _8382_/B _8382_/Y vdd gnd NOR2X1
XFILL_0__12207_ vdd gnd FILL
XFILL_1__11758_ vdd gnd FILL
XFILL_0__13187_ vdd gnd FILL
XFILL_0__10399_ vdd gnd FILL
X_7333_ _7333_/A _7333_/B _7333_/C _7333_/Y vdd gnd OAI21X1
XFILL_1__14477_ vdd gnd FILL
XFILL_0__12138_ vdd gnd FILL
XFILL_0__8725_ vdd gnd FILL
X_7264_ _7264_/A _7264_/B _7264_/Y vdd gnd NAND2X1
X_9003_ _9003_/A _9003_/B _9003_/C _9003_/Y vdd gnd OAI21X1
XFILL_0__12069_ vdd gnd FILL
XFILL_2__12979_ vdd gnd FILL
XFILL_0__8656_ vdd gnd FILL
X_7195_ _7195_/A _7195_/B _7195_/C _7195_/Y vdd gnd OAI21X1
XFILL_1__13359_ vdd gnd FILL
XFILL_0__7607_ vdd gnd FILL
XFILL_1__7380_ vdd gnd FILL
XFILL_0__8587_ vdd gnd FILL
XFILL_0__7538_ vdd gnd FILL
XFILL_1__9050_ vdd gnd FILL
X_9905_ _9905_/A _9905_/Y vdd gnd INVX8
XFILL_0__7469_ vdd gnd FILL
XFILL_1__8001_ vdd gnd FILL
XFILL_0__9208_ vdd gnd FILL
X_9836_ _9836_/D _9836_/CLK _9836_/Q vdd gnd DFFPOSX1
XFILL_0__9139_ vdd gnd FILL
X_9767_ _9767_/D _9767_/CLK _9767_/Q vdd gnd DFFPOSX1
XFILL_1__9952_ vdd gnd FILL
X_8718_ _8718_/A _8718_/B _8718_/Y vdd gnd NAND2X1
X_9698_ _9698_/A _9698_/B _9698_/C _9698_/Y vdd gnd OAI21X1
X_10580_ _10580_/A _10580_/B _10580_/Y vdd gnd NAND2X1
X_8649_ _8649_/A _8649_/B _8649_/Y vdd gnd NOR2X1
XFILL_1__9883_ vdd gnd FILL
XFILL_1__8834_ vdd gnd FILL
X_12250_ _12250_/A _12250_/B _12250_/C _12250_/Y vdd gnd AOI21X1
XFILL_1__8765_ vdd gnd FILL
X_11201_ _11201_/A _11201_/B _11201_/Y vdd gnd NOR2X1
X_12181_ _12181_/A _12181_/B _12181_/C _12181_/Y vdd gnd NAND3X1
XFILL_1__7716_ vdd gnd FILL
XFILL_1__8696_ vdd gnd FILL
X_11132_ _11132_/A _11132_/B _11132_/Y vdd gnd NAND2X1
XFILL_1__7647_ vdd gnd FILL
X_11063_ _11063_/A _11063_/Y vdd gnd INVX1
XFILL_1__7578_ vdd gnd FILL
X_10014_ _10014_/A _10014_/B _10014_/Y vdd gnd NOR2X1
XFILL_1__9317_ vdd gnd FILL
XFILL_2__8110_ vdd gnd FILL
XFILL257250x57750 vdd gnd FILL
X_14822_ _14822_/A _14822_/B _14822_/Y vdd gnd NOR2X1
XFILL_2__8041_ vdd gnd FILL
XFILL_1__9248_ vdd gnd FILL
X_14753_ _14753_/A _14753_/B _14753_/Y vdd gnd NAND2X1
XFILL_2__10330_ vdd gnd FILL
X_11965_ _11965_/A _11965_/B _11965_/C _11965_/Y vdd gnd OAI21X1
XFILL_1__9179_ vdd gnd FILL
X_13704_ _13704_/A _13704_/B _13704_/C _13704_/Y vdd gnd OAI21X1
X_10916_ _10916_/A _10916_/B _10916_/C _10916_/Y vdd gnd AOI21X1
X_14684_ _14684_/A _14684_/B _14684_/C _14684_/Y vdd gnd NAND3X1
X_11896_ _11896_/A _11896_/B _11896_/C _11896_/Y vdd gnd AOI21X1
XFILL_0__11440_ vdd gnd FILL
XFILL_1__10991_ vdd gnd FILL
X_13635_ _13635_/A _13635_/B _13635_/C _13635_/Y vdd gnd NAND3X1
XFILL_2__12000_ vdd gnd FILL
X_10847_ _10847_/A _10847_/Y vdd gnd INVX1
XFILL_2__8943_ vdd gnd FILL
XFILL_1__12730_ vdd gnd FILL
XFILL_0_BUFX2_insert111 vdd gnd FILL
XFILL_0__11371_ vdd gnd FILL
XFILL_0_BUFX2_insert122 vdd gnd FILL
XFILL_0_BUFX2_insert133 vdd gnd FILL
X_13566_ _13566_/A _13566_/B _13566_/Y vdd gnd NAND2X1
XFILL_0__13110_ vdd gnd FILL
XFILL_0_BUFX2_insert144 vdd gnd FILL
X_10778_ _10778_/A _10778_/B _10778_/C _10778_/D _10778_/Y vdd gnd AOI22X1
XFILL_1__12661_ vdd gnd FILL
XFILL_0__10322_ vdd gnd FILL
XFILL_0__14090_ vdd gnd FILL
XFILL_0_BUFX2_insert155 vdd gnd FILL
X_12517_ _12517_/A _12517_/Y vdd gnd INVX1
XFILL_0_BUFX2_insert166 vdd gnd FILL
XFILL_0_BUFX2_insert177 vdd gnd FILL
XFILL_0_BUFX2_insert188 vdd gnd FILL
XFILL_2__7825_ vdd gnd FILL
XFILL_1__14400_ vdd gnd FILL
X_13497_ _13497_/D _13497_/CLK _13497_/Q vdd gnd DFFPOSX1
XFILL_2__13951_ vdd gnd FILL
XFILL_0__13041_ vdd gnd FILL
XFILL_0_BUFX2_insert199 vdd gnd FILL
XFILL_0__10253_ vdd gnd FILL
X_12448_ _12448_/A _12448_/B _12448_/C _12448_/Y vdd gnd OAI21X1
XFILL_1__14331_ vdd gnd FILL
XFILL_2__7756_ vdd gnd FILL
XFILL_1__11543_ vdd gnd FILL
XFILL_2__13882_ vdd gnd FILL
XFILL_0__10184_ vdd gnd FILL
X_12379_ _12379_/A _12379_/B _12379_/Y vdd gnd NAND2X1
XFILL_1__14262_ vdd gnd FILL
XFILL_1_CLKBUF1_insert391 vdd gnd FILL
XFILL_2__7687_ vdd gnd FILL
XFILL_1__11474_ vdd gnd FILL
XFILL_0__8510_ vdd gnd FILL
X_14118_ _14118_/A _14118_/B _14118_/Y vdd gnd AND2X2
XFILL_1__13213_ vdd gnd FILL
XFILL_0__9490_ vdd gnd FILL
XFILL_1__10425_ vdd gnd FILL
XFILL_0__13943_ vdd gnd FILL
XFILL_2__12764_ vdd gnd FILL
XFILL_0__8441_ vdd gnd FILL
X_14049_ _14049_/A _14049_/Y vdd gnd INVX1
XFILL_1__13144_ vdd gnd FILL
XFILL_2__9357_ vdd gnd FILL
XFILL_1__10356_ vdd gnd FILL
XFILL_0__13874_ vdd gnd FILL
XFILL_2__12695_ vdd gnd FILL
XFILL_0__8372_ vdd gnd FILL
XFILL_2__8308_ vdd gnd FILL
XFILL_1__13075_ vdd gnd FILL
XFILL_2__9288_ vdd gnd FILL
XFILL_0__12825_ vdd gnd FILL
XFILL256950x223350 vdd gnd FILL
XFILL_1__10287_ vdd gnd FILL
XFILL257550x208950 vdd gnd FILL
XFILL_0__7323_ vdd gnd FILL
X_7951_ _7951_/D _7951_/CLK _7951_/Q vdd gnd DFFPOSX1
XFILL_1__12026_ vdd gnd FILL
XFILL_2__11577_ vdd gnd FILL
XFILL_0__12756_ vdd gnd FILL
XFILL_0__7254_ vdd gnd FILL
X_7882_ _7882_/A _7882_/B _7882_/C _7882_/Y vdd gnd OAI21X1
XFILL_0__11707_ vdd gnd FILL
XFILL_0__12687_ vdd gnd FILL
XFILL_0__7185_ vdd gnd FILL
X_9621_ _9621_/A _9621_/B _9621_/Y vdd gnd NAND2X1
XFILL_0__14426_ vdd gnd FILL
XFILL_1__13977_ vdd gnd FILL
X_9552_ _9552_/A _9552_/B _9552_/Y vdd gnd NOR2X1
XFILL_1__12928_ vdd gnd FILL
XFILL_0__14357_ vdd gnd FILL
X_8503_ _8503_/A _8503_/Y vdd gnd INVX1
XFILL_0__11569_ vdd gnd FILL
X_9483_ _9483_/A _9483_/Y vdd gnd INVX1
XFILL_2__12129_ vdd gnd FILL
XFILL_0__13308_ vdd gnd FILL
XBUFX2_insert17 BUFX2_insert17/A BUFX2_insert17/Y vdd gnd BUFX2
XFILL_0__14288_ vdd gnd FILL
XFILL_1__12859_ vdd gnd FILL
X_8434_ _8434_/A _8434_/B _8434_/Y vdd gnd NAND2X1
XBUFX2_insert28 BUFX2_insert28/A BUFX2_insert28/Y vdd gnd BUFX2
XFILL_0__13239_ vdd gnd FILL
X_8365_ _8365_/A _8365_/B _8365_/C _8365_/D _8365_/Y vdd gnd AOI22X1
X_7316_ _7316_/A _7316_/B _7316_/C _7316_/Y vdd gnd OAI21X1
XFILL_0__9757_ vdd gnd FILL
XFILL_1__8550_ vdd gnd FILL
X_8296_ _8296_/A _8296_/B _8296_/Y vdd gnd AND2X2
XFILL_1__7501_ vdd gnd FILL
XFILL_0__8708_ vdd gnd FILL
X_7247_ _7247_/A _7247_/Y vdd gnd INVX1
XFILL_0__9688_ vdd gnd FILL
XFILL_1__8481_ vdd gnd FILL
XFILL_1__7432_ vdd gnd FILL
XFILL_0__8639_ vdd gnd FILL
X_7178_ _7178_/A _7178_/B _7178_/S _7178_/Y vdd gnd MUX2X1
XCLKBUF1_insert390 CLKBUF1_insert390/A CLKBUF1_insert390/Y vdd gnd CLKBUF1
XFILL_1__7363_ vdd gnd FILL
XFILL257250x150 vdd gnd FILL
XFILL_2_BUFX2_insert206 vdd gnd FILL
XFILL_1__9102_ vdd gnd FILL
XFILL257550x118950 vdd gnd FILL
XFILL_2_BUFX2_insert239 vdd gnd FILL
XFILL_1__7294_ vdd gnd FILL
XFILL_1__9033_ vdd gnd FILL
X_11750_ _11750_/A _11750_/Y vdd gnd INVX1
X_9819_ _9819_/D _9819_/CLK _9819_/Q vdd gnd DFFPOSX1
X_10701_ _10701_/D _10701_/CLK _10701_/Q vdd gnd DFFPOSX1
X_11681_ _11681_/D _11681_/CLK _11681_/Q vdd gnd DFFPOSX1
XBUFX2_insert205 BUFX2_insert205/A BUFX2_insert205/Y vdd gnd BUFX2
XBUFX2_insert216 BUFX2_insert216/A BUFX2_insert216/Y vdd gnd BUFX2
X_13420_ _13420_/A _13420_/B _13420_/C _13420_/Y vdd gnd OAI21X1
XBUFX2_insert227 BUFX2_insert227/A BUFX2_insert227/Y vdd gnd BUFX2
X_10632_ _10632_/A _10632_/B _10632_/Y vdd gnd NAND2X1
XBUFX2_insert238 BUFX2_insert238/A BUFX2_insert238/Y vdd gnd BUFX2
XFILL_1__9935_ vdd gnd FILL
XBUFX2_insert249 BUFX2_insert249/A BUFX2_insert249/Y vdd gnd BUFX2
X_10563_ _10563_/A _10563_/B _10563_/Y vdd gnd OR2X2
X_13351_ _13351_/A _13351_/Y vdd gnd INVX1
XFILL_1__9866_ vdd gnd FILL
X_12302_ _12302_/A _12302_/B _12302_/Y vdd gnd AND2X2
XFILL_2__7610_ vdd gnd FILL
X_10494_ _10494_/A _10494_/B _10494_/Y vdd gnd NAND2X1
XFILL_1__8817_ vdd gnd FILL
X_13282_ _13282_/A _13282_/Y vdd gnd INVX1
X_12233_ _12233_/A _12233_/B _12233_/Y vdd gnd NAND2X1
XFILL_2__7541_ vdd gnd FILL
XFILL_1__8748_ vdd gnd FILL
X_12164_ _12164_/A _12164_/B _12164_/C _12164_/Y vdd gnd OAI21X1
XFILL_2__7472_ vdd gnd FILL
XFILL_1__8679_ vdd gnd FILL
X_11115_ _11115_/A _11115_/Y vdd gnd INVX1
X_12095_ _12095_/A _12095_/B _12095_/S _12095_/Y vdd gnd MUX2X1
XFILL_1__10210_ vdd gnd FILL
XFILL_0__10940_ vdd gnd FILL
XFILL_1__11190_ vdd gnd FILL
X_11046_ _11046_/A _11046_/B _11046_/C _11046_/Y vdd gnd OAI21X1
XFILL_1__10141_ vdd gnd FILL
XFILL_0__10871_ vdd gnd FILL
XFILL_1__10072_ vdd gnd FILL
X_14805_ _14805_/A _14805_/B _14805_/C _14805_/Y vdd gnd OAI21X1
XFILL_0__13590_ vdd gnd FILL
XFILL_2__8024_ vdd gnd FILL
XFILL_1__13900_ vdd gnd FILL
X_12997_ _12997_/A _12997_/B _12997_/C _12997_/Y vdd gnd OAI21X1
X_14736_ _14736_/A _14736_/B _14736_/C _14736_/Y vdd gnd NAND3X1
XFILL_2__10313_ vdd gnd FILL
X_11948_ _11948_/A _11948_/Y vdd gnd INVX1
XFILL_1__13831_ vdd gnd FILL
XFILL_0__12472_ vdd gnd FILL
X_14667_ _14667_/A _14667_/Y vdd gnd INVX1
XFILL_2__10244_ vdd gnd FILL
X_11879_ _11879_/A _11879_/Y vdd gnd INVX1
XFILL_0__11423_ vdd gnd FILL
XFILL_1__13762_ vdd gnd FILL
XFILL_1__10974_ vdd gnd FILL
X_13618_ _13618_/A _13618_/Y vdd gnd INVX1
XFILL_0__8990_ vdd gnd FILL
X_14598_ _14598_/A _14598_/B _14598_/Y vdd gnd NOR2X1
XFILL_2__8926_ vdd gnd FILL
XFILL_2__10175_ vdd gnd FILL
XFILL_1__12713_ vdd gnd FILL
XFILL_0__14142_ vdd gnd FILL
XFILL_0__11354_ vdd gnd FILL
XFILL_1__13693_ vdd gnd FILL
X_13549_ _13549_/A _13549_/B _13549_/Y vdd gnd NAND2X1
XFILL_1__12644_ vdd gnd FILL
XFILL_0__10305_ vdd gnd FILL
XFILL_0__14073_ vdd gnd FILL
XFILL_0__11285_ vdd gnd FILL
XFILL_0__7872_ vdd gnd FILL
XFILL_2__7808_ vdd gnd FILL
XFILL_0__13024_ vdd gnd FILL
XFILL_0__10236_ vdd gnd FILL
XFILL_0__9611_ vdd gnd FILL
X_8150_ _8150_/A _8150_/B _8150_/C _8150_/Y vdd gnd OAI21X1
XFILL_2__7739_ vdd gnd FILL
XFILL_1__14314_ vdd gnd FILL
XFILL_1__11526_ vdd gnd FILL
X_7101_ _7101_/A _7101_/B _7101_/C _7101_/Y vdd gnd OAI21X1
XFILL_0__10167_ vdd gnd FILL
XFILL_0__9542_ vdd gnd FILL
X_8081_ _8081_/A _8081_/Y vdd gnd INVX8
XFILL_1__14245_ vdd gnd FILL
XFILL_1__11457_ vdd gnd FILL
XFILL_2__13796_ vdd gnd FILL
XFILL_0__10098_ vdd gnd FILL
XFILL_0__9473_ vdd gnd FILL
XFILL_1__10408_ vdd gnd FILL
XFILL_1__11388_ vdd gnd FILL
XFILL_0__13926_ vdd gnd FILL
XFILL_0__8424_ vdd gnd FILL
XFILL_1__13127_ vdd gnd FILL
XFILL_1__10339_ vdd gnd FILL
XFILL_0__13857_ vdd gnd FILL
XFILL_0__8355_ vdd gnd FILL
X_8983_ _8983_/A _8983_/B _8983_/Y vdd gnd NAND2X1
XFILL_1__13058_ vdd gnd FILL
XFILL_0__12808_ vdd gnd FILL
XFILL_0__7306_ vdd gnd FILL
XFILL_0__13788_ vdd gnd FILL
X_7934_ _7934_/D _7934_/CLK _7934_/Q vdd gnd DFFPOSX1
XFILL_1__12009_ vdd gnd FILL
XFILL_0__8286_ vdd gnd FILL
XFILL_0__12739_ vdd gnd FILL
XFILL_0__7237_ vdd gnd FILL
X_7865_ _7865_/A _7865_/B _7865_/C _7865_/Y vdd gnd OAI21X1
XFILL_0__7168_ vdd gnd FILL
X_9604_ _9604_/A _9604_/B _9604_/Y vdd gnd NAND2X1
X_7796_ _7796_/A _7796_/Y vdd gnd INVX1
XFILL_0__14409_ vdd gnd FILL
XFILL_0__7099_ vdd gnd FILL
X_9535_ _9535_/A _9535_/Y vdd gnd INVX1
XFILL_1__9720_ vdd gnd FILL
X_9466_ _9466_/A _9466_/B _9466_/C _9466_/D _9466_/Y vdd gnd AOI22X1
XFILL_1__9651_ vdd gnd FILL
X_8417_ _8417_/A _8417_/B _8417_/Y vdd gnd NAND2X1
X_9397_ _9397_/A _9397_/B _9397_/Y vdd gnd NAND2X1
XFILL_1__8602_ vdd gnd FILL
X_8348_ _8348_/A _8348_/Y vdd gnd INVX1
XFILL_1__9582_ vdd gnd FILL
XFILL_1__8533_ vdd gnd FILL
X_8279_ _8279_/A _8279_/Y vdd gnd INVX1
XFILL_1__8464_ vdd gnd FILL
XFILL_1__7415_ vdd gnd FILL
XFILL_1__8395_ vdd gnd FILL
X_12920_ _12920_/A _12920_/Y vdd gnd INVX1
XFILL_1__7346_ vdd gnd FILL
X_12851_ _12851_/A _12851_/B _12851_/C _12851_/Y vdd gnd AOI21X1
XFILL_1__7277_ vdd gnd FILL
X_11802_ _11802_/A _11802_/Y vdd gnd INVX1
XFILL_1__9016_ vdd gnd FILL
X_12782_ _12782_/A _12782_/B _12782_/C _12782_/Y vdd gnd OAI21X1
X_14521_ _14521_/D _14521_/CLK _14521_/Q vdd gnd DFFPOSX1
X_11733_ _11733_/A _11733_/B _11733_/Y vdd gnd NAND2X1
X_14452_ _14452_/A _14452_/B _14452_/Y vdd gnd NAND2X1
X_11664_ _11664_/D _11664_/CLK _11664_/Q vdd gnd DFFPOSX1
XFILL_2__9760_ vdd gnd FILL
X_13403_ _13403_/A _13403_/B _13403_/C _13403_/Y vdd gnd OAI21X1
X_10615_ _10615_/A _10615_/Y vdd gnd INVX1
XFILL_1__9918_ vdd gnd FILL
X_14383_ _14383_/A _14383_/B _14383_/Y vdd gnd NAND2X1
X_11595_ _11595_/A _11595_/B _11595_/C _11595_/Y vdd gnd OAI21X1
XFILL_2__9691_ vdd gnd FILL
X_13334_ _13334_/A _13334_/B _13334_/C _13334_/Y vdd gnd NAND3X1
X_10546_ _10546_/A _10546_/B _10546_/Y vdd gnd OR2X2
XFILL_1__9849_ vdd gnd FILL
XFILL_0__11070_ vdd gnd FILL
X_13265_ _13265_/A _13265_/Y vdd gnd INVX1
X_10477_ _10477_/A _10477_/B _10477_/Y vdd gnd NAND2X1
XFILL_0__10021_ vdd gnd FILL
XFILL_1__12360_ vdd gnd FILL
XFILL_2__10931_ vdd gnd FILL
X_12216_ _12216_/A _12216_/B _12216_/C _12216_/Y vdd gnd OAI21X1
X_13196_ _13196_/A _13196_/B _13196_/C _13196_/Y vdd gnd OAI21X1
XFILL_2__7524_ vdd gnd FILL
XFILL_1__11311_ vdd gnd FILL
XFILL_1__12291_ vdd gnd FILL
XFILL_2__10862_ vdd gnd FILL
X_12147_ _12147_/A _12147_/B _12147_/Y vdd gnd NAND2X1
XFILL_1__14030_ vdd gnd FILL
XFILL_2__7455_ vdd gnd FILL
XFILL_1__11242_ vdd gnd FILL
XFILL_0__14760_ vdd gnd FILL
XFILL_2__10793_ vdd gnd FILL
XFILL_0__11972_ vdd gnd FILL
X_12078_ _12078_/A _12078_/B _12078_/Y vdd gnd NOR2X1
XFILL_2__12532_ vdd gnd FILL
XFILL_0__13711_ vdd gnd FILL
XFILL_2__7386_ vdd gnd FILL
XFILL_0__10923_ vdd gnd FILL
XFILL_1__11173_ vdd gnd FILL
XFILL_0__14691_ vdd gnd FILL
X_11029_ _11029_/A _11029_/B _11029_/C _11029_/Y vdd gnd OAI21X1
XFILL_1__10124_ vdd gnd FILL
XFILL_2__12463_ vdd gnd FILL
XFILL_0__13642_ vdd gnd FILL
XFILL_0__10854_ vdd gnd FILL
XFILL_0__8140_ vdd gnd FILL
XFILL_1__10055_ vdd gnd FILL
XFILL_2__12394_ vdd gnd FILL
XFILL_0__13573_ vdd gnd FILL
XFILL_0__8071_ vdd gnd FILL
XFILL_0__10785_ vdd gnd FILL
XFILL_2__8007_ vdd gnd FILL
XFILL_0__12524_ vdd gnd FILL
XFILL_1__14863_ vdd gnd FILL
X_14719_ _14719_/A _14719_/B _14719_/Y vdd gnd NAND2X1
X_7650_ _7650_/A _7650_/B _7650_/Y vdd gnd NAND2X1
XFILL_1__13814_ vdd gnd FILL
XFILL_0__12455_ vdd gnd FILL
XFILL_1__14794_ vdd gnd FILL
X_7581_ _7581_/A _7581_/B _7581_/Y vdd gnd NAND2X1
XFILL_2__10227_ vdd gnd FILL
XFILL_2__13015_ vdd gnd FILL
XFILL_0__11406_ vdd gnd FILL
XFILL_1__13745_ vdd gnd FILL
XFILL_1__10957_ vdd gnd FILL
X_9320_ _9320_/A _9320_/B _9320_/C _9320_/Y vdd gnd OAI21X1
XFILL_0__12386_ vdd gnd FILL
XFILL_0__8973_ vdd gnd FILL
XFILL_2__10158_ vdd gnd FILL
XFILL_0__14125_ vdd gnd FILL
XFILL_0__11337_ vdd gnd FILL
XFILL_1__10888_ vdd gnd FILL
XFILL_1__13676_ vdd gnd FILL
X_9251_ _9251_/A _9251_/Y vdd gnd INVX1
XFILL_2__10089_ vdd gnd FILL
XFILL_1__12627_ vdd gnd FILL
XFILL_0__14056_ vdd gnd FILL
X_8202_ _8202_/A _8202_/B _8202_/C _8202_/D _8202_/Y vdd gnd AOI22X1
XFILL_0__11268_ vdd gnd FILL
X_9182_ _9182_/A _9182_/B _9182_/C _9182_/Y vdd gnd NAND3X1
XFILL_0__7855_ vdd gnd FILL
XFILL_0__13007_ vdd gnd FILL
XFILL_0__10219_ vdd gnd FILL
X_8133_ _8133_/A _8133_/B _8133_/S _8133_/Y vdd gnd MUX2X1
XFILL_0__11199_ vdd gnd FILL
XFILL_0__7786_ vdd gnd FILL
XFILL_1__11509_ vdd gnd FILL
XFILL_1__12489_ vdd gnd FILL
XFILL_0__9525_ vdd gnd FILL
X_8064_ _8064_/A _8064_/B _8064_/S _8064_/Y vdd gnd MUX2X1
XFILL_1__14228_ vdd gnd FILL
XFILL_0__9456_ vdd gnd FILL
XFILL_0__13909_ vdd gnd FILL
XFILL_1__7200_ vdd gnd FILL
XFILL_0__8407_ vdd gnd FILL
XFILL_0__9387_ vdd gnd FILL
XFILL_1__8180_ vdd gnd FILL
XFILL_1__7131_ vdd gnd FILL
XFILL_0__8338_ vdd gnd FILL
X_8966_ _8966_/A _8966_/B _8966_/Y vdd gnd NAND2X1
X_7917_ _7917_/D _7917_/CLK _7917_/Q vdd gnd DFFPOSX1
XFILL_0__8269_ vdd gnd FILL
X_8897_ _8897_/D _8897_/CLK _8897_/Q vdd gnd DFFPOSX1
XFILL_0_CLKBUF1_insert103 vdd gnd FILL
X_7848_ _7848_/A _7848_/B _7848_/C _7848_/Y vdd gnd OAI21X1
X_7779_ _7779_/A _7779_/B _7779_/Y vdd gnd NAND2X1
X_9518_ _9518_/A _9518_/B _9518_/Y vdd gnd NAND2X1
X_10400_ _10400_/A _10400_/B _10400_/C _10400_/Y vdd gnd OAI21X1
XFILL_1__9703_ vdd gnd FILL
X_11380_ _11380_/A _11380_/B _11380_/C _11380_/Y vdd gnd OAI21X1
X_9449_ _9449_/A _9449_/B _9449_/Y vdd gnd NAND2X1
XFILL_1__7895_ vdd gnd FILL
X_10331_ _10331_/A _10331_/B _10331_/C _10331_/Y vdd gnd NAND3X1
XFILL_1__9634_ vdd gnd FILL
X_10262_ _10262_/A _10262_/B _10262_/Y vdd gnd NAND2X1
X_13050_ _13050_/A _13050_/B _13050_/Y vdd gnd NOR2X1
XFILL_1__9565_ vdd gnd FILL
X_12001_ _12001_/A _12001_/B _12001_/C _12001_/Y vdd gnd OAI21X1
X_10193_ _10193_/A _10193_/Y vdd gnd INVX1
XFILL_1__8516_ vdd gnd FILL
XFILL_1__9496_ vdd gnd FILL
XFILL_1__8447_ vdd gnd FILL
X_13952_ _13952_/A _13952_/B _13952_/C _13952_/Y vdd gnd OAI21X1
XFILL_1__8378_ vdd gnd FILL
X_12903_ _12903_/A _12903_/B _12903_/Y vdd gnd AND2X2
XFILL_1__7329_ vdd gnd FILL
X_13883_ _13883_/A _13883_/B _13883_/C _13883_/Y vdd gnd OAI21X1
X_12834_ _12834_/A _12834_/B _12834_/C _12834_/Y vdd gnd OAI21X1
XFILL_0__10570_ vdd gnd FILL
X_12765_ _12765_/A _12765_/Y vdd gnd INVX2
XFILL_1__11860_ vdd gnd FILL
X_14504_ _14504_/D _14504_/CLK _14504_/Q vdd gnd DFFPOSX1
X_11716_ _11716_/A _11716_/Y vdd gnd INVX1
X_12696_ _12696_/A _12696_/B _12696_/Y vdd gnd NOR2X1
XFILL_0__12240_ vdd gnd FILL
XFILL_1__10811_ vdd gnd FILL
XFILL_1__11791_ vdd gnd FILL
X_14435_ _14435_/A _14435_/B _14435_/Y vdd gnd AND2X2
X_11647_ _11647_/D _11647_/CLK _11647_/Q vdd gnd DFFPOSX1
XFILL_2__9743_ vdd gnd FILL
XFILL_1__13530_ vdd gnd FILL
XFILL_0__12171_ vdd gnd FILL
X_14366_ _14366_/A _14366_/B _14366_/C _14366_/Y vdd gnd NAND3X1
XFILL_2__14820_ vdd gnd FILL
X_11578_ _11578_/A _11578_/B _11578_/C _11578_/Y vdd gnd OAI21X1
XFILL_2__9674_ vdd gnd FILL
XFILL_0__11122_ vdd gnd FILL
XFILL_1__10673_ vdd gnd FILL
X_13317_ _13317_/A _13317_/B _13317_/C _13317_/Y vdd gnd NAND3X1
X_10529_ _10529_/A _10529_/Y vdd gnd INVX1
XFILL_2_CLKBUF1_insert34 vdd gnd FILL
X_14297_ _14297_/A _14297_/B _14297_/Y vdd gnd NAND2X1
XFILL_2__14751_ vdd gnd FILL
XFILL_1__12412_ vdd gnd FILL
XFILL_0__11053_ vdd gnd FILL
XFILL_1__13392_ vdd gnd FILL
XFILL_2_CLKBUF1_insert67 vdd gnd FILL
XFILL_0__7640_ vdd gnd FILL
X_13248_ _13248_/A _13248_/Y vdd gnd INVX1
XFILL_2_CLKBUF1_insert89 vdd gnd FILL
XFILL_0__10004_ vdd gnd FILL
XFILL_1__12343_ vdd gnd FILL
XFILL_2__14682_ vdd gnd FILL
X_13179_ _13179_/A _13179_/B _13179_/C _13179_/Y vdd gnd OAI21X1
XFILL_0__7571_ vdd gnd FILL
XFILL_0__14812_ vdd gnd FILL
XFILL_1__12274_ vdd gnd FILL
XFILL_0__9310_ vdd gnd FILL
XFILL_1__14013_ vdd gnd FILL
XFILL_1__11225_ vdd gnd FILL
XFILL_0__14743_ vdd gnd FILL
XFILL_0__11955_ vdd gnd FILL
XFILL_0__9241_ vdd gnd FILL
XFILL_0_BUFX2_insert16 vdd gnd FILL
XFILL_2__12515_ vdd gnd FILL
XFILL_0_BUFX2_insert27 vdd gnd FILL
XFILL_0_CLKBUF1_insert60 vdd gnd FILL
XFILL_0_CLKBUF1_insert71 vdd gnd FILL
XFILL_0__10906_ vdd gnd FILL
XFILL_1__11156_ vdd gnd FILL
XFILL_0_CLKBUF1_insert82 vdd gnd FILL
XFILL_0__14674_ vdd gnd FILL
XFILL_0_CLKBUF1_insert93 vdd gnd FILL
XFILL_0__11886_ vdd gnd FILL
XFILL_0__9172_ vdd gnd FILL
X_8820_ _8820_/A _8820_/B _8820_/C _8820_/Y vdd gnd OAI21X1
XFILL_1__10107_ vdd gnd FILL
XFILL_2__12446_ vdd gnd FILL
XFILL_1__11087_ vdd gnd FILL
XFILL_0__10837_ vdd gnd FILL
XFILL_0__13625_ vdd gnd FILL
XFILL_0__8123_ vdd gnd FILL
X_8751_ _8751_/A _8751_/B _8751_/C _8751_/Y vdd gnd OAI21X1
XFILL_1__14915_ vdd gnd FILL
XFILL_1__10038_ vdd gnd FILL
XFILL_2__12377_ vdd gnd FILL
XFILL_0__13556_ vdd gnd FILL
XFILL_0__10768_ vdd gnd FILL
X_7702_ _7702_/A _7702_/B _7702_/C _7702_/Y vdd gnd OAI21X1
XFILL_0__8054_ vdd gnd FILL
XFILL_2__14116_ vdd gnd FILL
X_8682_ _8682_/A _8682_/B _8682_/Y vdd gnd NOR2X1
XFILL_0__12507_ vdd gnd FILL
XFILL_1__14846_ vdd gnd FILL
X_7633_ _7633_/A _7633_/B _7633_/C _7633_/Y vdd gnd AOI21X1
XFILL_2__14047_ vdd gnd FILL
XFILL_0__12438_ vdd gnd FILL
XFILL_1__14777_ vdd gnd FILL
XFILL_1__11989_ vdd gnd FILL
X_7564_ _7564_/A _7564_/B _7564_/C _7564_/Y vdd gnd AOI21X1
XFILL_1__13728_ vdd gnd FILL
XFILL_0__12369_ vdd gnd FILL
X_9303_ _9303_/A _9303_/B _9303_/C _9303_/Y vdd gnd OAI21X1
XFILL_0__8956_ vdd gnd FILL
X_7495_ _7495_/A _7495_/B _7495_/C _7495_/Y vdd gnd AOI21X1
XFILL_0__14108_ vdd gnd FILL
XFILL_1__13659_ vdd gnd FILL
XFILL_0__7907_ vdd gnd FILL
X_9234_ _9234_/A _9234_/B _9234_/C _9234_/Y vdd gnd NAND3X1
XFILL_1__7680_ vdd gnd FILL
XFILL_0__14039_ vdd gnd FILL
X_9165_ _9165_/A _9165_/B _9165_/Y vdd gnd NAND2X1
XFILL_0__7838_ vdd gnd FILL
X_8116_ _8116_/A _8116_/B _8116_/S _8116_/Y vdd gnd MUX2X1
XFILL_1__9350_ vdd gnd FILL
X_9096_ _9096_/A _9096_/Y vdd gnd INVX1
XFILL_0__7769_ vdd gnd FILL
XFILL_0__9508_ vdd gnd FILL
XFILL_1__8301_ vdd gnd FILL
X_8047_ _8047_/A _8047_/Y vdd gnd INVX1
XFILL_1__9281_ vdd gnd FILL
XFILL_0__9439_ vdd gnd FILL
XFILL_1__8232_ vdd gnd FILL
XFILL_1__8163_ vdd gnd FILL
X_9998_ _9998_/A _9998_/B _9998_/C _9998_/Y vdd gnd OAI21X1
XFILL_1__7114_ vdd gnd FILL
X_10880_ _10880_/A _10880_/B _10880_/C _10880_/Y vdd gnd OAI21X1
X_8949_ _8949_/A _8949_/B _8949_/C _8949_/Y vdd gnd OAI21X1
XFILL_1__8094_ vdd gnd FILL
X_12550_ _12550_/D _12550_/CLK _12550_/Q vdd gnd DFFPOSX1
X_11501_ _11501_/A _11501_/B _11501_/C _11501_/Y vdd gnd OAI21X1
X_12481_ _12481_/A _12481_/B _12481_/C _12481_/Y vdd gnd OAI21X1
XFILL_1__8996_ vdd gnd FILL
X_14220_ _14220_/A _14220_/B _14220_/Y vdd gnd NAND2X1
X_11432_ _11432_/A _11432_/B _11432_/Y vdd gnd NAND2X1
X_14151_ _14151_/A _14151_/B _14151_/C _14151_/Y vdd gnd OAI21X1
X_11363_ _11363_/A _11363_/B _11363_/Y vdd gnd AND2X2
XFILL_1__7878_ vdd gnd FILL
X_13102_ _13102_/A _13102_/Y vdd gnd INVX1
X_10314_ _10314_/A _10314_/B _10314_/C _10314_/Y vdd gnd NAND3X1
XFILL_1__9617_ vdd gnd FILL
XFILL_2__8410_ vdd gnd FILL
X_14082_ _14082_/A _14082_/B _14082_/Y vdd gnd NOR2X1
X_11294_ _11294_/A _11294_/B _11294_/C _11294_/Y vdd gnd OAI21X1
X_13033_ _13033_/A _13033_/Y vdd gnd INVX1
X_10245_ _10245_/A _10245_/B _10245_/C _10245_/Y vdd gnd NAND3X1
XFILL_1__9548_ vdd gnd FILL
XFILL_2__8341_ vdd gnd FILL
X_10176_ _10176_/A _10176_/B _10176_/Y vdd gnd AND2X2
XFILL_1__9479_ vdd gnd FILL
XFILL_2__10630_ vdd gnd FILL
XFILL_2__8272_ vdd gnd FILL
XFILL_1__11010_ vdd gnd FILL
XFILL_2__10561_ vdd gnd FILL
XFILL_0__11740_ vdd gnd FILL
X_13935_ _13935_/A _13935_/B _13935_/C _13935_/Y vdd gnd AOI21X1
XFILL_2__10492_ vdd gnd FILL
X_13866_ _13866_/A _13866_/B _13866_/Y vdd gnd NAND2X1
XFILL_0__13410_ vdd gnd FILL
XFILL_0__10622_ vdd gnd FILL
XFILL_1__12961_ vdd gnd FILL
XFILL_0__14390_ vdd gnd FILL
X_12817_ _12817_/A _12817_/Y vdd gnd INVX1
XFILL_1_BUFX2_insert330 vdd gnd FILL
XFILL_1_BUFX2_insert341 vdd gnd FILL
XFILL_1__14700_ vdd gnd FILL
X_13797_ _13797_/A _13797_/Y vdd gnd INVX1
XFILL_1__11912_ vdd gnd FILL
XFILL_0__13341_ vdd gnd FILL
XFILL_1_BUFX2_insert352 vdd gnd FILL
XFILL_1_BUFX2_insert363 vdd gnd FILL
XFILL_0__10553_ vdd gnd FILL
XFILL_1_BUFX2_insert374 vdd gnd FILL
XFILL_1__12892_ vdd gnd FILL
X_12748_ _12748_/A _12748_/B _12748_/S _12748_/Y vdd gnd MUX2X1
XFILL_2__11113_ vdd gnd FILL
XFILL_1__14631_ vdd gnd FILL
XFILL_2__12093_ vdd gnd FILL
XFILL_1__11843_ vdd gnd FILL
XFILL_0__13272_ vdd gnd FILL
XFILL_0__10484_ vdd gnd FILL
X_12679_ _12679_/A _12679_/B _12679_/Y vdd gnd NAND2X1
XFILL_0__12223_ vdd gnd FILL
XFILL_1__14562_ vdd gnd FILL
X_14418_ _14418_/A _14418_/B _14418_/C _14418_/Y vdd gnd NAND3X1
XFILL_0__8810_ vdd gnd FILL
XFILL_1__11774_ vdd gnd FILL
XFILL_1__13513_ vdd gnd FILL
XFILL_0__12154_ vdd gnd FILL
XFILL_1__14493_ vdd gnd FILL
XFILL_0__8741_ vdd gnd FILL
X_14349_ _14349_/A _14349_/B _14349_/C _14349_/Y vdd gnd OAI21X1
X_7280_ _7280_/A _7280_/Y vdd gnd INVX1
XFILL_2__14803_ vdd gnd FILL
XFILL_0__11105_ vdd gnd FILL
XFILL_1__10656_ vdd gnd FILL
XFILL_0__12085_ vdd gnd FILL
XFILL_2__8608_ vdd gnd FILL
XFILL_0__8672_ vdd gnd FILL
XFILL_2__14734_ vdd gnd FILL
XFILL_0__11036_ vdd gnd FILL
XFILL_2__11946_ vdd gnd FILL
XFILL_1__10587_ vdd gnd FILL
XFILL_1__13375_ vdd gnd FILL
XFILL_0__7623_ vdd gnd FILL
XFILL_2__8539_ vdd gnd FILL
XFILL257250x219750 vdd gnd FILL
XFILL_2__14665_ vdd gnd FILL
XFILL_1__12326_ vdd gnd FILL
XFILL_2__11877_ vdd gnd FILL
XFILL_0__7554_ vdd gnd FILL
XFILL_1__12257_ vdd gnd FILL
XFILL_2__14596_ vdd gnd FILL
X_9921_ _9921_/A _9921_/B _9921_/Y vdd gnd NOR2X1
XFILL_0__12987_ vdd gnd FILL
XFILL_0__7485_ vdd gnd FILL
XFILL_1__11208_ vdd gnd FILL
XFILL_0__14726_ vdd gnd FILL
XFILL_1__12188_ vdd gnd FILL
XFILL_0__9224_ vdd gnd FILL
XFILL_0__11938_ vdd gnd FILL
X_9852_ _9852_/A _9852_/Y vdd gnd INVX2
XFILL_1__11139_ vdd gnd FILL
XFILL_0__14657_ vdd gnd FILL
XFILL_0__11869_ vdd gnd FILL
XFILL_0__9155_ vdd gnd FILL
X_8803_ _8803_/A _8803_/B _8803_/C _8803_/Y vdd gnd OAI21X1
X_9783_ _9783_/D _9783_/CLK _9783_/Q vdd gnd DFFPOSX1
XFILL_2__12429_ vdd gnd FILL
XFILL_0__13608_ vdd gnd FILL
XFILL_0__8106_ vdd gnd FILL
XFILL_0__14588_ vdd gnd FILL
XFILL_0__9086_ vdd gnd FILL
X_8734_ _8734_/A _8734_/B _8734_/C _8734_/Y vdd gnd AOI21X1
XFILL_0__13539_ vdd gnd FILL
XFILL_0__8037_ vdd gnd FILL
X_8665_ _8665_/A _8665_/B _8665_/Y vdd gnd OR2X2
XFILL_1__14829_ vdd gnd FILL
X_7616_ _7616_/A _7616_/Y vdd gnd INVX1
X_8596_ _8596_/A _8596_/B _8596_/Y vdd gnd NOR2X1
XFILL_1__7801_ vdd gnd FILL
X_7547_ _7547_/A _7547_/B _7547_/Y vdd gnd OR2X2
XFILL_0__9988_ vdd gnd FILL
XFILL_1__8781_ vdd gnd FILL
XFILL_0__8939_ vdd gnd FILL
XFILL_1__7732_ vdd gnd FILL
X_7478_ _7478_/A _7478_/Y vdd gnd INVX1
X_9217_ _9217_/A _9217_/B _9217_/C _9217_/Y vdd gnd OAI21X1
XFILL_1__7663_ vdd gnd FILL
XFILL_1__9402_ vdd gnd FILL
XFILL256650x144150 vdd gnd FILL
X_9148_ _9148_/A _9148_/Y vdd gnd INVX1
XFILL257250x129750 vdd gnd FILL
XFILL_1__7594_ vdd gnd FILL
X_10030_ _10030_/A _10030_/Y vdd gnd INVX1
XFILL_1__9333_ vdd gnd FILL
X_9079_ _9079_/A _9079_/Y vdd gnd INVX1
XFILL_1__9264_ vdd gnd FILL
XFILL_1__8215_ vdd gnd FILL
X_11981_ _11981_/A _11981_/B _11981_/C _11981_/Y vdd gnd OAI21X1
XFILL_1__9195_ vdd gnd FILL
X_13720_ _13720_/A _13720_/Y vdd gnd INVX1
X_10932_ _10932_/A _10932_/B _10932_/C _10932_/Y vdd gnd NAND3X1
XFILL_1__8146_ vdd gnd FILL
XFILL_0_BUFX2_insert8 vdd gnd FILL
X_13651_ _13651_/A _13651_/Y vdd gnd INVX1
X_10863_ _10863_/A _10863_/B _10863_/C _10863_/Y vdd gnd NAND3X1
XFILL_1__8077_ vdd gnd FILL
X_12602_ _12602_/D _12602_/CLK _12602_/Q vdd gnd DFFPOSX1
X_13582_ _13582_/A _13582_/B _13582_/C _13582_/Y vdd gnd NAND3X1
X_10794_ _10794_/A _10794_/B _10794_/C _10794_/Y vdd gnd AOI21X1
XFILL_0_BUFX2_insert304 vdd gnd FILL
XFILL_0_BUFX2_insert315 vdd gnd FILL
XFILL_0_BUFX2_insert326 vdd gnd FILL
X_12533_ _12533_/A _12533_/B _12533_/C _12533_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert337 vdd gnd FILL
XFILL_2__7841_ vdd gnd FILL
XFILL_0_BUFX2_insert348 vdd gnd FILL
XFILL_0_BUFX2_insert359 vdd gnd FILL
X_12464_ _12464_/A _12464_/B _12464_/C _12464_/Y vdd gnd OAI21X1
XFILL_2__7772_ vdd gnd FILL
XFILL_1__8979_ vdd gnd FILL
X_14203_ _14203_/D _14203_/CLK _14203_/Q vdd gnd DFFPOSX1
X_11415_ _11415_/A _11415_/B _11415_/Y vdd gnd NAND2X1
XFILL_1__10510_ vdd gnd FILL
X_12395_ _12395_/A _12395_/B _12395_/Y vdd gnd NAND2X1
XFILL_1__11490_ vdd gnd FILL
X_14134_ _14134_/A _14134_/B _14134_/C _14134_/Y vdd gnd OAI21X1
X_11346_ _11346_/A _11346_/B _11346_/Y vdd gnd NAND2X1
XFILL_2__11800_ vdd gnd FILL
XFILL_1__10441_ vdd gnd FILL
X_14065_ _14065_/A _14065_/B _14065_/Y vdd gnd AND2X2
X_11277_ _11277_/A _11277_/B _11277_/Y vdd gnd NAND2X1
XFILL_1__13160_ vdd gnd FILL
XFILL_2__11731_ vdd gnd FILL
XFILL_1__10372_ vdd gnd FILL
XFILL_0__12910_ vdd gnd FILL
X_13016_ _13016_/A _13016_/B _13016_/C _13016_/Y vdd gnd NAND3X1
XFILL_0__13890_ vdd gnd FILL
X_10228_ _10228_/A _10228_/B _10228_/C _10228_/Y vdd gnd OAI21X1
XFILL_2__8324_ vdd gnd FILL
XFILL_1__12111_ vdd gnd FILL
XFILL_1__13091_ vdd gnd FILL
XFILL_0__12841_ vdd gnd FILL
X_10159_ _10159_/A _10159_/B _10159_/C _10159_/Y vdd gnd OAI21X1
XFILL_2__13401_ vdd gnd FILL
XFILL_2__10613_ vdd gnd FILL
XFILL_2__8255_ vdd gnd FILL
XFILL_1__12042_ vdd gnd FILL
XFILL_0__12772_ vdd gnd FILL
XFILL_0__7270_ vdd gnd FILL
XFILL_2__13332_ vdd gnd FILL
XFILL_2__10544_ vdd gnd FILL
XFILL_0__11723_ vdd gnd FILL
XFILL_2__8186_ vdd gnd FILL
X_13918_ _13918_/A _13918_/B _13918_/Y vdd gnd AND2X2
X_14898_ _14898_/D _14898_/CLK _14898_/Q vdd gnd DFFPOSX1
XFILL_2__10475_ vdd gnd FILL
XFILL_0__14442_ vdd gnd FILL
XFILL_1__13993_ vdd gnd FILL
X_13849_ _13849_/A _13849_/Y vdd gnd INVX1
XFILL_0__10605_ vdd gnd FILL
XFILL_1__12944_ vdd gnd FILL
XFILL_0__14373_ vdd gnd FILL
XFILL_1_BUFX2_insert160 vdd gnd FILL
XFILL_0__11585_ vdd gnd FILL
XFILL_1_BUFX2_insert171 vdd gnd FILL
XFILL_1_BUFX2_insert182 vdd gnd FILL
XFILL_0__13324_ vdd gnd FILL
XFILL_0__10536_ vdd gnd FILL
XFILL_1_BUFX2_insert193 vdd gnd FILL
XFILL_0__9911_ vdd gnd FILL
XFILL_1__12875_ vdd gnd FILL
X_8450_ _8450_/A _8450_/B _8450_/Y vdd gnd NAND2X1
XFILL_1__14614_ vdd gnd FILL
XFILL_1__11826_ vdd gnd FILL
XFILL_0__13255_ vdd gnd FILL
XFILL_0__10467_ vdd gnd FILL
X_7401_ _7401_/A _7401_/B _7401_/C _7401_/Y vdd gnd OAI21X1
X_8381_ _8381_/A _8381_/B _8381_/Y vdd gnd NAND2X1
XFILL_2__11027_ vdd gnd FILL
XFILL_0__12206_ vdd gnd FILL
XFILL_0__13186_ vdd gnd FILL
XFILL_1__11757_ vdd gnd FILL
XFILL_0__10398_ vdd gnd FILL
X_7332_ _7332_/A _7332_/Y vdd gnd INVX1
XFILL_0__12137_ vdd gnd FILL
XFILL_1__14476_ vdd gnd FILL
XFILL_0__8724_ vdd gnd FILL
X_7263_ _7263_/A _7263_/B _7263_/C _7263_/Y vdd gnd OAI21X1
XFILL_1__13427_ vdd gnd FILL
XFILL_1__10639_ vdd gnd FILL
XFILL_0__12068_ vdd gnd FILL
X_9002_ _9002_/A _9002_/Y vdd gnd INVX2
XFILL_0__8655_ vdd gnd FILL
X_7194_ _7194_/A _7194_/B _7194_/S _7194_/Y vdd gnd MUX2X1
XFILL_2__14717_ vdd gnd FILL
XFILL_0__11019_ vdd gnd FILL
XFILL_2__11929_ vdd gnd FILL
XFILL_1__13358_ vdd gnd FILL
XFILL_0__7606_ vdd gnd FILL
XFILL_0__8586_ vdd gnd FILL
XFILL_2__14648_ vdd gnd FILL
XFILL_1__12309_ vdd gnd FILL
XFILL_1__13289_ vdd gnd FILL
XFILL_0__7537_ vdd gnd FILL
XFILL_2__14579_ vdd gnd FILL
X_9904_ _9904_/A _9904_/Y vdd gnd INVX8
XFILL_0__7468_ vdd gnd FILL
XFILL_0__14709_ vdd gnd FILL
XFILL_0__9207_ vdd gnd FILL
XFILL_1__8000_ vdd gnd FILL
X_9835_ _9835_/D _9835_/CLK _9835_/Q vdd gnd DFFPOSX1
XFILL_0__7399_ vdd gnd FILL
XFILL_0__9138_ vdd gnd FILL
X_9766_ _9766_/D _9766_/CLK _9766_/Q vdd gnd DFFPOSX1
XFILL_0__9069_ vdd gnd FILL
XFILL_1__9951_ vdd gnd FILL
XFILL257250x104550 vdd gnd FILL
X_8717_ _8717_/A _8717_/B _8717_/C _8717_/D _8717_/Y vdd gnd AOI22X1
X_9697_ _9697_/A _9697_/B _9697_/Y vdd gnd NAND2X1
XFILL_1__9882_ vdd gnd FILL
X_8648_ _8648_/A _8648_/Y vdd gnd INVX1
XFILL_1__8833_ vdd gnd FILL
X_8579_ _8579_/A _8579_/Y vdd gnd INVX1
XFILL_1__8764_ vdd gnd FILL
X_11200_ _11200_/A _11200_/B _11200_/Y vdd gnd AND2X2
XFILL_1__7715_ vdd gnd FILL
X_12180_ _12180_/A _12180_/B _12180_/Y vdd gnd NOR2X1
XFILL_1__8695_ vdd gnd FILL
X_11131_ _11131_/A _11131_/Y vdd gnd INVX1
XFILL_1__7646_ vdd gnd FILL
X_11062_ _11062_/A _11062_/B _11062_/Y vdd gnd AND2X2
XFILL_1__7577_ vdd gnd FILL
X_10013_ _10013_/A _10013_/B _10013_/C _10013_/Y vdd gnd OAI21X1
XFILL_1__9316_ vdd gnd FILL
X_14821_ _14821_/A _14821_/B _14821_/Y vdd gnd NOR2X1
XFILL_1__9247_ vdd gnd FILL
X_14752_ _14752_/A _14752_/B _14752_/Y vdd gnd OR2X2
X_11964_ _11964_/A _11964_/B _11964_/Y vdd gnd NOR2X1
XFILL_1__9178_ vdd gnd FILL
X_13703_ _13703_/A _13703_/Y vdd gnd INVX1
X_10915_ _10915_/A _10915_/B _10915_/Y vdd gnd NAND2X1
X_14683_ _14683_/A _14683_/B _14683_/Y vdd gnd NOR2X1
XFILL_1__8129_ vdd gnd FILL
XFILL_2__10260_ vdd gnd FILL
X_11895_ _11895_/A _11895_/B _11895_/Y vdd gnd NAND2X1
X_13634_ _13634_/A _13634_/B _13634_/C _13634_/Y vdd gnd AOI21X1
XFILL_1__10990_ vdd gnd FILL
X_10846_ _10846_/A _10846_/B _10846_/Y vdd gnd NAND2X1
XFILL_2__10191_ vdd gnd FILL
XFILL_0__11370_ vdd gnd FILL
XFILL_0_BUFX2_insert112 vdd gnd FILL
X_13565_ _13565_/A _13565_/Y vdd gnd INVX1
XFILL_0_BUFX2_insert123 vdd gnd FILL
X_10777_ _10777_/A _10777_/B _10777_/Y vdd gnd AND2X2
XFILL_0_BUFX2_insert134 vdd gnd FILL
XFILL_0__10321_ vdd gnd FILL
XFILL_0_BUFX2_insert145 vdd gnd FILL
XFILL_1__12660_ vdd gnd FILL
X_12516_ _12516_/A _12516_/B _12516_/C _12516_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert156 vdd gnd FILL
XFILL_0_BUFX2_insert167 vdd gnd FILL
X_13496_ _13496_/D _13496_/CLK _13496_/Q vdd gnd DFFPOSX1
XFILL_0_BUFX2_insert178 vdd gnd FILL
XFILL_1__11611_ vdd gnd FILL
XFILL_0__13040_ vdd gnd FILL
XFILL_0_BUFX2_insert189 vdd gnd FILL
XFILL_0__10252_ vdd gnd FILL
X_12447_ _12447_/A _12447_/B _12447_/C _12447_/Y vdd gnd OAI21X1
XFILL_1__14330_ vdd gnd FILL
XFILL_1__11542_ vdd gnd FILL
XFILL_0__10183_ vdd gnd FILL
X_12378_ _12378_/A _12378_/B _12378_/Y vdd gnd NOR2X1
XFILL_1__14261_ vdd gnd FILL
XFILL_1__11473_ vdd gnd FILL
X_14117_ _14117_/A _14117_/B _14117_/C _14117_/Y vdd gnd OAI21X1
X_11329_ _11329_/A _11329_/B _11329_/C _11329_/Y vdd gnd AOI21X1
XFILL_1__13212_ vdd gnd FILL
XFILL_1__10424_ vdd gnd FILL
XFILL_0__13942_ vdd gnd FILL
XFILL_0__8440_ vdd gnd FILL
X_14048_ _14048_/A _14048_/B _14048_/C _14048_/Y vdd gnd OAI21X1
XFILL_2__11714_ vdd gnd FILL
XFILL_1__13143_ vdd gnd FILL
XFILL_1__10355_ vdd gnd FILL
XFILL_0__13873_ vdd gnd FILL
XFILL_0__8371_ vdd gnd FILL
XFILL_2__14433_ vdd gnd FILL
XFILL_1__10286_ vdd gnd FILL
XFILL_0__12824_ vdd gnd FILL
XFILL_1__13074_ vdd gnd FILL
XFILL_0__7322_ vdd gnd FILL
X_7950_ _7950_/D _7950_/CLK _7950_/Q vdd gnd DFFPOSX1
XFILL_2__8238_ vdd gnd FILL
XFILL_1__12025_ vdd gnd FILL
XFILL_0__12755_ vdd gnd FILL
XFILL_0__7253_ vdd gnd FILL
XFILL_2__13315_ vdd gnd FILL
X_7881_ _7881_/A _7881_/B _7881_/C _7881_/Y vdd gnd OAI21X1
XFILL_2__10527_ vdd gnd FILL
XFILL_2__8169_ vdd gnd FILL
XFILL_0__11706_ vdd gnd FILL
X_9620_ _9620_/A _9620_/B _9620_/Y vdd gnd NAND2X1
XFILL_0__12686_ vdd gnd FILL
XFILL_0__7184_ vdd gnd FILL
XFILL_2__13246_ vdd gnd FILL
XFILL_2__10458_ vdd gnd FILL
XFILL_0__14425_ vdd gnd FILL
XFILL_1__13976_ vdd gnd FILL
X_9551_ _9551_/A _9551_/B _9551_/Y vdd gnd NAND2X1
XFILL_2__13177_ vdd gnd FILL
XFILL_1__12927_ vdd gnd FILL
XFILL_2__10389_ vdd gnd FILL
XFILL_0__14356_ vdd gnd FILL
XFILL_0__11568_ vdd gnd FILL
X_8502_ _8502_/A _8502_/B _8502_/C _8502_/Y vdd gnd NOR3X1
X_9482_ _9482_/A _9482_/B _9482_/C _9482_/Y vdd gnd OAI21X1
XFILL_0__10519_ vdd gnd FILL
XFILL_0__13307_ vdd gnd FILL
XFILL_1__12858_ vdd gnd FILL
XFILL_0__14287_ vdd gnd FILL
XBUFX2_insert18 BUFX2_insert18/A BUFX2_insert18/Y vdd gnd BUFX2
XFILL_0__11499_ vdd gnd FILL
X_8433_ _8433_/A _8433_/Y vdd gnd INVX1
XFILL_1__11809_ vdd gnd FILL
XFILL_0__13238_ vdd gnd FILL
XFILL_1__12789_ vdd gnd FILL
X_8364_ _8364_/A _8364_/B _8364_/Y vdd gnd NOR2X1
XFILL_0__13169_ vdd gnd FILL
X_7315_ _7315_/A _7315_/B _7315_/Y vdd gnd NOR2X1
XFILL_0__9756_ vdd gnd FILL
X_8295_ _8295_/A _8295_/B _8295_/Y vdd gnd NAND2X1
XFILL_1__14459_ vdd gnd FILL
XFILL_1__7500_ vdd gnd FILL
XFILL_0__8707_ vdd gnd FILL
X_7246_ _7246_/A _7246_/B _7246_/C _7246_/Y vdd gnd NAND3X1
XFILL_0__9687_ vdd gnd FILL
XFILL_1__8480_ vdd gnd FILL
XFILL_1__7431_ vdd gnd FILL
XFILL_0__8638_ vdd gnd FILL
X_7177_ _7177_/A _7177_/B _7177_/C _7177_/Y vdd gnd OAI21X1
XFILL_1__7362_ vdd gnd FILL
XFILL_0__8569_ vdd gnd FILL
XCLKBUF1_insert391 CLKBUF1_insert391/A CLKBUF1_insert391/Y vdd gnd CLKBUF1
XFILL_1__9101_ vdd gnd FILL
XFILL_2_BUFX2_insert218 vdd gnd FILL
XFILL_2_BUFX2_insert229 vdd gnd FILL
XFILL_1__7293_ vdd gnd FILL
XFILL_1__9032_ vdd gnd FILL
X_9818_ _9818_/D _9818_/CLK _9818_/Q vdd gnd DFFPOSX1
X_10700_ _10700_/D _10700_/CLK _10700_/Q vdd gnd DFFPOSX1
X_11680_ _11680_/D _11680_/CLK _11680_/Q vdd gnd DFFPOSX1
X_9749_ _9749_/A _9749_/B _9749_/C _9749_/Y vdd gnd OAI21X1
XBUFX2_insert206 BUFX2_insert206/A BUFX2_insert206/Y vdd gnd BUFX2
X_10631_ _10631_/A _10631_/B _10631_/C _10631_/Y vdd gnd OAI21X1
XBUFX2_insert217 BUFX2_insert217/A BUFX2_insert217/Y vdd gnd BUFX2
XBUFX2_insert228 BUFX2_insert228/A BUFX2_insert228/Y vdd gnd BUFX2
XFILL_1__9934_ vdd gnd FILL
XBUFX2_insert239 BUFX2_insert239/A BUFX2_insert239/Y vdd gnd BUFX2
X_13350_ _13350_/A _13350_/B _13350_/C _13350_/Y vdd gnd OAI21X1
X_10562_ _10562_/A _10562_/B _10562_/Y vdd gnd NAND2X1
XFILL_1__9865_ vdd gnd FILL
X_12301_ _12301_/A _12301_/B _12301_/Y vdd gnd NOR2X1
X_13281_ _13281_/A _13281_/B _13281_/Y vdd gnd NAND2X1
X_10493_ _10493_/A _10493_/B _10493_/Y vdd gnd NOR2X1
XFILL_1__8816_ vdd gnd FILL
X_12232_ _12232_/A _12232_/B _12232_/C _12232_/Y vdd gnd NAND3X1
XFILL_1__8747_ vdd gnd FILL
X_12163_ _12163_/A _12163_/B _12163_/Y vdd gnd OR2X2
XFILL_1__8678_ vdd gnd FILL
X_11114_ _11114_/A _11114_/B _11114_/Y vdd gnd NAND2X1
XFILL_2__9210_ vdd gnd FILL
XFILL_1__7629_ vdd gnd FILL
X_12094_ _12094_/A _12094_/B _12094_/S _12094_/Y vdd gnd MUX2X1
X_11045_ _11045_/A _11045_/B _11045_/C _11045_/Y vdd gnd OAI21X1
XFILL_2__9141_ vdd gnd FILL
XFILL_1__10140_ vdd gnd FILL
XFILL_0__10870_ vdd gnd FILL
XFILL_2__11430_ vdd gnd FILL
XFILL_1__10071_ vdd gnd FILL
X_14804_ _14804_/A _14804_/B _14804_/C _14804_/Y vdd gnd AOI21X1
X_12996_ _12996_/A _12996_/B _12996_/Y vdd gnd NAND2X1
XFILL_2__13100_ vdd gnd FILL
X_14735_ _14735_/A _14735_/B _14735_/Y vdd gnd NOR2X1
X_11947_ _11947_/A _11947_/B _11947_/C _11947_/Y vdd gnd AOI21X1
XFILL_2__14080_ vdd gnd FILL
XFILL_1__13830_ vdd gnd FILL
XFILL_0__12471_ vdd gnd FILL
X_14666_ _14666_/A _14666_/Y vdd gnd INVX1
X_11878_ _11878_/A _11878_/Y vdd gnd INVX1
XFILL_2__13031_ vdd gnd FILL
XFILL_0__11422_ vdd gnd FILL
XFILL_2__9974_ vdd gnd FILL
XFILL_1__13761_ vdd gnd FILL
XFILL_1__10973_ vdd gnd FILL
X_13617_ _13617_/A _13617_/B _13617_/C _13617_/Y vdd gnd OAI21X1
X_10829_ _10829_/A _10829_/Y vdd gnd INVX8
X_14597_ _14597_/A _14597_/B _14597_/Y vdd gnd AND2X2
XFILL_1__12712_ vdd gnd FILL
XFILL_0__11353_ vdd gnd FILL
XFILL_0__14141_ vdd gnd FILL
XFILL_1__13692_ vdd gnd FILL
X_13548_ _13548_/A _13548_/Y vdd gnd INVX1
XFILL_0__10304_ vdd gnd FILL
XFILL_1__12643_ vdd gnd FILL
XFILL_0__14072_ vdd gnd FILL
XFILL_0__11284_ vdd gnd FILL
XFILL_0__7871_ vdd gnd FILL
X_13479_ _13479_/D _13479_/CLK _13479_/Q vdd gnd DFFPOSX1
XFILL_0__13023_ vdd gnd FILL
XFILL_0__10235_ vdd gnd FILL
XFILL_2__8787_ vdd gnd FILL
XFILL_0__9610_ vdd gnd FILL
XFILL_1__14313_ vdd gnd FILL
XFILL_1__11525_ vdd gnd FILL
XFILL_0__10166_ vdd gnd FILL
X_7100_ _7100_/A _7100_/B _7100_/Y vdd gnd NAND2X1
XFILL_0__9541_ vdd gnd FILL
X_8080_ _8080_/A _8080_/B _8080_/C _8080_/Y vdd gnd OAI21X1
XFILL_1__14244_ vdd gnd FILL
XFILL_1__11456_ vdd gnd FILL
XFILL_0__10097_ vdd gnd FILL
XFILL_0__9472_ vdd gnd FILL
XFILL_1__10407_ vdd gnd FILL
XFILL_0__13925_ vdd gnd FILL
XFILL_0__8423_ vdd gnd FILL
XFILL_1__11387_ vdd gnd FILL
XFILL_1__13126_ vdd gnd FILL
XFILL_1__10338_ vdd gnd FILL
XFILL_0__13856_ vdd gnd FILL
XFILL_0__8354_ vdd gnd FILL
XFILL_2__14416_ vdd gnd FILL
X_8982_ _8982_/A _8982_/Y vdd gnd INVX1
XFILL_1__13057_ vdd gnd FILL
XFILL_1__10269_ vdd gnd FILL
XFILL_0__12807_ vdd gnd FILL
XFILL_0__7305_ vdd gnd FILL
XFILL_0__13787_ vdd gnd FILL
X_7933_ _7933_/D _7933_/CLK _7933_/Q vdd gnd DFFPOSX1
XFILL_0__8285_ vdd gnd FILL
XFILL_0__10999_ vdd gnd FILL
XFILL_2__14347_ vdd gnd FILL
XFILL_1__12008_ vdd gnd FILL
XFILL_0__12738_ vdd gnd FILL
XFILL_0__7236_ vdd gnd FILL
X_7864_ _7864_/A _7864_/B _7864_/Y vdd gnd NAND2X1
XFILL_2__14278_ vdd gnd FILL
X_9603_ _9603_/A _9603_/B _9603_/Y vdd gnd NAND2X1
XFILL_0__12669_ vdd gnd FILL
XFILL_0__7167_ vdd gnd FILL
XFILL_2__13229_ vdd gnd FILL
X_7795_ _7795_/A _7795_/B _7795_/Y vdd gnd NOR2X1
XFILL_0__14408_ vdd gnd FILL
XFILL_1__13959_ vdd gnd FILL
X_9534_ _9534_/A _9534_/B _9534_/C _9534_/Y vdd gnd OAI21X1
XFILL_0__7098_ vdd gnd FILL
XFILL_0__14339_ vdd gnd FILL
X_9465_ _9465_/A _9465_/B _9465_/C _9465_/Y vdd gnd AOI21X1
XFILL_1__9650_ vdd gnd FILL
X_8416_ _8416_/A _8416_/B _8416_/Y vdd gnd NAND2X1
X_9396_ _9396_/A _9396_/B _9396_/Y vdd gnd NAND2X1
XFILL_1__8601_ vdd gnd FILL
XFILL_1__9581_ vdd gnd FILL
X_8347_ _8347_/A _8347_/B _8347_/Y vdd gnd NAND2X1
XFILL_1__8532_ vdd gnd FILL
XFILL_0__9739_ vdd gnd FILL
X_8278_ _8278_/A _8278_/B _8278_/C _8278_/Y vdd gnd AOI21X1
X_7229_ _7229_/A _7229_/B _7229_/C _7229_/Y vdd gnd OAI21X1
XFILL_1__8463_ vdd gnd FILL
XFILL_1__7414_ vdd gnd FILL
XFILL_1__8394_ vdd gnd FILL
XFILL_1__7345_ vdd gnd FILL
X_12850_ _12850_/A _12850_/B _12850_/Y vdd gnd NAND2X1
XFILL_1__7276_ vdd gnd FILL
X_11801_ _11801_/A _11801_/B _11801_/C _11801_/Y vdd gnd OAI21X1
XFILL_1__9015_ vdd gnd FILL
X_12781_ _12781_/A _12781_/B _12781_/C _12781_/D _12781_/Y vdd gnd AOI22X1
X_14520_ _14520_/D _14520_/CLK _14520_/Q vdd gnd DFFPOSX1
X_11732_ _11732_/A _11732_/B _11732_/C _11732_/D _11732_/Y vdd gnd AOI22X1
X_14451_ _14451_/A _14451_/B _14451_/C _14451_/Y vdd gnd OAI21X1
X_11663_ _11663_/D _11663_/CLK _11663_/Q vdd gnd DFFPOSX1
X_13402_ _13402_/A _13402_/B _13402_/Y vdd gnd NAND2X1
X_10614_ _10614_/A _10614_/B _10614_/C _10614_/Y vdd gnd OAI21X1
X_14382_ _14382_/A _14382_/B _14382_/Y vdd gnd NOR2X1
XFILL_1__9917_ vdd gnd FILL
XFILL_2__8710_ vdd gnd FILL
X_11594_ _11594_/A _11594_/B _11594_/C _11594_/Y vdd gnd OAI21X1
X_13333_ _13333_/A _13333_/B _13333_/C _13333_/Y vdd gnd OAI21X1
X_10545_ _10545_/A _10545_/B _10545_/Y vdd gnd NAND2X1
XFILL_2__8641_ vdd gnd FILL
XFILL_1__9848_ vdd gnd FILL
X_13264_ _13264_/A _13264_/B _13264_/Y vdd gnd NOR2X1
X_10476_ _10476_/A _10476_/B _10476_/Y vdd gnd NOR2X1
XFILL_0__10020_ vdd gnd FILL
XFILL_2__8572_ vdd gnd FILL
X_12215_ _12215_/A _12215_/B _12215_/Y vdd gnd NOR2X1
X_13195_ _13195_/A _13195_/B _13195_/C _13195_/Y vdd gnd NAND3X1
XFILL_1__11310_ vdd gnd FILL
XFILL_1__12290_ vdd gnd FILL
X_12146_ _12146_/A _12146_/B _12146_/Y vdd gnd NAND2X1
XFILL_1__11241_ vdd gnd FILL
XFILL_2__13580_ vdd gnd FILL
XFILL_0__11971_ vdd gnd FILL
X_12077_ _12077_/A _12077_/B _12077_/Y vdd gnd NAND2X1
XFILL_0__13710_ vdd gnd FILL
XFILL_1__11172_ vdd gnd FILL
XFILL_0__10922_ vdd gnd FILL
X_11028_ _11028_/A _11028_/Y vdd gnd INVX1
XFILL_0__14690_ vdd gnd FILL
XFILL_2__9124_ vdd gnd FILL
XFILL_1__10123_ vdd gnd FILL
XFILL_0__13641_ vdd gnd FILL
XFILL_0__10853_ vdd gnd FILL
XFILL_2__9055_ vdd gnd FILL
XFILL_2__11413_ vdd gnd FILL
XFILL_1__10054_ vdd gnd FILL
XFILL_0__10784_ vdd gnd FILL
XFILL_0__13572_ vdd gnd FILL
XFILL_0__8070_ vdd gnd FILL
X_12979_ _12979_/A _12979_/B _12979_/C _12979_/Y vdd gnd NAND3X1
XFILL_2__14132_ vdd gnd FILL
XFILL_2__11344_ vdd gnd FILL
XFILL_1__14862_ vdd gnd FILL
XFILL_0__12523_ vdd gnd FILL
X_14718_ _14718_/A _14718_/B _14718_/Y vdd gnd NOR2X1
XFILL_2__14063_ vdd gnd FILL
XFILL_1__13813_ vdd gnd FILL
XFILL_2__11275_ vdd gnd FILL
XFILL_1__14793_ vdd gnd FILL
XFILL_0__12454_ vdd gnd FILL
X_14649_ _14649_/A _14649_/B _14649_/Y vdd gnd AND2X2
X_7580_ _7580_/A _7580_/B _7580_/C _7580_/Y vdd gnd OAI21X1
XFILL_2__9957_ vdd gnd FILL
XFILL_0__11405_ vdd gnd FILL
XFILL_1__13744_ vdd gnd FILL
XFILL_1__10956_ vdd gnd FILL
XFILL_0__12385_ vdd gnd FILL
XFILL_0__8972_ vdd gnd FILL
XFILL_0__11336_ vdd gnd FILL
XFILL_0__14124_ vdd gnd FILL
XFILL_2__9888_ vdd gnd FILL
XFILL_1__13675_ vdd gnd FILL
XFILL_1__10887_ vdd gnd FILL
X_9250_ _9250_/A _9250_/B _9250_/Y vdd gnd NAND2X1
XFILL_2__8839_ vdd gnd FILL
XFILL_1__12626_ vdd gnd FILL
XFILL_0__11267_ vdd gnd FILL
XFILL_0__14055_ vdd gnd FILL
X_8201_ _8201_/A _8201_/B _8201_/C _8201_/Y vdd gnd OAI21X1
XFILL_0__7854_ vdd gnd FILL
X_9181_ _9181_/A _9181_/B _9181_/C _9181_/Y vdd gnd OAI21X1
XFILL_2__13916_ vdd gnd FILL
XFILL_0__10218_ vdd gnd FILL
XFILL_0__13006_ vdd gnd FILL
XFILL_0__11198_ vdd gnd FILL
X_8132_ _8132_/A _8132_/B _8132_/C _8132_/Y vdd gnd AOI21X1
XFILL_0__7785_ vdd gnd FILL
XFILL_1__11508_ vdd gnd FILL
XFILL_0__10149_ vdd gnd FILL
XFILL_0__9524_ vdd gnd FILL
XFILL_1__12488_ vdd gnd FILL
X_8063_ _8063_/A _8063_/B _8063_/C _8063_/Y vdd gnd OAI21X1
XFILL_1__14227_ vdd gnd FILL
XFILL_1__11439_ vdd gnd FILL
XFILL_0__9455_ vdd gnd FILL
XFILL_2__12729_ vdd gnd FILL
XFILL_0__13908_ vdd gnd FILL
XFILL_1__14158_ vdd gnd FILL
XFILL_0__8406_ vdd gnd FILL
XFILL_0__9386_ vdd gnd FILL
XFILL_1__13109_ vdd gnd FILL
XFILL_1__14089_ vdd gnd FILL
XFILL_0__13839_ vdd gnd FILL
XFILL_1__7130_ vdd gnd FILL
XFILL_0__8337_ vdd gnd FILL
X_8965_ _8965_/A _8965_/Y vdd gnd INVX1
X_7916_ _7916_/D _7916_/CLK _7916_/Q vdd gnd DFFPOSX1
XFILL_0__8268_ vdd gnd FILL
X_8896_ _8896_/D _8896_/CLK _8896_/Q vdd gnd DFFPOSX1
XFILL_0__7219_ vdd gnd FILL
X_7847_ _7847_/A _7847_/B _7847_/Y vdd gnd NAND2X1
XFILL_0__8199_ vdd gnd FILL
XFILL_0_CLKBUF1_insert104 vdd gnd FILL
X_7778_ _7778_/A _7778_/B _7778_/Y vdd gnd NAND2X1
X_9517_ _9517_/A _9517_/B _9517_/C _9517_/Y vdd gnd OAI21X1
XFILL_1__9702_ vdd gnd FILL
X_9448_ _9448_/A _9448_/Y vdd gnd INVX1
XFILL_1__7894_ vdd gnd FILL
X_10330_ _10330_/A _10330_/Y vdd gnd INVX1
XFILL_1__9633_ vdd gnd FILL
X_9379_ _9379_/A _9379_/B _9379_/C _9379_/Y vdd gnd OAI21X1
X_10261_ _10261_/A _10261_/B _10261_/C _10261_/Y vdd gnd OAI21X1
XFILL_1__9564_ vdd gnd FILL
X_12000_ _12000_/A _12000_/Y vdd gnd INVX1
XFILL_1__8515_ vdd gnd FILL
X_10192_ _10192_/A _10192_/B _10192_/Y vdd gnd NAND2X1
XFILL_1__9495_ vdd gnd FILL
XFILL_1__8446_ vdd gnd FILL
X_13951_ _13951_/A _13951_/B _13951_/C _13951_/Y vdd gnd NAND3X1
XFILL_1__8377_ vdd gnd FILL
X_12902_ _12902_/A _12902_/B _12902_/C _12902_/Y vdd gnd NAND3X1
XFILL_1__7328_ vdd gnd FILL
X_13882_ _13882_/A _13882_/B _13882_/Y vdd gnd NAND2X1
X_12833_ _12833_/A _12833_/B _12833_/C _12833_/Y vdd gnd OAI21X1
XFILL_1__7259_ vdd gnd FILL
X_12764_ _12764_/A _12764_/B _12764_/C _12764_/Y vdd gnd AOI21X1
X_14503_ _14503_/D _14503_/CLK _14503_/Q vdd gnd DFFPOSX1
X_11715_ _11715_/A _11715_/B _11715_/Y vdd gnd NAND2X1
X_12695_ _12695_/A _12695_/B _12695_/Y vdd gnd NAND2X1
XFILL_2__11060_ vdd gnd FILL
XFILL_1__10810_ vdd gnd FILL
XFILL_1__11790_ vdd gnd FILL
X_14434_ _14434_/A _14434_/B _14434_/Y vdd gnd NOR2X1
X_11646_ _11646_/D _11646_/CLK _11646_/Q vdd gnd DFFPOSX1
XFILL_0__12170_ vdd gnd FILL
X_14365_ _14365_/A _14365_/B _14365_/Y vdd gnd OR2X2
X_11577_ _11577_/A _11577_/B _11577_/C _11577_/Y vdd gnd OAI21X1
XFILL_0__11121_ vdd gnd FILL
XFILL_1__10672_ vdd gnd FILL
X_13316_ _13316_/A _13316_/Y vdd gnd INVX1
X_10528_ _10528_/A _10528_/B _10528_/Y vdd gnd NAND2X1
X_14296_ _14296_/A _14296_/B _14296_/Y vdd gnd NAND2X1
XFILL_2__8624_ vdd gnd FILL
XFILL_1__12411_ vdd gnd FILL
XFILL_0__11052_ vdd gnd FILL
XFILL_2_CLKBUF1_insert46 vdd gnd FILL
XFILL_2__11962_ vdd gnd FILL
XFILL_1__13391_ vdd gnd FILL
X_13247_ _13247_/A _13247_/B _13247_/Y vdd gnd NAND2X1
X_10459_ _10459_/A _10459_/Y vdd gnd INVX1
XFILL_2__13701_ vdd gnd FILL
XFILL_2_CLKBUF1_insert79 vdd gnd FILL
XFILL_0__10003_ vdd gnd FILL
XFILL_2__8555_ vdd gnd FILL
XFILL_1__12342_ vdd gnd FILL
XFILL_2__11893_ vdd gnd FILL
X_13178_ _13178_/A _13178_/B _13178_/Y vdd gnd NOR2X1
XFILL_0__7570_ vdd gnd FILL
XFILL_2__13632_ vdd gnd FILL
XFILL_0__14811_ vdd gnd FILL
XFILL_2__8486_ vdd gnd FILL
XFILL_1__12273_ vdd gnd FILL
X_12129_ _12129_/A _12129_/Y vdd gnd INVX1
XFILL_1__14012_ vdd gnd FILL
XFILL_1__11224_ vdd gnd FILL
XFILL_2__13563_ vdd gnd FILL
XFILL_0__14742_ vdd gnd FILL
XFILL_0__9240_ vdd gnd FILL
XFILL_0__11954_ vdd gnd FILL
XFILL_0_CLKBUF1_insert50 vdd gnd FILL
XFILL256350x57750 vdd gnd FILL
XFILL_0_CLKBUF1_insert61 vdd gnd FILL
XFILL_0_BUFX2_insert17 vdd gnd FILL
XFILL_0_BUFX2_insert28 vdd gnd FILL
XFILL_0__10905_ vdd gnd FILL
XFILL_1__11155_ vdd gnd FILL
XFILL_0__14673_ vdd gnd FILL
XFILL_0_CLKBUF1_insert72 vdd gnd FILL
XFILL_0__9171_ vdd gnd FILL
XFILL_0_CLKBUF1_insert83 vdd gnd FILL
XFILL_0__11885_ vdd gnd FILL
XFILL_2__9107_ vdd gnd FILL
XFILL_0_CLKBUF1_insert94 vdd gnd FILL
XFILL_1__10106_ vdd gnd FILL
XFILL_0__13624_ vdd gnd FILL
XFILL_1__11086_ vdd gnd FILL
XFILL_0__8122_ vdd gnd FILL
XFILL_0__10836_ vdd gnd FILL
XFILL_2__9038_ vdd gnd FILL
X_8750_ _8750_/A _8750_/B _8750_/Y vdd gnd AND2X2
XFILL_1__10037_ vdd gnd FILL
XFILL_1__14914_ vdd gnd FILL
XFILL_0__13555_ vdd gnd FILL
X_7701_ _7701_/A _7701_/B _7701_/Y vdd gnd OR2X2
XFILL_0__8053_ vdd gnd FILL
X_8681_ _8681_/A _8681_/Y vdd gnd INVX1
XFILL_2__11327_ vdd gnd FILL
XFILL_1__14845_ vdd gnd FILL
XFILL_0__12506_ vdd gnd FILL
X_7632_ _7632_/A _7632_/B _7632_/Y vdd gnd NAND2X1
XFILL_2__11258_ vdd gnd FILL
XFILL_1__14776_ vdd gnd FILL
XFILL_0__12437_ vdd gnd FILL
XFILL_1__11988_ vdd gnd FILL
X_7563_ _7563_/A _7563_/B _7563_/Y vdd gnd NAND2X1
XFILL_1__13727_ vdd gnd FILL
XFILL_1__10939_ vdd gnd FILL
XFILL_2__11189_ vdd gnd FILL
X_9302_ _9302_/A _9302_/B _9302_/C _9302_/Y vdd gnd OAI21X1
XFILL_0__12368_ vdd gnd FILL
XFILL_0__8955_ vdd gnd FILL
X_7494_ _7494_/A _7494_/B _7494_/Y vdd gnd NAND2X1
XFILL_0__14107_ vdd gnd FILL
XFILL_1__13658_ vdd gnd FILL
XFILL_0__11319_ vdd gnd FILL
X_9233_ _9233_/A _9233_/B _9233_/C _9233_/Y vdd gnd NAND3X1
XFILL_0__7906_ vdd gnd FILL
XFILL_0__12299_ vdd gnd FILL
XFILL_0__14038_ vdd gnd FILL
XFILL_1__13589_ vdd gnd FILL
XFILL_0__7837_ vdd gnd FILL
X_9164_ _9164_/A _9164_/B _9164_/C _9164_/Y vdd gnd OAI21X1
X_8115_ _8115_/A _8115_/B _8115_/S _8115_/Y vdd gnd MUX2X1
XFILL_0__7768_ vdd gnd FILL
X_9095_ _9095_/A _9095_/Y vdd gnd INVX1
XFILL_1__8300_ vdd gnd FILL
XFILL_0__9507_ vdd gnd FILL
XFILL_1__9280_ vdd gnd FILL
X_8046_ _8046_/A _8046_/B _8046_/Y vdd gnd NAND2X1
XFILL_0__7699_ vdd gnd FILL
XFILL_0__9438_ vdd gnd FILL
XFILL_1__8231_ vdd gnd FILL
XFILL_0__9369_ vdd gnd FILL
XFILL_1__8162_ vdd gnd FILL
X_9997_ _9997_/A _9997_/Y vdd gnd INVX1
XFILL_1__7113_ vdd gnd FILL
X_8948_ _8948_/A _8948_/B _8948_/Y vdd gnd NAND2X1
XFILL_1__8093_ vdd gnd FILL
X_8879_ _8879_/D _8879_/CLK _8879_/Q vdd gnd DFFPOSX1
X_11500_ _11500_/A _11500_/B _11500_/C _11500_/Y vdd gnd NAND3X1
X_12480_ _12480_/A _12480_/B _12480_/Y vdd gnd NAND2X1
XFILL_1__8995_ vdd gnd FILL
X_11431_ _11431_/A _11431_/B _11431_/Y vdd gnd NOR2X1
X_14150_ _14150_/A _14150_/B _14150_/C _14150_/Y vdd gnd OAI21X1
X_11362_ _11362_/A _11362_/B _11362_/C _11362_/Y vdd gnd NAND3X1
XFILL_1__7877_ vdd gnd FILL
X_13101_ _13101_/A _13101_/B _13101_/C _13101_/Y vdd gnd AOI21X1
X_10313_ _10313_/A _10313_/B _10313_/C _10313_/Y vdd gnd OAI21X1
X_14081_ _14081_/A _14081_/B _14081_/Y vdd gnd AND2X2
XFILL_1__9616_ vdd gnd FILL
X_11293_ _11293_/A _11293_/B _11293_/Y vdd gnd NAND2X1
X_13032_ _13032_/A _13032_/B _13032_/C _13032_/Y vdd gnd AOI21X1
X_10244_ _10244_/A _10244_/B _10244_/C _10244_/Y vdd gnd OAI21X1
XFILL_1__9547_ vdd gnd FILL
X_10175_ _10175_/A _10175_/Y vdd gnd INVX1
XFILL_1__9478_ vdd gnd FILL
XFILL_2__7222_ vdd gnd FILL
XFILL_1__8429_ vdd gnd FILL
X_13934_ _13934_/A _13934_/B _13934_/C _13934_/Y vdd gnd OAI21X1
XFILL_2__7153_ vdd gnd FILL
X_13865_ _13865_/A _13865_/B _13865_/Y vdd gnd NAND2X1
XFILL_2__7084_ vdd gnd FILL
XFILL_0__10621_ vdd gnd FILL
XFILL_1__12960_ vdd gnd FILL
XFILL_1_BUFX2_insert320 vdd gnd FILL
X_12816_ _12816_/A _12816_/B _12816_/C _12816_/Y vdd gnd OAI21X1
XFILL_1_BUFX2_insert331 vdd gnd FILL
XFILL_1_BUFX2_insert342 vdd gnd FILL
XFILL_1__11911_ vdd gnd FILL
X_13796_ _13796_/A _13796_/B _13796_/C _13796_/Y vdd gnd NAND3X1
XFILL_0__13340_ vdd gnd FILL
XFILL_1_BUFX2_insert353 vdd gnd FILL
XFILL_0__10552_ vdd gnd FILL
XFILL_1_BUFX2_insert364 vdd gnd FILL
XFILL_1__12891_ vdd gnd FILL
XFILL_1_BUFX2_insert375 vdd gnd FILL
X_12747_ _12747_/A _12747_/B _12747_/S _12747_/Y vdd gnd MUX2X1
XFILL_1__14630_ vdd gnd FILL
XFILL_1__11842_ vdd gnd FILL
XFILL_0__10483_ vdd gnd FILL
XFILL_0__13271_ vdd gnd FILL
X_12678_ _12678_/A _12678_/Y vdd gnd INVX1
XFILL256950x36150 vdd gnd FILL
XFILL_2__11043_ vdd gnd FILL
XFILL_1__14561_ vdd gnd FILL
XFILL_0__12222_ vdd gnd FILL
XFILL_1__11773_ vdd gnd FILL
X_14417_ _14417_/A _14417_/B _14417_/Y vdd gnd NAND2X1
X_11629_ _11629_/D _11629_/CLK _11629_/Q vdd gnd DFFPOSX1
XFILL_1__13512_ vdd gnd FILL
XFILL_1__14492_ vdd gnd FILL
XFILL_0__12153_ vdd gnd FILL
XFILL_0__8740_ vdd gnd FILL
X_14348_ _14348_/A _14348_/B _14348_/Y vdd gnd NAND2X1
XFILL_0__11104_ vdd gnd FILL
XFILL_1__10655_ vdd gnd FILL
XFILL_0__12084_ vdd gnd FILL
X_14279_ _14279_/A _14279_/B _14279_/C _14279_/Y vdd gnd NAND3X1
XFILL_0__8671_ vdd gnd FILL
XFILL256950x208950 vdd gnd FILL
XFILL_0__11035_ vdd gnd FILL
XFILL_1__13374_ vdd gnd FILL
XFILL_0__7622_ vdd gnd FILL
XFILL_1__10586_ vdd gnd FILL
XFILL_1__12325_ vdd gnd FILL
XFILL_0__7553_ vdd gnd FILL
XFILL_2__13615_ vdd gnd FILL
XFILL_2__10827_ vdd gnd FILL
XFILL_1__12256_ vdd gnd FILL
XFILL_0__12986_ vdd gnd FILL
X_9920_ _9920_/A _9920_/B _9920_/S _9920_/Y vdd gnd MUX2X1
XFILL_0__7484_ vdd gnd FILL
XFILL_1__11207_ vdd gnd FILL
XFILL_2__13546_ vdd gnd FILL
XFILL_0__14725_ vdd gnd FILL
XFILL_0__9223_ vdd gnd FILL
XFILL_0__11937_ vdd gnd FILL
XFILL_1__12187_ vdd gnd FILL
X_9851_ _9851_/A _9851_/B _9851_/C _9851_/Y vdd gnd OAI21X1
XFILL_1__11138_ vdd gnd FILL
XFILL_0__14656_ vdd gnd FILL
XFILL_0__9154_ vdd gnd FILL
XFILL_0__11868_ vdd gnd FILL
X_8802_ _8802_/A _8802_/B _8802_/Y vdd gnd NAND2X1
X_9782_ _9782_/D _9782_/CLK _9782_/Q vdd gnd DFFPOSX1
XFILL_0__13607_ vdd gnd FILL
XFILL_1__11069_ vdd gnd FILL
XFILL_0__8105_ vdd gnd FILL
XFILL_0__10819_ vdd gnd FILL
XFILL_0__14587_ vdd gnd FILL
XFILL_0__9085_ vdd gnd FILL
X_8733_ _8733_/A _8733_/B _8733_/C _8733_/Y vdd gnd OAI21X1
XFILL_0__11799_ vdd gnd FILL
XFILL_0__13538_ vdd gnd FILL
XFILL_0__8036_ vdd gnd FILL
X_8664_ _8664_/A _8664_/B _8664_/C _8664_/Y vdd gnd OAI21X1
XFILL_1__14828_ vdd gnd FILL
X_7615_ _7615_/A _7615_/B _7615_/Y vdd gnd NOR2X1
X_8595_ _8595_/A _8595_/B _8595_/Y vdd gnd AND2X2
XFILL_1__14759_ vdd gnd FILL
XFILL_1__7800_ vdd gnd FILL
X_7546_ _7546_/A _7546_/B _7546_/Y vdd gnd NAND2X1
XFILL_1__8780_ vdd gnd FILL
XFILL_0__9987_ vdd gnd FILL
XFILL_1__7731_ vdd gnd FILL
XFILL_0__8938_ vdd gnd FILL
X_7477_ _7477_/A _7477_/B _7477_/C _7477_/Y vdd gnd AOI21X1
X_9216_ _9216_/A _9216_/B _9216_/C _9216_/Y vdd gnd AOI21X1
XFILL_1__7662_ vdd gnd FILL
XFILL_1__9401_ vdd gnd FILL
X_9147_ _9147_/A _9147_/Y vdd gnd INVX1
XFILL_1__7593_ vdd gnd FILL
XFILL_1__9332_ vdd gnd FILL
X_9078_ _9078_/A _9078_/B _9078_/C _9078_/Y vdd gnd OAI21X1
XFILL_1__9263_ vdd gnd FILL
X_8029_ _8029_/A _8029_/Y vdd gnd INVX1
XFILL_1__8214_ vdd gnd FILL
X_11980_ _11980_/A _11980_/Y vdd gnd INVX1
XFILL_1__9194_ vdd gnd FILL
X_10931_ _10931_/A _10931_/Y vdd gnd INVX1
XFILL_1__8145_ vdd gnd FILL
XFILL_0_BUFX2_insert9 vdd gnd FILL
X_10862_ _10862_/A _10862_/B _10862_/C _10862_/Y vdd gnd NAND3X1
X_13650_ _13650_/A _13650_/B _13650_/C _13650_/Y vdd gnd NAND3X1
XFILL_1__8076_ vdd gnd FILL
X_12601_ _12601_/D _12601_/CLK _12601_/Q vdd gnd DFFPOSX1
X_13581_ _13581_/A _13581_/B _13581_/C _13581_/Y vdd gnd NAND3X1
X_10793_ _10793_/A _10793_/B _10793_/C _10793_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert305 vdd gnd FILL
XFILL_0_BUFX2_insert316 vdd gnd FILL
X_12532_ _12532_/A _12532_/B _12532_/Y vdd gnd NAND2X1
XFILL_0_BUFX2_insert327 vdd gnd FILL
XFILL_0_BUFX2_insert338 vdd gnd FILL
XFILL_0_BUFX2_insert349 vdd gnd FILL
X_12463_ _12463_/A _12463_/Y vdd gnd INVX1
XFILL_1__8978_ vdd gnd FILL
X_14202_ _14202_/D _14202_/CLK _14202_/Q vdd gnd DFFPOSX1
X_11414_ _11414_/A _11414_/B _11414_/Y vdd gnd NAND2X1
XFILL_2__9510_ vdd gnd FILL
X_12394_ _12394_/A _12394_/B _12394_/Y vdd gnd OR2X2
X_14133_ _14133_/A _14133_/B _14133_/Y vdd gnd NAND2X1
X_11345_ _11345_/A _11345_/B _11345_/Y vdd gnd NAND2X1
XFILL_2__9441_ vdd gnd FILL
XFILL_1__10440_ vdd gnd FILL
X_14064_ _14064_/A _14064_/B _14064_/Y vdd gnd NAND2X1
X_11276_ _11276_/A _11276_/B _11276_/C _11276_/Y vdd gnd OAI21X1
XFILL_2__9372_ vdd gnd FILL
XFILL_1__10371_ vdd gnd FILL
X_13015_ _13015_/A _13015_/Y vdd gnd INVX1
X_10227_ _10227_/A _10227_/B _10227_/C _10227_/Y vdd gnd OAI21X1
XFILL_1__12110_ vdd gnd FILL
XFILL_1__13090_ vdd gnd FILL
XFILL_0__12840_ vdd gnd FILL
X_10158_ _10158_/A _10158_/B _10158_/C _10158_/Y vdd gnd NAND3X1
XFILL_2__14380_ vdd gnd FILL
XFILL_1__12041_ vdd gnd FILL
XFILL_2__11592_ vdd gnd FILL
XFILL_0__12771_ vdd gnd FILL
XFILL_2__7205_ vdd gnd FILL
X_10089_ _10089_/A _10089_/B _10089_/Y vdd gnd NAND2X1
XFILL_0__11722_ vdd gnd FILL
X_13917_ _13917_/A _13917_/B _13917_/Y vdd gnd NOR2X1
XFILL_2__7136_ vdd gnd FILL
X_14897_ _14897_/D _14897_/CLK _14897_/Q vdd gnd DFFPOSX1
XFILL_2__13262_ vdd gnd FILL
XFILL_0__14441_ vdd gnd FILL
XFILL_1__13992_ vdd gnd FILL
XFILL_2__12213_ vdd gnd FILL
X_13848_ _13848_/A _13848_/B _13848_/Y vdd gnd NAND2X1
XFILL_2__13193_ vdd gnd FILL
XFILL_1__12943_ vdd gnd FILL
XFILL_0__10604_ vdd gnd FILL
XFILL_0__14372_ vdd gnd FILL
XFILL_1_BUFX2_insert150 vdd gnd FILL
XFILL_0__11584_ vdd gnd FILL
XFILL_1_BUFX2_insert161 vdd gnd FILL
XFILL_1_BUFX2_insert172 vdd gnd FILL
X_13779_ _13779_/A _13779_/B _13779_/C _13779_/Y vdd gnd NAND3X1
XFILL_1_BUFX2_insert183 vdd gnd FILL
XFILL_0__13323_ vdd gnd FILL
XFILL_0__10535_ vdd gnd FILL
XFILL_1__12874_ vdd gnd FILL
XFILL_0__9910_ vdd gnd FILL
XFILL_1_BUFX2_insert194 vdd gnd FILL
XFILL_1__14613_ vdd gnd FILL
XFILL_1__11825_ vdd gnd FILL
XFILL_0__13254_ vdd gnd FILL
X_7400_ _7400_/A _7400_/B _7400_/Y vdd gnd NAND2X1
XFILL_0__10466_ vdd gnd FILL
X_8380_ _8380_/A _8380_/B _8380_/C _8380_/Y vdd gnd OAI21X1
XFILL_0__12205_ vdd gnd FILL
XFILL_1__11756_ vdd gnd FILL
XFILL_0__13185_ vdd gnd FILL
XFILL_0__10397_ vdd gnd FILL
X_7331_ _7331_/A _7331_/B _7331_/Y vdd gnd NOR2X1
XFILL_2__9708_ vdd gnd FILL
XFILL_0__12136_ vdd gnd FILL
XFILL_1__14475_ vdd gnd FILL
XFILL_0__8723_ vdd gnd FILL
X_7262_ _7262_/A _7262_/B _7262_/Y vdd gnd NAND2X1
XFILL_2__9639_ vdd gnd FILL
XFILL_1__13426_ vdd gnd FILL
XFILL_1__10638_ vdd gnd FILL
X_9001_ _9001_/A _9001_/B _9001_/C _9001_/Y vdd gnd OAI21X1
XFILL_0__12067_ vdd gnd FILL
XFILL_2__12977_ vdd gnd FILL
XFILL_0__8654_ vdd gnd FILL
X_7193_ _7193_/A _7193_/B _7193_/S _7193_/Y vdd gnd MUX2X1
XFILL_0__11018_ vdd gnd FILL
XFILL_1__13357_ vdd gnd FILL
XFILL_1__10569_ vdd gnd FILL
XFILL_0__7605_ vdd gnd FILL
XFILL_0__8585_ vdd gnd FILL
XFILL_1__12308_ vdd gnd FILL
XFILL_1__13288_ vdd gnd FILL
XFILL_0__7536_ vdd gnd FILL
XFILL_1__12239_ vdd gnd FILL
XFILL_0__12969_ vdd gnd FILL
XFILL_0__7467_ vdd gnd FILL
X_9903_ _9903_/A _9903_/Y vdd gnd INVX1
XFILL_0__14708_ vdd gnd FILL
XFILL_0__9206_ vdd gnd FILL
X_9834_ _9834_/D _9834_/CLK _9834_/Q vdd gnd DFFPOSX1
XFILL_0__7398_ vdd gnd FILL
XFILL_0__14639_ vdd gnd FILL
XFILL_0__9137_ vdd gnd FILL
X_9765_ _9765_/D _9765_/CLK _9765_/Q vdd gnd DFFPOSX1
XFILL_0__9068_ vdd gnd FILL
X_8716_ _8716_/A _8716_/B _8716_/C _8716_/Y vdd gnd AOI21X1
XFILL_1__9950_ vdd gnd FILL
X_9696_ _9696_/A _9696_/B _9696_/C _9696_/Y vdd gnd OAI21X1
XFILL_0__8019_ vdd gnd FILL
X_8647_ _8647_/A _8647_/Y vdd gnd INVX1
XFILL_1__9881_ vdd gnd FILL
XFILL_1__8832_ vdd gnd FILL
X_8578_ _8578_/A _8578_/Y vdd gnd INVX1
X_7529_ _7529_/A _7529_/B _7529_/C _7529_/Y vdd gnd AOI21X1
XFILL_1__8763_ vdd gnd FILL
XFILL_1__7714_ vdd gnd FILL
XFILL_1__8694_ vdd gnd FILL
X_11130_ _11130_/A _11130_/B _11130_/Y vdd gnd NAND2X1
XFILL_1__7645_ vdd gnd FILL
X_11061_ _11061_/A _11061_/B _11061_/C _11061_/Y vdd gnd NAND3X1
XFILL_1__7576_ vdd gnd FILL
X_10012_ _10012_/A _10012_/B _10012_/Y vdd gnd NAND2X1
XFILL_1__9315_ vdd gnd FILL
X_14820_ _14820_/A _14820_/Y vdd gnd INVX1
XFILL_1__9246_ vdd gnd FILL
X_14751_ _14751_/A _14751_/B _14751_/Y vdd gnd NAND2X1
XFILL_1__9177_ vdd gnd FILL
X_11963_ _11963_/A _11963_/Y vdd gnd INVX1
X_13702_ _13702_/A _13702_/B _13702_/C _13702_/Y vdd gnd NOR3X1
XFILL_1__8128_ vdd gnd FILL
X_10914_ _10914_/A _10914_/B _10914_/C _10914_/Y vdd gnd OAI21X1
X_14682_ _14682_/A _14682_/B _14682_/Y vdd gnd NOR2X1
X_11894_ _11894_/A _11894_/B _11894_/C _11894_/Y vdd gnd OAI21X1
XFILL_2__9990_ vdd gnd FILL
X_13633_ _13633_/A _13633_/B _13633_/Y vdd gnd NAND2X1
X_10845_ _10845_/A _10845_/B _10845_/Y vdd gnd NOR2X1
XFILL_1__8059_ vdd gnd FILL
X_13564_ _13564_/A _13564_/B _13564_/Y vdd gnd NAND2X1
X_10776_ _10776_/A _10776_/Y vdd gnd INVX2
XFILL_0_BUFX2_insert113 vdd gnd FILL
XFILL_0_BUFX2_insert124 vdd gnd FILL
XFILL_0_BUFX2_insert135 vdd gnd FILL
XFILL_0__10320_ vdd gnd FILL
XFILL_0_BUFX2_insert146 vdd gnd FILL
X_12515_ _12515_/A _12515_/B _12515_/C _12515_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert157 vdd gnd FILL
X_13495_ _13495_/D _13495_/CLK _13495_/Q vdd gnd DFFPOSX1
XFILL_0_BUFX2_insert168 vdd gnd FILL
XFILL_1__11610_ vdd gnd FILL
XFILL_0_BUFX2_insert179 vdd gnd FILL
XFILL_0__10251_ vdd gnd FILL
X_12446_ _12446_/A _12446_/B _12446_/Y vdd gnd AND2X2
XFILL_2__12900_ vdd gnd FILL
XFILL_1__11541_ vdd gnd FILL
XFILL_0__10182_ vdd gnd FILL
XFILL_2__13880_ vdd gnd FILL
X_12377_ _12377_/A _12377_/Y vdd gnd INVX1
XFILL_1__14260_ vdd gnd FILL
XFILL_2__12831_ vdd gnd FILL
XFILL_1__11472_ vdd gnd FILL
X_14116_ _14116_/A _14116_/B _14116_/Y vdd gnd NAND2X1
X_11328_ _11328_/A _11328_/B _11328_/Y vdd gnd NAND2X1
XFILL_1__13211_ vdd gnd FILL
XFILL_2__9424_ vdd gnd FILL
XFILL_1__10423_ vdd gnd FILL
XFILL_2__12762_ vdd gnd FILL
XFILL_0__13941_ vdd gnd FILL
X_14047_ _14047_/A _14047_/B _14047_/C _14047_/Y vdd gnd AOI21X1
X_11259_ _11259_/A _11259_/B _11259_/Y vdd gnd NAND2X1
XFILL_1__13142_ vdd gnd FILL
XFILL_2__9355_ vdd gnd FILL
XFILL_1__10354_ vdd gnd FILL
XFILL_2__12693_ vdd gnd FILL
XFILL_0__13872_ vdd gnd FILL
XFILL_0__8370_ vdd gnd FILL
XFILL_1__13073_ vdd gnd FILL
XFILL_2__9286_ vdd gnd FILL
XFILL_0__12823_ vdd gnd FILL
XFILL_0__7321_ vdd gnd FILL
XFILL_1__10285_ vdd gnd FILL
XFILL_1__12024_ vdd gnd FILL
XFILL_2__14363_ vdd gnd FILL
XFILL_2__11575_ vdd gnd FILL
XFILL_0__12754_ vdd gnd FILL
XFILL_0__7252_ vdd gnd FILL
X_7880_ _7880_/A _7880_/B _7880_/Y vdd gnd NAND2X1
XFILL_2__14294_ vdd gnd FILL
XFILL_0__11705_ vdd gnd FILL
XFILL_0__12685_ vdd gnd FILL
XFILL_0__7183_ vdd gnd FILL
XFILL_2__7119_ vdd gnd FILL
XFILL_0__14424_ vdd gnd FILL
XFILL_1__13975_ vdd gnd FILL
X_9550_ _9550_/A _9550_/B _9550_/C _9550_/Y vdd gnd OAI21X1
XFILL_1__12926_ vdd gnd FILL
XFILL_0__14355_ vdd gnd FILL
X_8501_ _8501_/A _8501_/B _8501_/C _8501_/Y vdd gnd NAND3X1
XFILL_0__11567_ vdd gnd FILL
X_9481_ _9481_/A _9481_/B _9481_/C _9481_/Y vdd gnd AOI21X1
XFILL_2__12127_ vdd gnd FILL
XFILL_0__13306_ vdd gnd FILL
XFILL_0__10518_ vdd gnd FILL
XFILL_1__12857_ vdd gnd FILL
XFILL_0__14286_ vdd gnd FILL
X_8432_ _8432_/A _8432_/B _8432_/C _8432_/Y vdd gnd OAI21X1
XFILL_0__11498_ vdd gnd FILL
XBUFX2_insert19 BUFX2_insert19/A BUFX2_insert19/Y vdd gnd BUFX2
XFILL_2__12058_ vdd gnd FILL
XFILL_1__11808_ vdd gnd FILL
XFILL_0__13237_ vdd gnd FILL
XFILL_0__10449_ vdd gnd FILL
XFILL_1__12788_ vdd gnd FILL
X_8363_ _8363_/A _8363_/B _8363_/Y vdd gnd NOR2X1
XFILL_1__11739_ vdd gnd FILL
XFILL_0__13168_ vdd gnd FILL
X_7314_ _7314_/A _7314_/B _7314_/C _7314_/Y vdd gnd AOI21X1
XFILL_0__9755_ vdd gnd FILL
X_8294_ _8294_/A _8294_/B _8294_/C _8294_/D _8294_/Y vdd gnd AOI22X1
XFILL_1__14458_ vdd gnd FILL
XFILL_0__12119_ vdd gnd FILL
XFILL_0__13099_ vdd gnd FILL
XFILL_0__8706_ vdd gnd FILL
X_7245_ _7245_/A _7245_/B _7245_/C _7245_/Y vdd gnd OAI21X1
XFILL_0__9686_ vdd gnd FILL
XFILL_1__13409_ vdd gnd FILL
XFILL_1__14389_ vdd gnd FILL
XFILL_1__7430_ vdd gnd FILL
XFILL_0__8637_ vdd gnd FILL
X_7176_ _7176_/A _7176_/B _7176_/Y vdd gnd NAND2X1
XFILL_1__7361_ vdd gnd FILL
XFILL_0__8568_ vdd gnd FILL
XFILL_1__9100_ vdd gnd FILL
XFILL_2_BUFX2_insert208 vdd gnd FILL
XFILL_0__7519_ vdd gnd FILL
XFILL_1__7292_ vdd gnd FILL
XFILL_0__8499_ vdd gnd FILL
XFILL_1__9031_ vdd gnd FILL
X_9817_ _9817_/D _9817_/CLK _9817_/Q vdd gnd DFFPOSX1
X_9748_ _9748_/A _9748_/B _9748_/Y vdd gnd NAND2X1
X_10630_ _10630_/A _10630_/B _10630_/C _10630_/Y vdd gnd OAI21X1
XBUFX2_insert207 BUFX2_insert207/A BUFX2_insert207/Y vdd gnd BUFX2
XBUFX2_insert218 BUFX2_insert218/A BUFX2_insert218/Y vdd gnd BUFX2
XFILL_1__9933_ vdd gnd FILL
XBUFX2_insert229 BUFX2_insert229/A BUFX2_insert229/Y vdd gnd BUFX2
X_9679_ _9679_/A _9679_/B _9679_/C _9679_/Y vdd gnd OAI21X1
X_10561_ _10561_/A _10561_/B _10561_/Y vdd gnd NAND2X1
XFILL_1__9864_ vdd gnd FILL
X_12300_ _12300_/A _12300_/B _12300_/C _12300_/Y vdd gnd AOI21X1
X_13280_ _13280_/A _13280_/B _13280_/Y vdd gnd NAND2X1
X_10492_ _10492_/A _10492_/B _10492_/C _10492_/D _10492_/Y vdd gnd OAI22X1
XFILL_1__8815_ vdd gnd FILL
X_12231_ _12231_/A _12231_/B _12231_/Y vdd gnd NAND2X1
XFILL_1__8746_ vdd gnd FILL
X_12162_ _12162_/A _12162_/B _12162_/C _12162_/Y vdd gnd NAND3X1
XFILL_2__7470_ vdd gnd FILL
XFILL_1__8677_ vdd gnd FILL
X_11113_ _11113_/A _11113_/B _11113_/C _11113_/D _11113_/Y vdd gnd AOI22X1
X_12093_ _12093_/A _12093_/B _12093_/C _12093_/Y vdd gnd NAND3X1
XFILL_1__7628_ vdd gnd FILL
X_11044_ _11044_/A _11044_/Y vdd gnd INVX1
XFILL_1__7559_ vdd gnd FILL
XFILL_2__9071_ vdd gnd FILL
XFILL_1__10070_ vdd gnd FILL
X_14803_ _14803_/A _14803_/B _14803_/C _14803_/Y vdd gnd OAI21X1
XFILL257550x86550 vdd gnd FILL
XFILL_2__8022_ vdd gnd FILL
XFILL_1__9229_ vdd gnd FILL
XFILL_2__11360_ vdd gnd FILL
X_12995_ _12995_/A _12995_/B _12995_/Y vdd gnd NOR2X1
X_14734_ _14734_/A _14734_/B _14734_/Y vdd gnd NAND2X1
XFILL_2__10311_ vdd gnd FILL
X_11946_ _11946_/A _11946_/B _11946_/C _11946_/Y vdd gnd OAI21X1
XFILL_2__11291_ vdd gnd FILL
XFILL_0__12470_ vdd gnd FILL
X_14665_ _14665_/A _14665_/B _14665_/Y vdd gnd OR2X2
X_11877_ _11877_/A _11877_/B _11877_/C _11877_/Y vdd gnd AOI21X1
XFILL_0__11421_ vdd gnd FILL
XFILL_1__13760_ vdd gnd FILL
XFILL_1__10972_ vdd gnd FILL
X_13616_ _13616_/A _13616_/B _13616_/C _13616_/Y vdd gnd AOI21X1
X_10828_ _10828_/A _10828_/Y vdd gnd INVX8
X_14596_ _14596_/A _14596_/B _14596_/Y vdd gnd AND2X2
XFILL_2__8924_ vdd gnd FILL
XFILL_1__12711_ vdd gnd FILL
XFILL_0__14140_ vdd gnd FILL
XFILL_0__11352_ vdd gnd FILL
XFILL_1__13691_ vdd gnd FILL
X_13547_ _13547_/A _13547_/Y vdd gnd INVX8
X_10759_ _10759_/D _10759_/CLK _10759_/Q vdd gnd DFFPOSX1
XFILL_1__12642_ vdd gnd FILL
XFILL_0__10303_ vdd gnd FILL
XFILL_0__14071_ vdd gnd FILL
XFILL_0__11283_ vdd gnd FILL
XFILL_0__7870_ vdd gnd FILL
XFILL_2__7806_ vdd gnd FILL
X_13478_ _13478_/D _13478_/CLK _13478_/Q vdd gnd DFFPOSX1
XFILL_2__13932_ vdd gnd FILL
XFILL_0__13022_ vdd gnd FILL
XFILL_0__10234_ vdd gnd FILL
X_12429_ _12429_/A _12429_/B _12429_/C _12429_/Y vdd gnd OAI21X1
XFILL_1__14312_ vdd gnd FILL
XFILL_2__7737_ vdd gnd FILL
XFILL_1__11524_ vdd gnd FILL
XFILL_2__13863_ vdd gnd FILL
XFILL_0__10165_ vdd gnd FILL
XFILL_0__9540_ vdd gnd FILL
XFILL_1__14243_ vdd gnd FILL
XFILL_2__12814_ vdd gnd FILL
XFILL_1__11455_ vdd gnd FILL
XFILL_0__10096_ vdd gnd FILL
XFILL_2__13794_ vdd gnd FILL
XFILL_0__9471_ vdd gnd FILL
XFILL_2__9407_ vdd gnd FILL
XFILL_1__10406_ vdd gnd FILL
XFILL_2__12745_ vdd gnd FILL
XFILL_0__13924_ vdd gnd FILL
XFILL_1__11386_ vdd gnd FILL
XFILL_0__8422_ vdd gnd FILL
XFILL_1__13125_ vdd gnd FILL
XFILL_2__9338_ vdd gnd FILL
XFILL_1__10337_ vdd gnd FILL
XFILL_0__13855_ vdd gnd FILL
XFILL_2__12676_ vdd gnd FILL
XFILL_0__8353_ vdd gnd FILL
X_8981_ _8981_/A _8981_/Y vdd gnd INVX8
XFILL_1__13056_ vdd gnd FILL
XFILL_2__9269_ vdd gnd FILL
XFILL_0__12806_ vdd gnd FILL
XFILL_1__10268_ vdd gnd FILL
XFILL_0__7304_ vdd gnd FILL
XFILL_0__13786_ vdd gnd FILL
XFILL_0__10998_ vdd gnd FILL
X_7932_ _7932_/D _7932_/CLK _7932_/Q vdd gnd DFFPOSX1
XFILL_0__8284_ vdd gnd FILL
XFILL_1__12007_ vdd gnd FILL
XFILL_2__11558_ vdd gnd FILL
XFILL_0__12737_ vdd gnd FILL
XFILL_0__7235_ vdd gnd FILL
XFILL_1__10199_ vdd gnd FILL
X_7863_ _7863_/A _7863_/B _7863_/C _7863_/Y vdd gnd OAI21X1
XFILL_2__11489_ vdd gnd FILL
XFILL_0__12668_ vdd gnd FILL
XFILL_0__7166_ vdd gnd FILL
X_9602_ _9602_/A _9602_/B _9602_/Y vdd gnd OR2X2
X_7794_ _7794_/A _7794_/B _7794_/Y vdd gnd NAND2X1
XFILL_0__14407_ vdd gnd FILL
XFILL_1__13958_ vdd gnd FILL
X_9533_ _9533_/A _9533_/B _9533_/C _9533_/Y vdd gnd OAI21X1
XFILL_0__7097_ vdd gnd FILL
XFILL_0__14338_ vdd gnd FILL
XFILL_1__12909_ vdd gnd FILL
XFILL_1__13889_ vdd gnd FILL
X_9464_ _9464_/A _9464_/Y vdd gnd INVX1
XFILL_0__14269_ vdd gnd FILL
X_8415_ _8415_/A _8415_/B _8415_/C _8415_/Y vdd gnd OAI21X1
X_9395_ _9395_/A _9395_/B _9395_/Y vdd gnd OR2X2
XFILL_1__8600_ vdd gnd FILL
X_8346_ _8346_/A _8346_/B _8346_/Y vdd gnd NAND2X1
XFILL_1__9580_ vdd gnd FILL
XFILL_0__7999_ vdd gnd FILL
XFILL_0__9738_ vdd gnd FILL
XFILL_1__8531_ vdd gnd FILL
X_8277_ _8277_/A _8277_/B _8277_/Y vdd gnd NOR2X1
X_7228_ _7228_/A _7228_/Y vdd gnd INVX2
XFILL_0__9669_ vdd gnd FILL
XFILL_1__8462_ vdd gnd FILL
XFILL_1__7413_ vdd gnd FILL
X_7159_ _7159_/A _7159_/B _7159_/Y vdd gnd NOR2X1
XFILL_1__8393_ vdd gnd FILL
XFILL_1__7344_ vdd gnd FILL
XFILL_1__7275_ vdd gnd FILL
X_11800_ _11800_/A _11800_/B _11800_/Y vdd gnd NAND2X1
XFILL_1__9014_ vdd gnd FILL
X_12780_ _12780_/A _12780_/B _12780_/Y vdd gnd NOR2X1
XFILL257550x18150 vdd gnd FILL
X_11731_ _11731_/A _11731_/B _11731_/C _11731_/Y vdd gnd OAI21X1
X_14450_ _14450_/A _14450_/B _14450_/Y vdd gnd NAND2X1
X_11662_ _11662_/D _11662_/CLK _11662_/Q vdd gnd DFFPOSX1
X_13401_ _13401_/A _13401_/B _13401_/C _13401_/Y vdd gnd OAI21X1
X_10613_ _10613_/A _10613_/B _10613_/C _10613_/Y vdd gnd OAI21X1
XFILL_1__9916_ vdd gnd FILL
X_14381_ _14381_/A _14381_/B _14381_/C _14381_/D _14381_/Y vdd gnd AOI22X1
X_11593_ _11593_/A _11593_/Y vdd gnd INVX1
X_10544_ _10544_/A _10544_/B _10544_/Y vdd gnd NAND2X1
X_13332_ _13332_/A _13332_/B _13332_/C _13332_/D _13332_/Y vdd gnd OAI22X1
XFILL_1__9847_ vdd gnd FILL
XFILL257550x61350 vdd gnd FILL
X_10475_ _10475_/A _10475_/B _10475_/Y vdd gnd NAND2X1
X_13263_ _13263_/A _13263_/B _13263_/C _13263_/Y vdd gnd AOI21X1
X_12214_ _12214_/A _12214_/B _12214_/C _12214_/Y vdd gnd OAI21X1
X_13194_ _13194_/A _13194_/B _13194_/Y vdd gnd NOR2X1
XFILL_2__7522_ vdd gnd FILL
XFILL_1__8729_ vdd gnd FILL
XFILL_2__10860_ vdd gnd FILL
X_12145_ _12145_/A _12145_/B _12145_/Y vdd gnd OR2X2
XFILL_2__7453_ vdd gnd FILL
XFILL_1__11240_ vdd gnd FILL
XFILL_2__10791_ vdd gnd FILL
XFILL_0__11970_ vdd gnd FILL
X_12076_ _12076_/A _12076_/B _12076_/C _12076_/Y vdd gnd OAI21X1
XFILL_2__7384_ vdd gnd FILL
XFILL_2__12530_ vdd gnd FILL
XFILL_1__11171_ vdd gnd FILL
XFILL_0__10921_ vdd gnd FILL
X_11027_ _11027_/A _11027_/B _11027_/Y vdd gnd NOR2X1
XFILL_1__10122_ vdd gnd FILL
XFILL_0__13640_ vdd gnd FILL
XFILL_0__10852_ vdd gnd FILL
XFILL_1__10053_ vdd gnd FILL
XFILL_0__13571_ vdd gnd FILL
XFILL_0__10783_ vdd gnd FILL
XFILL_2__8005_ vdd gnd FILL
X_12978_ _12978_/A _12978_/B _12978_/C _12978_/D _12978_/Y vdd gnd AOI22X1
XFILL_0__12522_ vdd gnd FILL
XFILL_1__14861_ vdd gnd FILL
X_14717_ _14717_/A _14717_/B _14717_/Y vdd gnd NOR2X1
X_11929_ _11929_/A _11929_/B _11929_/C _11929_/Y vdd gnd NAND3X1
XFILL_1__13812_ vdd gnd FILL
XFILL_0__12453_ vdd gnd FILL
XFILL_1__14792_ vdd gnd FILL
X_14648_ _14648_/A _14648_/B _14648_/C _14648_/Y vdd gnd AOI21X1
XFILL_2__10225_ vdd gnd FILL
XFILL_0__11404_ vdd gnd FILL
XFILL_1__10955_ vdd gnd FILL
XFILL_1__13743_ vdd gnd FILL
XFILL_0__12384_ vdd gnd FILL
XFILL_0__8971_ vdd gnd FILL
X_14579_ _14579_/A _14579_/B _14579_/C _14579_/Y vdd gnd OAI21X1
XFILL_2__10156_ vdd gnd FILL
XFILL_0__14123_ vdd gnd FILL
XFILL_0__11335_ vdd gnd FILL
XFILL_1__13674_ vdd gnd FILL
XFILL256650x219750 vdd gnd FILL
XFILL_1__10886_ vdd gnd FILL
XFILL_1__12625_ vdd gnd FILL
XFILL_2__10087_ vdd gnd FILL
XFILL_0__14054_ vdd gnd FILL
X_8200_ _8200_/A _8200_/B _8200_/C _8200_/Y vdd gnd AOI21X1
XFILL_0__11266_ vdd gnd FILL
XFILL_0__7853_ vdd gnd FILL
X_9180_ _9180_/A _9180_/Y vdd gnd INVX1
XFILL_0__13005_ vdd gnd FILL
XFILL_0__10217_ vdd gnd FILL
X_8131_ _8131_/A _8131_/B _8131_/Y vdd gnd NAND2X1
XFILL_0__11197_ vdd gnd FILL
XFILL_0__7784_ vdd gnd FILL
XFILL_1__11507_ vdd gnd FILL
XFILL_2__13846_ vdd gnd FILL
XFILL_0__10148_ vdd gnd FILL
XFILL_1__12487_ vdd gnd FILL
XFILL_0__9523_ vdd gnd FILL
X_8062_ _8062_/A _8062_/B _8062_/Y vdd gnd NAND2X1
XFILL_1__14226_ vdd gnd FILL
XFILL_1__11438_ vdd gnd FILL
XFILL_2__13777_ vdd gnd FILL
XFILL_2__10989_ vdd gnd FILL
XFILL_0__10079_ vdd gnd FILL
XFILL_0__9454_ vdd gnd FILL
XFILL_1__14157_ vdd gnd FILL
XFILL_0__13907_ vdd gnd FILL
XFILL_1__11369_ vdd gnd FILL
XFILL_0__8405_ vdd gnd FILL
XFILL_1__13108_ vdd gnd FILL
XFILL_0__9385_ vdd gnd FILL
XFILL_1__14088_ vdd gnd FILL
XFILL_0__13838_ vdd gnd FILL
XFILL_0__8336_ vdd gnd FILL
X_8964_ _8964_/A _8964_/B _8964_/C _8964_/Y vdd gnd AOI21X1
XFILL_1__13039_ vdd gnd FILL
XFILL_0__13769_ vdd gnd FILL
X_7915_ _7915_/A _7915_/B _7915_/C _7915_/Y vdd gnd OAI21X1
XFILL_0__8267_ vdd gnd FILL
X_8895_ _8895_/D _8895_/CLK _8895_/Q vdd gnd DFFPOSX1
XFILL_0__7218_ vdd gnd FILL
X_7846_ _7846_/A _7846_/B _7846_/Y vdd gnd NAND2X1
XFILL_0__8198_ vdd gnd FILL
XFILL_0_CLKBUF1_insert105 vdd gnd FILL
XFILL_0__7149_ vdd gnd FILL
X_7777_ _7777_/A _7777_/B _7777_/Y vdd gnd NOR2X1
X_9516_ _9516_/A _9516_/B _9516_/Y vdd gnd NOR2X1
XFILL_1__9701_ vdd gnd FILL
X_9447_ _9447_/A _9447_/Y vdd gnd INVX1
XFILL_1__7893_ vdd gnd FILL
XFILL_1__9632_ vdd gnd FILL
X_9378_ _9378_/A _9378_/B _9378_/Y vdd gnd NAND2X1
X_10260_ _10260_/A _10260_/B _10260_/Y vdd gnd NAND2X1
X_8329_ _8329_/A _8329_/B _8329_/Y vdd gnd NAND2X1
XFILL_1__9563_ vdd gnd FILL
X_10191_ _10191_/A _10191_/Y vdd gnd INVX1
XFILL_1__8514_ vdd gnd FILL
XFILL_1__9494_ vdd gnd FILL
XFILL_1__8445_ vdd gnd FILL
X_13950_ _13950_/A _13950_/Y vdd gnd INVX1
XFILL_1__8376_ vdd gnd FILL
X_12901_ _12901_/A _12901_/B _12901_/C _12901_/Y vdd gnd OAI21X1
X_13881_ _13881_/A _13881_/Y vdd gnd INVX1
XFILL_1__7327_ vdd gnd FILL
X_12832_ _12832_/A _12832_/B _12832_/Y vdd gnd AND2X2
XFILL_1__7258_ vdd gnd FILL
X_12763_ _12763_/A _12763_/B _12763_/C _12763_/Y vdd gnd OAI21X1
XFILL_1__7189_ vdd gnd FILL
X_14502_ _14502_/D _14502_/CLK _14502_/Q vdd gnd DFFPOSX1
X_11714_ _11714_/A _11714_/B _11714_/C _11714_/D _11714_/Y vdd gnd AOI22X1
X_12694_ _12694_/A _12694_/Y vdd gnd INVX8
X_14433_ _14433_/A _14433_/Y vdd gnd INVX2
XFILL_2__10010_ vdd gnd FILL
X_11645_ _11645_/D _11645_/CLK _11645_/Q vdd gnd DFFPOSX1
XFILL_2__9741_ vdd gnd FILL
X_14364_ _14364_/A _14364_/B _14364_/Y vdd gnd NAND2X1
X_11576_ _11576_/A _11576_/B _11576_/Y vdd gnd NAND2X1
XFILL_2__9672_ vdd gnd FILL
XFILL_0__11120_ vdd gnd FILL
XFILL_1__10671_ vdd gnd FILL
X_13315_ _13315_/A _13315_/B _13315_/Y vdd gnd NOR2X1
X_10527_ _10527_/A _10527_/B _10527_/Y vdd gnd NAND2X1
X_14295_ _14295_/A _14295_/Y vdd gnd INVX1
XFILL_1__12410_ vdd gnd FILL
XFILL_0__11051_ vdd gnd FILL
XFILL_2_CLKBUF1_insert36 vdd gnd FILL
XFILL_1__13390_ vdd gnd FILL
X_10458_ _10458_/A _10458_/B _10458_/C _10458_/Y vdd gnd OAI21X1
XFILL_2_CLKBUF1_insert58 vdd gnd FILL
X_13246_ _13246_/A _13246_/B _13246_/Y vdd gnd OR2X2
XFILL_0__10002_ vdd gnd FILL
XFILL_1__12341_ vdd gnd FILL
XFILL_2__10912_ vdd gnd FILL
X_13177_ _13177_/A _13177_/B _13177_/Y vdd gnd NOR2X1
X_10389_ _10389_/A _10389_/B _10389_/C _10389_/Y vdd gnd AOI21X1
XFILL_2__7505_ vdd gnd FILL
XFILL_0__14810_ vdd gnd FILL
XFILL_1__12272_ vdd gnd FILL
XFILL_2__10843_ vdd gnd FILL
X_12128_ _12128_/A _12128_/B _12128_/C _12128_/Y vdd gnd OAI21X1
XFILL_1__14011_ vdd gnd FILL
XFILL_2__7436_ vdd gnd FILL
XFILL_1__11223_ vdd gnd FILL
XFILL_0__14741_ vdd gnd FILL
XFILL_2__10774_ vdd gnd FILL
XFILL_0__11953_ vdd gnd FILL
X_12059_ _12059_/A _12059_/B _12059_/Y vdd gnd NOR2X1
XFILL_0_CLKBUF1_insert40 vdd gnd FILL
XFILL_2__12513_ vdd gnd FILL
XFILL_2__7367_ vdd gnd FILL
XFILL_0_BUFX2_insert18 vdd gnd FILL
XFILL_0_CLKBUF1_insert51 vdd gnd FILL
XFILL_1__11154_ vdd gnd FILL
XFILL_0__10904_ vdd gnd FILL
XFILL_0__14672_ vdd gnd FILL
XFILL_0_CLKBUF1_insert62 vdd gnd FILL
XFILL_0_CLKBUF1_insert73 vdd gnd FILL
XFILL_0__9170_ vdd gnd FILL
XFILL_0__11884_ vdd gnd FILL
XFILL_0_CLKBUF1_insert84 vdd gnd FILL
XFILL_1__10105_ vdd gnd FILL
XFILL_2__12444_ vdd gnd FILL
XFILL_0_CLKBUF1_insert95 vdd gnd FILL
XFILL_0__13623_ vdd gnd FILL
XFILL_1__11085_ vdd gnd FILL
XFILL_2__7298_ vdd gnd FILL
XFILL_0__10835_ vdd gnd FILL
XFILL_0__8121_ vdd gnd FILL
XFILL_2_BUFX2_insert380 vdd gnd FILL
XFILL_1__10036_ vdd gnd FILL
XFILL_1__14913_ vdd gnd FILL
XFILL_2__12375_ vdd gnd FILL
XFILL_0__13554_ vdd gnd FILL
X_7700_ _7700_/A _7700_/B _7700_/Y vdd gnd OR2X2
XFILL_0__8052_ vdd gnd FILL
X_8680_ _8680_/A _8680_/B _8680_/Y vdd gnd NAND2X1
XFILL_0__12505_ vdd gnd FILL
XFILL_1__14844_ vdd gnd FILL
X_7631_ _7631_/A _7631_/B _7631_/C _7631_/Y vdd gnd NAND3X1
XFILL_0__12436_ vdd gnd FILL
XFILL_1__14775_ vdd gnd FILL
XFILL_1__11987_ vdd gnd FILL
X_7562_ _7562_/A _7562_/B _7562_/C _7562_/Y vdd gnd OAI21X1
XFILL_2__10208_ vdd gnd FILL
XFILL_1__10938_ vdd gnd FILL
XFILL_1__13726_ vdd gnd FILL
X_9301_ _9301_/A _9301_/B _9301_/Y vdd gnd NAND2X1
XFILL_0__12367_ vdd gnd FILL
XFILL_0__8954_ vdd gnd FILL
X_7493_ _7493_/A _7493_/B _7493_/Y vdd gnd NAND2X1
XFILL_2__10139_ vdd gnd FILL
XFILL_0__14106_ vdd gnd FILL
XFILL_0__11318_ vdd gnd FILL
XFILL_1__13657_ vdd gnd FILL
XFILL_1__10869_ vdd gnd FILL
X_9232_ _9232_/A _9232_/B _9232_/C _9232_/Y vdd gnd OAI21X1
XFILL_0__7905_ vdd gnd FILL
XFILL_0__12298_ vdd gnd FILL
XFILL_0__14037_ vdd gnd FILL
XFILL_0__11249_ vdd gnd FILL
XFILL_1__13588_ vdd gnd FILL
X_9163_ _9163_/A _9163_/B _9163_/Y vdd gnd NOR2X1
XFILL_0__7836_ vdd gnd FILL
X_8114_ _8114_/A _8114_/B _8114_/S _8114_/Y vdd gnd MUX2X1
X_9094_ _9094_/A _9094_/B _9094_/C _9094_/Y vdd gnd NAND3X1
XFILL_0__7767_ vdd gnd FILL
XFILL_0__9506_ vdd gnd FILL
X_8045_ _8045_/A _8045_/B _8045_/C _8045_/D _8045_/Y vdd gnd AOI22X1
XFILL_0__7698_ vdd gnd FILL
XFILL_0__9437_ vdd gnd FILL
XFILL_1__8230_ vdd gnd FILL
XFILL_0__9368_ vdd gnd FILL
XFILL_1__8161_ vdd gnd FILL
X_9996_ _9996_/A _9996_/B _9996_/Y vdd gnd NOR2X1
XFILL_1__7112_ vdd gnd FILL
XFILL_0__8319_ vdd gnd FILL
XFILL_1__8092_ vdd gnd FILL
X_8947_ _8947_/A _8947_/Y vdd gnd INVX1
XFILL_0__9299_ vdd gnd FILL
X_8878_ _8878_/D _8878_/CLK _8878_/Q vdd gnd DFFPOSX1
X_7829_ _7829_/A _7829_/B _7829_/Y vdd gnd NAND2X1
XFILL_1__8994_ vdd gnd FILL
X_11430_ _11430_/A _11430_/B _11430_/C _11430_/Y vdd gnd AOI21X1
X_11361_ _11361_/A _11361_/B _11361_/Y vdd gnd OR2X2
XFILL_1__7876_ vdd gnd FILL
X_13100_ _13100_/A _13100_/B _13100_/Y vdd gnd NAND2X1
X_10312_ _10312_/A _10312_/B _10312_/Y vdd gnd NOR2X1
XFILL_1__9615_ vdd gnd FILL
X_14080_ _14080_/A _14080_/B _14080_/C _14080_/Y vdd gnd NAND3X1
X_11292_ _11292_/A _11292_/B _11292_/C _11292_/Y vdd gnd OAI21X1
XFILL257550x169350 vdd gnd FILL
X_10243_ _10243_/A _10243_/B _10243_/C _10243_/Y vdd gnd OAI21X1
X_13031_ _13031_/A _13031_/B _13031_/Y vdd gnd NAND2X1
XFILL_1__9546_ vdd gnd FILL
X_10174_ _10174_/A _10174_/B _10174_/Y vdd gnd NAND2X1
XFILL_1__9477_ vdd gnd FILL
XFILL_1__8428_ vdd gnd FILL
X_13933_ _13933_/A _13933_/B _13933_/Y vdd gnd OR2X2
XFILL_1__8359_ vdd gnd FILL
X_13864_ _13864_/A _13864_/B _13864_/Y vdd gnd NOR2X1
XFILL_0__10620_ vdd gnd FILL
XFILL_1_BUFX2_insert310 vdd gnd FILL
X_12815_ _12815_/A _12815_/B _12815_/C _12815_/D _12815_/Y vdd gnd AOI22X1
XFILL_1_BUFX2_insert321 vdd gnd FILL
XFILL_2__12160_ vdd gnd FILL
XFILL_1_BUFX2_insert332 vdd gnd FILL
X_13795_ _13795_/A _13795_/B _13795_/C _13795_/Y vdd gnd OAI21X1
XFILL_1__11910_ vdd gnd FILL
XFILL_1_BUFX2_insert343 vdd gnd FILL
XFILL_0__10551_ vdd gnd FILL
XFILL_1__12890_ vdd gnd FILL
XFILL_1_BUFX2_insert354 vdd gnd FILL
XFILL_1_BUFX2_insert365 vdd gnd FILL
X_12746_ _12746_/A _12746_/B _12746_/S _12746_/Y vdd gnd MUX2X1
XFILL_1_BUFX2_insert376 vdd gnd FILL
XFILL_1__11841_ vdd gnd FILL
XFILL_2__12091_ vdd gnd FILL
XFILL_0__13270_ vdd gnd FILL
XFILL_0__10482_ vdd gnd FILL
X_12677_ _12677_/A _12677_/B _12677_/S _12677_/Y vdd gnd MUX2X1
XFILL_0__12221_ vdd gnd FILL
XFILL_1__14560_ vdd gnd FILL
XFILL_1__11772_ vdd gnd FILL
X_14416_ _14416_/A _14416_/B _14416_/Y vdd gnd NAND2X1
X_11628_ _11628_/D _11628_/CLK _11628_/Q vdd gnd DFFPOSX1
XFILL_2__9724_ vdd gnd FILL
XFILL_1__13511_ vdd gnd FILL
XFILL_1__14491_ vdd gnd FILL
XFILL_0__12152_ vdd gnd FILL
X_14347_ _14347_/A _14347_/B _14347_/Y vdd gnd NAND2X1
XFILL_2__14801_ vdd gnd FILL
X_11559_ _11559_/A _11559_/B _11559_/C _11559_/Y vdd gnd OAI21X1
XFILL_2__9655_ vdd gnd FILL
XFILL_0__11103_ vdd gnd FILL
XFILL_1__10654_ vdd gnd FILL
XFILL_0__12083_ vdd gnd FILL
XFILL_2__12993_ vdd gnd FILL
XFILL_0__8670_ vdd gnd FILL
X_14278_ _14278_/A _14278_/B _14278_/Y vdd gnd NAND2X1
XFILL_2__14732_ vdd gnd FILL
XFILL_0__11034_ vdd gnd FILL
XFILL_2__9586_ vdd gnd FILL
XFILL_1__13373_ vdd gnd FILL
XFILL_1__10585_ vdd gnd FILL
XFILL_0__7621_ vdd gnd FILL
X_13229_ _13229_/A _13229_/B _13229_/Y vdd gnd NOR2X1
XFILL_1__12324_ vdd gnd FILL
XFILL_0__7552_ vdd gnd FILL
XFILL_1__12255_ vdd gnd FILL
XFILL_0__12985_ vdd gnd FILL
XFILL_1__11206_ vdd gnd FILL
XFILL_0__7483_ vdd gnd FILL
XFILL_0__14724_ vdd gnd FILL
XFILL_0__11936_ vdd gnd FILL
XFILL_1__12186_ vdd gnd FILL
XFILL_0__9222_ vdd gnd FILL
X_9850_ _9850_/A _9850_/B _9850_/Y vdd gnd NOR2X1
XFILL_1__11137_ vdd gnd FILL
XFILL_0__14655_ vdd gnd FILL
XFILL_0__11867_ vdd gnd FILL
XFILL_0__9153_ vdd gnd FILL
X_8801_ _8801_/A _8801_/B _8801_/C _8801_/Y vdd gnd OAI21X1
X_9781_ _9781_/D _9781_/CLK _9781_/Q vdd gnd DFFPOSX1
XFILL_2__12427_ vdd gnd FILL
XFILL_1__11068_ vdd gnd FILL
XFILL_0__10818_ vdd gnd FILL
XFILL_0__13606_ vdd gnd FILL
XFILL_0__14586_ vdd gnd FILL
XFILL_0__8104_ vdd gnd FILL
XFILL_0__11798_ vdd gnd FILL
XFILL_0__9084_ vdd gnd FILL
X_8732_ _8732_/A _8732_/B _8732_/Y vdd gnd NAND2X1
XFILL257550x234150 vdd gnd FILL
XFILL_1__10019_ vdd gnd FILL
XFILL_2__12358_ vdd gnd FILL
XFILL_0__13537_ vdd gnd FILL
XFILL_0__8035_ vdd gnd FILL
X_8663_ _8663_/A _8663_/B _8663_/C _8663_/Y vdd gnd OAI21X1
XFILL_1__14827_ vdd gnd FILL
XFILL_2__12289_ vdd gnd FILL
X_7614_ _7614_/A _7614_/B _7614_/C _7614_/Y vdd gnd OAI21X1
X_8594_ _8594_/A _8594_/B _8594_/Y vdd gnd NAND2X1
XFILL_2__14028_ vdd gnd FILL
XFILL_0__12419_ vdd gnd FILL
XFILL_1__14758_ vdd gnd FILL
XFILL_0__13399_ vdd gnd FILL
X_7545_ _7545_/A _7545_/B _7545_/C _7545_/Y vdd gnd NAND3X1
XFILL_0__9986_ vdd gnd FILL
XFILL_1__13709_ vdd gnd FILL
XFILL_1__14689_ vdd gnd FILL
XFILL_0__8937_ vdd gnd FILL
XFILL_1__7730_ vdd gnd FILL
X_7476_ _7476_/A _7476_/B _7476_/C _7476_/Y vdd gnd OAI21X1
X_9215_ _9215_/A _9215_/Y vdd gnd INVX1
XFILL_1__7661_ vdd gnd FILL
XFILL_1__9400_ vdd gnd FILL
X_9146_ _9146_/A _9146_/B _9146_/C _9146_/Y vdd gnd OAI21X1
XFILL_0__7819_ vdd gnd FILL
XFILL_1__7592_ vdd gnd FILL
XFILL_0__8799_ vdd gnd FILL
XFILL_1__9331_ vdd gnd FILL
X_9077_ _9077_/A _9077_/B _9077_/C _9077_/Y vdd gnd OAI21X1
X_8028_ _8028_/A _8028_/B _8028_/Y vdd gnd NAND2X1
XFILL_1__9262_ vdd gnd FILL
XFILL_1__8213_ vdd gnd FILL
XFILL_1__9193_ vdd gnd FILL
X_10930_ _10930_/A _10930_/Y vdd gnd INVX1
XFILL_1__8144_ vdd gnd FILL
X_9979_ _9979_/A _9979_/B _9979_/Y vdd gnd NAND2X1
X_10861_ _10861_/A _10861_/B _10861_/C _10861_/Y vdd gnd AOI21X1
XFILL_1__8075_ vdd gnd FILL
XFILL257550x144150 vdd gnd FILL
X_12600_ _12600_/D _12600_/CLK _12600_/Q vdd gnd DFFPOSX1
X_13580_ _13580_/A _13580_/B _13580_/C _13580_/Y vdd gnd NAND3X1
X_10792_ _10792_/A _10792_/Y vdd gnd INVX1
XFILL_0_BUFX2_insert306 vdd gnd FILL
X_12531_ _12531_/A _12531_/B _12531_/C _12531_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert317 vdd gnd FILL
XFILL_0_BUFX2_insert328 vdd gnd FILL
XFILL_0_BUFX2_insert339 vdd gnd FILL
X_12462_ _12462_/A _12462_/B _12462_/C _12462_/Y vdd gnd OAI21X1
XFILL_1__8977_ vdd gnd FILL
XFILL_2__7770_ vdd gnd FILL
X_14201_ _14201_/D _14201_/CLK _14201_/Q vdd gnd DFFPOSX1
X_11413_ _11413_/A _11413_/B _11413_/Y vdd gnd NOR2X1
X_12393_ _12393_/A _12393_/B _12393_/Y vdd gnd NAND2X1
X_14132_ _14132_/A _14132_/B _14132_/C _14132_/Y vdd gnd OAI21X1
X_11344_ _11344_/A _11344_/B _11344_/Y vdd gnd NAND2X1
XFILL_1__7859_ vdd gnd FILL
X_14063_ _14063_/A _14063_/B _14063_/Y vdd gnd NAND2X1
X_11275_ _11275_/A _11275_/Y vdd gnd INVX1
XFILL_1__10370_ vdd gnd FILL
X_13014_ _13014_/A _13014_/B _13014_/C _13014_/Y vdd gnd AOI21X1
X_10226_ _10226_/A _10226_/B _10226_/C _10226_/Y vdd gnd OAI21X1
XFILL_1__9529_ vdd gnd FILL
XFILL_2__8322_ vdd gnd FILL
X_10157_ _10157_/A _10157_/B _10157_/C _10157_/Y vdd gnd NAND3X1
XFILL_2__10611_ vdd gnd FILL
XFILL_1__12040_ vdd gnd FILL
XFILL_2__8253_ vdd gnd FILL
XFILL_0__12770_ vdd gnd FILL
X_10088_ _10088_/A _10088_/B _10088_/C _10088_/Y vdd gnd OAI21X1
XFILL_2__10542_ vdd gnd FILL
XFILL_2__8184_ vdd gnd FILL
XFILL_0__11721_ vdd gnd FILL
X_13916_ _13916_/A _13916_/B _13916_/C _13916_/Y vdd gnd AOI21X1
X_14896_ _14896_/D _14896_/CLK _14896_/Q vdd gnd DFFPOSX1
XFILL_2__10473_ vdd gnd FILL
XFILL_0__14440_ vdd gnd FILL
XFILL_1__13991_ vdd gnd FILL
X_13847_ _13847_/A _13847_/B _13847_/Y vdd gnd NAND2X1
XFILL_0__10603_ vdd gnd FILL
XFILL_1__12942_ vdd gnd FILL
XFILL_0__14371_ vdd gnd FILL
XFILL_1_BUFX2_insert140 vdd gnd FILL
XFILL_0__11583_ vdd gnd FILL
XFILL_1_BUFX2_insert151 vdd gnd FILL
X_13778_ _13778_/A _13778_/B _13778_/C _13778_/Y vdd gnd OAI21X1
XFILL_1_BUFX2_insert162 vdd gnd FILL
XFILL_2__12143_ vdd gnd FILL
XFILL_0__13322_ vdd gnd FILL
XFILL_0__10534_ vdd gnd FILL
XFILL_1_BUFX2_insert173 vdd gnd FILL
XFILL_1_BUFX2_insert184 vdd gnd FILL
XFILL_1__12873_ vdd gnd FILL
X_12729_ _12729_/A _12729_/B _12729_/S _12729_/Y vdd gnd MUX2X1
XFILL_1_BUFX2_insert195 vdd gnd FILL
XFILL_1__14612_ vdd gnd FILL
XFILL_2__12074_ vdd gnd FILL
XFILL_1__11824_ vdd gnd FILL
XFILL_0__13253_ vdd gnd FILL
XFILL_0__10465_ vdd gnd FILL
XFILL_0__12204_ vdd gnd FILL
XFILL_0__13184_ vdd gnd FILL
XFILL_1__11755_ vdd gnd FILL
XFILL_0__10396_ vdd gnd FILL
X_7330_ _7330_/A _7330_/Y vdd gnd INVX1
XFILL_0__12135_ vdd gnd FILL
XFILL_2__7899_ vdd gnd FILL
XFILL_1__14474_ vdd gnd FILL
XFILL_0__8722_ vdd gnd FILL
X_7261_ _7261_/A _7261_/B _7261_/C _7261_/Y vdd gnd OAI21X1
XFILL_1__10637_ vdd gnd FILL
XFILL_1__13425_ vdd gnd FILL
X_9000_ _9000_/A _9000_/B _9000_/Y vdd gnd NAND2X1
XFILL_0__12066_ vdd gnd FILL
XFILL_0__8653_ vdd gnd FILL
X_7192_ _7192_/A _7192_/B _7192_/S _7192_/Y vdd gnd MUX2X1
XFILL_2__14715_ vdd gnd FILL
XFILL_2__11927_ vdd gnd FILL
XFILL_0__11017_ vdd gnd FILL
XFILL_1__10568_ vdd gnd FILL
XFILL_1__13356_ vdd gnd FILL
XFILL_0__7604_ vdd gnd FILL
XFILL_0__8584_ vdd gnd FILL
XFILL_2__14646_ vdd gnd FILL
XFILL_1__12307_ vdd gnd FILL
XFILL_1__13287_ vdd gnd FILL
XFILL_1__10499_ vdd gnd FILL
XFILL_0__7535_ vdd gnd FILL
XFILL_1__12238_ vdd gnd FILL
XFILL_2__14577_ vdd gnd FILL
XFILL_0__12968_ vdd gnd FILL
X_9902_ _9902_/A _9902_/Y vdd gnd INVX1
XFILL_0__7466_ vdd gnd FILL
XFILL_0__14707_ vdd gnd FILL
XFILL_1__12169_ vdd gnd FILL
XFILL_0__9205_ vdd gnd FILL
XFILL_0__11919_ vdd gnd FILL
XFILL_0__12899_ vdd gnd FILL
X_9833_ _9833_/D _9833_/CLK _9833_/Q vdd gnd DFFPOSX1
XFILL_0__7397_ vdd gnd FILL
XFILL_0__14638_ vdd gnd FILL
XFILL_0__9136_ vdd gnd FILL
X_9764_ _9764_/D _9764_/CLK _9764_/Q vdd gnd DFFPOSX1
XFILL_0__14569_ vdd gnd FILL
XFILL_0__9067_ vdd gnd FILL
X_8715_ _8715_/A _8715_/B _8715_/Y vdd gnd OR2X2
X_9695_ _9695_/A _9695_/B _9695_/Y vdd gnd NAND2X1
XFILL_0__8018_ vdd gnd FILL
XFILL_1__9880_ vdd gnd FILL
X_8646_ _8646_/A _8646_/B _8646_/Y vdd gnd NAND2X1
XFILL_1__8831_ vdd gnd FILL
X_8577_ _8577_/A _8577_/B _8577_/C _8577_/Y vdd gnd OAI21X1
X_7528_ _7528_/A _7528_/B _7528_/C _7528_/D _7528_/Y vdd gnd AOI22X1
XFILL_0__9969_ vdd gnd FILL
XFILL_1__8762_ vdd gnd FILL
XFILL_1__7713_ vdd gnd FILL
X_7459_ _7459_/A _7459_/B _7459_/Y vdd gnd NAND2X1
XFILL_1__8693_ vdd gnd FILL
XFILL_1__7644_ vdd gnd FILL
X_11060_ _11060_/A _11060_/B _11060_/C _11060_/Y vdd gnd OAI21X1
X_9129_ _9129_/A _9129_/B _9129_/C _9129_/Y vdd gnd NAND3X1
XFILL_1__7575_ vdd gnd FILL
X_10011_ _10011_/A _10011_/B _10011_/C _10011_/Y vdd gnd OAI21X1
XFILL_1__9314_ vdd gnd FILL
XFILL_1__9245_ vdd gnd FILL
X_14750_ _14750_/A _14750_/B _14750_/C _14750_/Y vdd gnd OAI21X1
X_11962_ _11962_/A _11962_/B _11962_/Y vdd gnd NAND2X1
XFILL_1__9176_ vdd gnd FILL
X_13701_ _13701_/A _13701_/B _13701_/C _13701_/Y vdd gnd NAND3X1
X_10913_ _10913_/A _10913_/Y vdd gnd INVX1
X_14681_ _14681_/A _14681_/B _14681_/Y vdd gnd AND2X2
XFILL_1__8127_ vdd gnd FILL
X_11893_ _11893_/A _11893_/B _11893_/Y vdd gnd AND2X2
X_13632_ _13632_/A _13632_/B _13632_/C _13632_/Y vdd gnd OAI21X1
X_10844_ _10844_/A _10844_/B _10844_/S _10844_/Y vdd gnd MUX2X1
XFILL_2__8940_ vdd gnd FILL
XFILL_1__8058_ vdd gnd FILL
X_13563_ _13563_/A _13563_/B _13563_/Y vdd gnd NOR2X1
X_10775_ _10775_/A _10775_/B _10775_/C _10775_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert114 vdd gnd FILL
XFILL_0_BUFX2_insert125 vdd gnd FILL
XFILL_0_BUFX2_insert136 vdd gnd FILL
X_12514_ _12514_/A _12514_/Y vdd gnd INVX1
XFILL_0_BUFX2_insert147 vdd gnd FILL
XFILL_2__7822_ vdd gnd FILL
XFILL_0_BUFX2_insert158 vdd gnd FILL
X_13494_ _13494_/D _13494_/CLK _13494_/Q vdd gnd DFFPOSX1
XFILL_0__10250_ vdd gnd FILL
XFILL_0_BUFX2_insert169 vdd gnd FILL
X_12445_ _12445_/A _12445_/B _12445_/Y vdd gnd NAND2X1
XFILL_2__7753_ vdd gnd FILL
XFILL_1__11540_ vdd gnd FILL
XFILL_0__10181_ vdd gnd FILL
X_12376_ _12376_/A _12376_/B _12376_/Y vdd gnd NAND2X1
XFILL_2__7684_ vdd gnd FILL
XFILL_1__11471_ vdd gnd FILL
X_14115_ _14115_/A _14115_/B _14115_/C _14115_/Y vdd gnd OAI21X1
X_11327_ _11327_/A _11327_/B _11327_/C _11327_/Y vdd gnd NAND3X1
XFILL_1__13210_ vdd gnd FILL
XFILL_1__10422_ vdd gnd FILL
XFILL_0__13940_ vdd gnd FILL
X_14046_ _14046_/A _14046_/B _14046_/Y vdd gnd NAND2X1
X_11258_ _11258_/A _11258_/B _11258_/C _11258_/Y vdd gnd OAI21X1
XFILL_1__13141_ vdd gnd FILL
XFILL_2__11712_ vdd gnd FILL
XFILL_1__10353_ vdd gnd FILL
X_10209_ _10209_/A _10209_/B _10209_/C _10209_/Y vdd gnd OAI21X1
XFILL_0__13871_ vdd gnd FILL
XFILL_2__8305_ vdd gnd FILL
X_11189_ _11189_/A _11189_/B _11189_/Y vdd gnd NAND2X1
XFILL_1__13072_ vdd gnd FILL
XFILL_1__10284_ vdd gnd FILL
XFILL_0__12822_ vdd gnd FILL
XFILL_0__7320_ vdd gnd FILL
XFILL_1__12023_ vdd gnd FILL
XFILL_2__8236_ vdd gnd FILL
XFILL_0__12753_ vdd gnd FILL
XFILL_0__7251_ vdd gnd FILL
XFILL_2__13313_ vdd gnd FILL
XFILL_2__10525_ vdd gnd FILL
XFILL_0__11704_ vdd gnd FILL
XFILL_2__8167_ vdd gnd FILL
XFILL_0__12684_ vdd gnd FILL
XFILL_0__7182_ vdd gnd FILL
X_14879_ _14879_/D _14879_/CLK _14879_/Q vdd gnd DFFPOSX1
XFILL_2__10456_ vdd gnd FILL
XFILL_2__8098_ vdd gnd FILL
XFILL_0__14423_ vdd gnd FILL
XFILL_1__13974_ vdd gnd FILL
XFILL_2__10387_ vdd gnd FILL
XFILL_0__14354_ vdd gnd FILL
XFILL_1__12925_ vdd gnd FILL
XFILL_0__11566_ vdd gnd FILL
X_8500_ _8500_/A _8500_/B _8500_/C _8500_/Y vdd gnd OAI21X1
X_9480_ _9480_/A _9480_/B _9480_/Y vdd gnd NAND2X1
XFILL_0__13305_ vdd gnd FILL
XFILL_0__10517_ vdd gnd FILL
XFILL_0__14285_ vdd gnd FILL
XFILL_1__12856_ vdd gnd FILL
XFILL_0__11497_ vdd gnd FILL
X_8431_ _8431_/A _8431_/B _8431_/C _8431_/Y vdd gnd OAI21X1
XFILL_1__11807_ vdd gnd FILL
XFILL_0__13236_ vdd gnd FILL
XFILL_0__10448_ vdd gnd FILL
XFILL_1__12787_ vdd gnd FILL
X_8362_ _8362_/A _8362_/B _8362_/Y vdd gnd NAND2X1
XFILL_2__11008_ vdd gnd FILL
XFILL_0__13167_ vdd gnd FILL
XFILL_1__11738_ vdd gnd FILL
XFILL_0__10379_ vdd gnd FILL
X_7313_ _7313_/A _7313_/B _7313_/Y vdd gnd NAND2X1
XFILL_0__9754_ vdd gnd FILL
X_8293_ _8293_/A _8293_/B _8293_/C _8293_/Y vdd gnd OAI21X1
XFILL_0__12118_ vdd gnd FILL
XFILL_1__14457_ vdd gnd FILL
XFILL_0__8705_ vdd gnd FILL
XFILL_0__13098_ vdd gnd FILL
X_7244_ _7244_/A _7244_/B _7244_/C _7244_/D _7244_/Y vdd gnd AOI22X1
XFILL_0__9685_ vdd gnd FILL
XFILL_1__13408_ vdd gnd FILL
XFILL_0__12049_ vdd gnd FILL
XFILL_1__14388_ vdd gnd FILL
XFILL_0__8636_ vdd gnd FILL
X_7175_ _7175_/A _7175_/Y vdd gnd INVX1
XFILL_1__13339_ vdd gnd FILL
XFILL_1__7360_ vdd gnd FILL
XFILL_0__8567_ vdd gnd FILL
XFILL_2__14629_ vdd gnd FILL
XFILL_0__7518_ vdd gnd FILL
XFILL_1__7291_ vdd gnd FILL
XFILL_0__8498_ vdd gnd FILL
XFILL_1__9030_ vdd gnd FILL
XFILL_0__7449_ vdd gnd FILL
X_9816_ _9816_/D _9816_/CLK _9816_/Q vdd gnd DFFPOSX1
XFILL_0__9119_ vdd gnd FILL
X_9747_ _9747_/A _9747_/B _9747_/C _9747_/Y vdd gnd OAI21X1
XFILL_1__9932_ vdd gnd FILL
XBUFX2_insert208 BUFX2_insert208/A BUFX2_insert208/Y vdd gnd BUFX2
XBUFX2_insert219 BUFX2_insert219/A BUFX2_insert219/Y vdd gnd BUFX2
X_9678_ _9678_/A _9678_/B _9678_/C _9678_/Y vdd gnd OAI21X1
X_10560_ _10560_/A _10560_/Y vdd gnd INVX1
XFILL_1__9863_ vdd gnd FILL
X_8629_ _8629_/A _8629_/B _8629_/Y vdd gnd NAND2X1
XFILL_1__8814_ vdd gnd FILL
X_10491_ _10491_/A _10491_/B _10491_/Y vdd gnd NAND2X1
X_12230_ _12230_/A _12230_/B _12230_/C _12230_/Y vdd gnd NAND3X1
XFILL_1__8745_ vdd gnd FILL
X_12161_ _12161_/A _12161_/B _12161_/C _12161_/Y vdd gnd OAI21X1
XFILL_1__8676_ vdd gnd FILL
X_11112_ _11112_/A _11112_/B _11112_/Y vdd gnd OR2X2
XFILL_1__7627_ vdd gnd FILL
X_12092_ _12092_/A _12092_/B _12092_/C _12092_/Y vdd gnd OAI21X1
X_11043_ _11043_/A _11043_/B _11043_/C _11043_/Y vdd gnd OAI21X1
XFILL_1__7558_ vdd gnd FILL
XFILL_1__7489_ vdd gnd FILL
X_14802_ _14802_/A _14802_/B _14802_/Y vdd gnd AND2X2
XFILL_1__9228_ vdd gnd FILL
X_12994_ _12994_/A _12994_/B _12994_/Y vdd gnd NAND2X1
X_14733_ _14733_/A _14733_/B _14733_/C _14733_/Y vdd gnd AOI21X1
X_11945_ _11945_/A _11945_/B _11945_/C _11945_/Y vdd gnd AOI21X1
XFILL_1__9159_ vdd gnd FILL
X_14664_ _14664_/A _14664_/B _14664_/Y vdd gnd NAND2X1
XFILL_2__10241_ vdd gnd FILL
X_11876_ _11876_/A _11876_/B _11876_/C _11876_/D _11876_/Y vdd gnd AOI22X1
XFILL_0__11420_ vdd gnd FILL
XFILL_1__10971_ vdd gnd FILL
X_13615_ _13615_/A _13615_/B _13615_/Y vdd gnd OR2X2
X_10827_ _10827_/A _10827_/Y vdd gnd INVX1
X_14595_ _14595_/A _14595_/B _14595_/Y vdd gnd NOR2X1
XFILL_2__10172_ vdd gnd FILL
XFILL_1__12710_ vdd gnd FILL
XFILL_0__11351_ vdd gnd FILL
XFILL_1__13690_ vdd gnd FILL
X_13546_ _13546_/A _13546_/Y vdd gnd INVX4
X_10758_ _10758_/D _10758_/CLK _10758_/Q vdd gnd DFFPOSX1
XFILL_0__10302_ vdd gnd FILL
XFILL_0__14070_ vdd gnd FILL
XFILL_1__12641_ vdd gnd FILL
XFILL_0__11282_ vdd gnd FILL
X_13477_ _13477_/D _13477_/CLK _13477_/Q vdd gnd DFFPOSX1
X_10689_ _10689_/D _10689_/CLK _10689_/Q vdd gnd DFFPOSX1
XFILL_0__13021_ vdd gnd FILL
XFILL_0__10233_ vdd gnd FILL
X_12428_ _12428_/A _12428_/B _12428_/Y vdd gnd NAND2X1
XFILL_1__14311_ vdd gnd FILL
XFILL_1__11523_ vdd gnd FILL
XFILL_0__10164_ vdd gnd FILL
X_12359_ _12359_/A _12359_/B _12359_/C _12359_/Y vdd gnd OAI21X1
XFILL_2__7667_ vdd gnd FILL
XFILL_1__14242_ vdd gnd FILL
XFILL_1__11454_ vdd gnd FILL
XFILL_0__10095_ vdd gnd FILL
XFILL_2_BUFX2_insert1 vdd gnd FILL
XFILL_0__9470_ vdd gnd FILL
XFILL_1__10405_ vdd gnd FILL
XFILL_0__13923_ vdd gnd FILL
XFILL_2__7598_ vdd gnd FILL
XFILL_1__11385_ vdd gnd FILL
XFILL_0__8421_ vdd gnd FILL
X_14029_ _14029_/A _14029_/B _14029_/Y vdd gnd NOR2X1
XFILL_1__13124_ vdd gnd FILL
XFILL_1__10336_ vdd gnd FILL
XFILL_0__13854_ vdd gnd FILL
XFILL_0__8352_ vdd gnd FILL
XFILL_1__13055_ vdd gnd FILL
X_8980_ _8980_/A _8980_/Y vdd gnd INVX8
XFILL_1__10267_ vdd gnd FILL
XFILL_0__12805_ vdd gnd FILL
XFILL_0__7303_ vdd gnd FILL
XFILL_0__10997_ vdd gnd FILL
XFILL_0__13785_ vdd gnd FILL
X_7931_ _7931_/D _7931_/CLK _7931_/Q vdd gnd DFFPOSX1
XFILL_0__8283_ vdd gnd FILL
XFILL_2__8219_ vdd gnd FILL
XFILL_1__12006_ vdd gnd FILL
XFILL_1__10198_ vdd gnd FILL
XFILL_0__12736_ vdd gnd FILL
XFILL_0__7234_ vdd gnd FILL
X_7862_ _7862_/A _7862_/B _7862_/Y vdd gnd NAND2X1
XFILL_2__10508_ vdd gnd FILL
XFILL_0__12667_ vdd gnd FILL
X_9601_ _9601_/A _9601_/B _9601_/Y vdd gnd NAND2X1
XFILL_0__7165_ vdd gnd FILL
XFILL_2__13227_ vdd gnd FILL
XFILL_2__10439_ vdd gnd FILL
X_7793_ _7793_/A _7793_/B _7793_/C _7793_/D _7793_/Y vdd gnd AOI22X1
XFILL_0__14406_ vdd gnd FILL
XFILL_1__13957_ vdd gnd FILL
X_9532_ _9532_/A _9532_/B _9532_/C _9532_/Y vdd gnd OAI21X1
XFILL_0__7096_ vdd gnd FILL
XFILL_2__13158_ vdd gnd FILL
XFILL_1__12908_ vdd gnd FILL
XFILL_0__14337_ vdd gnd FILL
XFILL_0__11549_ vdd gnd FILL
XFILL_1__13888_ vdd gnd FILL
X_9463_ _9463_/A _9463_/B _9463_/Y vdd gnd NOR2X1
XFILL_2__13089_ vdd gnd FILL
XFILL_1__12839_ vdd gnd FILL
XFILL_0__14268_ vdd gnd FILL
X_8414_ _8414_/A _8414_/B _8414_/Y vdd gnd NAND2X1
X_9394_ _9394_/A _9394_/B _9394_/Y vdd gnd NAND2X1
XFILL_0__13219_ vdd gnd FILL
X_8345_ _8345_/A _8345_/Y vdd gnd INVX1
XFILL_0__7998_ vdd gnd FILL
XFILL_0__9737_ vdd gnd FILL
XFILL_1__8530_ vdd gnd FILL
X_8276_ _8276_/A _8276_/B _8276_/C _8276_/Y vdd gnd OAI21X1
X_7227_ _7227_/A _7227_/B _7227_/C _7227_/Y vdd gnd AOI21X1
XFILL_0__9668_ vdd gnd FILL
XFILL_1__8461_ vdd gnd FILL
XFILL_1__7412_ vdd gnd FILL
XFILL_0__8619_ vdd gnd FILL
X_7158_ _7158_/A _7158_/B _7158_/Y vdd gnd NAND2X1
XFILL_0__9599_ vdd gnd FILL
XFILL_1__8392_ vdd gnd FILL
XFILL_1__7343_ vdd gnd FILL
X_7089_ _7089_/A _7089_/B _7089_/C _7089_/Y vdd gnd AOI21X1
XFILL_1__7274_ vdd gnd FILL
XFILL_1__9013_ vdd gnd FILL
X_11730_ _11730_/A _11730_/B _11730_/C _11730_/Y vdd gnd OAI21X1
X_11661_ _11661_/D _11661_/CLK _11661_/Q vdd gnd DFFPOSX1
X_13400_ _13400_/A _13400_/B _13400_/Y vdd gnd NAND2X1
X_10612_ _10612_/A _10612_/B _10612_/Y vdd gnd OR2X2
X_14380_ _14380_/A _14380_/B _14380_/C _14380_/Y vdd gnd AOI21X1
XFILL_1__9915_ vdd gnd FILL
X_11592_ _11592_/A _11592_/B _11592_/C _11592_/Y vdd gnd OAI21X1
X_13331_ _13331_/A _13331_/B _13331_/C _13331_/Y vdd gnd OAI21X1
X_10543_ _10543_/A _10543_/B _10543_/C _10543_/Y vdd gnd OAI21X1
XFILL_1__9846_ vdd gnd FILL
X_13262_ _13262_/A _13262_/B _13262_/C _13262_/Y vdd gnd OAI21X1
X_10474_ _10474_/A _10474_/B _10474_/C _10474_/Y vdd gnd OAI21X1
XFILL_2__8570_ vdd gnd FILL
X_12213_ _12213_/A _12213_/B _12213_/C _12213_/Y vdd gnd AOI21X1
X_13193_ _13193_/A _13193_/B _13193_/C _13193_/Y vdd gnd AOI21X1
XFILL_1__8728_ vdd gnd FILL
X_12144_ _12144_/A _12144_/B _12144_/Y vdd gnd NAND2X1
XFILL_1__8659_ vdd gnd FILL
X_12075_ _12075_/A _12075_/B _12075_/C _12075_/Y vdd gnd OAI21X1
XFILL_1__11170_ vdd gnd FILL
XFILL_0__10920_ vdd gnd FILL
X_11026_ _11026_/A _11026_/Y vdd gnd INVX1
XFILL_2__9122_ vdd gnd FILL
XFILL_1__10121_ vdd gnd FILL
XFILL_2__12460_ vdd gnd FILL
XFILL_0__10851_ vdd gnd FILL
XFILL_1__10052_ vdd gnd FILL
XFILL_2__12391_ vdd gnd FILL
XFILL_0__13570_ vdd gnd FILL
XFILL_0__10782_ vdd gnd FILL
X_12977_ _12977_/A _12977_/B _12977_/Y vdd gnd NOR2X1
XFILL_2__14130_ vdd gnd FILL
XFILL_0__12521_ vdd gnd FILL
XFILL_1__14860_ vdd gnd FILL
X_14716_ _14716_/A _14716_/B _14716_/Y vdd gnd AND2X2
X_11928_ _11928_/A _11928_/B _11928_/Y vdd gnd NAND2X1
XFILL_2__14061_ vdd gnd FILL
XFILL_1__13811_ vdd gnd FILL
XFILL_0__12452_ vdd gnd FILL
XFILL_1__14791_ vdd gnd FILL
X_14647_ _14647_/A _14647_/B _14647_/C _14647_/Y vdd gnd AOI21X1
X_11859_ _11859_/A _11859_/B _11859_/C _11859_/Y vdd gnd OAI21X1
XFILL_2__13012_ vdd gnd FILL
XFILL_0__11403_ vdd gnd FILL
XFILL_2__9955_ vdd gnd FILL
XFILL_1__13742_ vdd gnd FILL
XFILL_0__12383_ vdd gnd FILL
XFILL_1__10954_ vdd gnd FILL
XFILL_0__8970_ vdd gnd FILL
X_14578_ _14578_/A _14578_/B _14578_/C _14578_/Y vdd gnd OAI21X1
XFILL_0__11334_ vdd gnd FILL
XFILL_0__14122_ vdd gnd FILL
XFILL256950x64950 vdd gnd FILL
XFILL_1__13673_ vdd gnd FILL
X_13529_ _13529_/A _13529_/B _13529_/C _13529_/Y vdd gnd OAI21X1
XFILL_1__10885_ vdd gnd FILL
XFILL_2__8837_ vdd gnd FILL
XFILL_0__14053_ vdd gnd FILL
XFILL_1__12624_ vdd gnd FILL
XFILL_0__11265_ vdd gnd FILL
XFILL_0__7852_ vdd gnd FILL
XFILL_0__13004_ vdd gnd FILL
XFILL_0__10216_ vdd gnd FILL
X_8130_ _8130_/A _8130_/B _8130_/C _8130_/Y vdd gnd OAI21X1
XFILL_0__11196_ vdd gnd FILL
XFILL_0__7783_ vdd gnd FILL
XFILL_1__11506_ vdd gnd FILL
XFILL_0__10147_ vdd gnd FILL
XFILL_0__9522_ vdd gnd FILL
XFILL_1__12486_ vdd gnd FILL
X_8061_ _8061_/A _8061_/Y vdd gnd INVX1
XFILL_1__14225_ vdd gnd FILL
XFILL_1__11437_ vdd gnd FILL
XFILL_0__10078_ vdd gnd FILL
XFILL_0__9453_ vdd gnd FILL
XFILL_0__13906_ vdd gnd FILL
XFILL_1__14156_ vdd gnd FILL
XFILL_0__8404_ vdd gnd FILL
XFILL_1__11368_ vdd gnd FILL
XFILL_0__9384_ vdd gnd FILL
XFILL_1__13107_ vdd gnd FILL
XFILL_1__10319_ vdd gnd FILL
XFILL_1__11299_ vdd gnd FILL
XFILL_1__14087_ vdd gnd FILL
XFILL_0__13837_ vdd gnd FILL
XFILL_0__8335_ vdd gnd FILL
X_8963_ _8963_/A _8963_/B _8963_/C _8963_/Y vdd gnd OAI21X1
XFILL_1__13038_ vdd gnd FILL
XFILL_0__13768_ vdd gnd FILL
X_7914_ _7914_/A _7914_/B _7914_/Y vdd gnd NAND2X1
XFILL_0__8266_ vdd gnd FILL
XFILL_2__14328_ vdd gnd FILL
X_8894_ _8894_/D _8894_/CLK _8894_/Q vdd gnd DFFPOSX1
XFILL_0__12719_ vdd gnd FILL
XFILL_0__7217_ vdd gnd FILL
XFILL_0__13699_ vdd gnd FILL
X_7845_ _7845_/A _7845_/B _7845_/C _7845_/Y vdd gnd OAI21X1
XFILL_0__8197_ vdd gnd FILL
XFILL_2__14259_ vdd gnd FILL
XFILL_0_CLKBUF1_insert106 vdd gnd FILL
XFILL_0__7148_ vdd gnd FILL
X_7776_ _7776_/A _7776_/Y vdd gnd INVX1
X_9515_ _9515_/A _9515_/B _9515_/Y vdd gnd AND2X2
XFILL_0__7079_ vdd gnd FILL
XFILL_1__9700_ vdd gnd FILL
X_9446_ _9446_/A _9446_/B _9446_/C _9446_/Y vdd gnd OAI21X1
XFILL_1__7892_ vdd gnd FILL
XFILL_1__9631_ vdd gnd FILL
X_9377_ _9377_/A _9377_/B _9377_/C _9377_/Y vdd gnd AOI21X1
XFILL_1__9562_ vdd gnd FILL
X_8328_ _8328_/A _8328_/B _8328_/Y vdd gnd AND2X2
X_10190_ _10190_/A _10190_/B _10190_/Y vdd gnd NAND2X1
XFILL_1__8513_ vdd gnd FILL
XFILL_1__9493_ vdd gnd FILL
X_8259_ _8259_/A _8259_/Y vdd gnd INVX1
XFILL_1__8444_ vdd gnd FILL
XFILL_1__8375_ vdd gnd FILL
X_12900_ _12900_/A _12900_/B _12900_/C _12900_/Y vdd gnd NAND3X1
XFILL_1__7326_ vdd gnd FILL
X_13880_ _13880_/A _13880_/B _13880_/C _13880_/Y vdd gnd OAI21X1
X_12831_ _12831_/A _12831_/B _12831_/Y vdd gnd NAND2X1
XFILL_1__7257_ vdd gnd FILL
X_12762_ _12762_/A _12762_/Y vdd gnd INVX1
XFILL_1__7188_ vdd gnd FILL
X_14501_ _14501_/D _14501_/CLK _14501_/Q vdd gnd DFFPOSX1
X_11713_ _11713_/A _11713_/B _11713_/C _11713_/Y vdd gnd OAI21X1
X_12693_ _12693_/A _12693_/B _12693_/C _12693_/Y vdd gnd OAI21X1
X_14432_ _14432_/A _14432_/B _14432_/Y vdd gnd NAND2X1
X_11644_ _11644_/D _11644_/CLK _11644_/Q vdd gnd DFFPOSX1
X_14363_ _14363_/A _14363_/B _14363_/C _14363_/Y vdd gnd OAI21X1
X_11575_ _11575_/A _11575_/B _11575_/C _11575_/Y vdd gnd OAI21X1
XFILL_1__10670_ vdd gnd FILL
X_13314_ _13314_/A _13314_/B _13314_/C _13314_/D _13314_/Y vdd gnd AOI22X1
X_10526_ _10526_/A _10526_/B _10526_/Y vdd gnd OR2X2
X_14294_ _14294_/A _14294_/B _14294_/C _14294_/Y vdd gnd NAND3X1
XFILL_2__8622_ vdd gnd FILL
XFILL_0__11050_ vdd gnd FILL
XFILL_2__11960_ vdd gnd FILL
XFILL_2_CLKBUF1_insert48 vdd gnd FILL
X_13245_ _13245_/A _13245_/B _13245_/Y vdd gnd NAND2X1
X_10457_ _10457_/A _10457_/B _10457_/C _10457_/Y vdd gnd OAI21X1
XFILL_0__10001_ vdd gnd FILL
XFILL_2__8553_ vdd gnd FILL
XFILL_1__12340_ vdd gnd FILL
XFILL_2__11891_ vdd gnd FILL
X_13176_ _13176_/A _13176_/B _13176_/Y vdd gnd NAND2X1
XFILL_2__13630_ vdd gnd FILL
X_10388_ _10388_/A _10388_/Y vdd gnd INVX1
XFILL_2__8484_ vdd gnd FILL
XFILL_1__12271_ vdd gnd FILL
X_12127_ _12127_/A _12127_/B _12127_/C _12127_/Y vdd gnd OAI21X1
XFILL_1__14010_ vdd gnd FILL
XFILL_1__11222_ vdd gnd FILL
XFILL_0__14740_ vdd gnd FILL
XFILL_0__11952_ vdd gnd FILL
X_12058_ _12058_/A _12058_/B _12058_/Y vdd gnd NAND2X1
XFILL_0_CLKBUF1_insert30 vdd gnd FILL
XFILL_0_CLKBUF1_insert41 vdd gnd FILL
XFILL_1__11153_ vdd gnd FILL
XFILL_0_CLKBUF1_insert52 vdd gnd FILL
XFILL_0__10903_ vdd gnd FILL
X_11009_ _11009_/A _11009_/B _11009_/Y vdd gnd NAND2X1
XFILL_0__14671_ vdd gnd FILL
XFILL_0_BUFX2_insert19 vdd gnd FILL
XFILL_2__9105_ vdd gnd FILL
XFILL_0__11883_ vdd gnd FILL
XFILL_0_CLKBUF1_insert63 vdd gnd FILL
XFILL_1__10104_ vdd gnd FILL
XFILL_0_CLKBUF1_insert74 vdd gnd FILL
XFILL_0_CLKBUF1_insert85 vdd gnd FILL
XFILL_0__13622_ vdd gnd FILL
XFILL_1__11084_ vdd gnd FILL
XFILL_0_CLKBUF1_insert96 vdd gnd FILL
XFILL_0__8120_ vdd gnd FILL
XFILL_0__10834_ vdd gnd FILL
XFILL_2__9036_ vdd gnd FILL
XFILL_2_BUFX2_insert370 vdd gnd FILL
XFILL_1__10035_ vdd gnd FILL
XFILL_1__14912_ vdd gnd FILL
XFILL_0__13553_ vdd gnd FILL
XFILL_0__8051_ vdd gnd FILL
XFILL_2__14113_ vdd gnd FILL
XFILL_2__11325_ vdd gnd FILL
XFILL_1__14843_ vdd gnd FILL
XFILL_0__12504_ vdd gnd FILL
X_7630_ _7630_/A _7630_/B _7630_/C _7630_/Y vdd gnd AOI21X1
XFILL_2__14044_ vdd gnd FILL
XFILL_2__11256_ vdd gnd FILL
XFILL_1__14774_ vdd gnd FILL
XFILL_0__12435_ vdd gnd FILL
XFILL_1__11986_ vdd gnd FILL
X_7561_ _7561_/A _7561_/B _7561_/C _7561_/Y vdd gnd NAND3X1
XFILL_2__9938_ vdd gnd FILL
XFILL_1__13725_ vdd gnd FILL
XFILL_1__10937_ vdd gnd FILL
XFILL_0__12366_ vdd gnd FILL
X_9300_ _9300_/A _9300_/B _9300_/Y vdd gnd NAND2X1
XFILL_0__8953_ vdd gnd FILL
X_7492_ _7492_/A _7492_/B _7492_/Y vdd gnd NAND2X1
XFILL_0__11317_ vdd gnd FILL
XBUFX2_insert380 BUFX2_insert380/A BUFX2_insert380/Y vdd gnd BUFX2
XFILL_0__14105_ vdd gnd FILL
XFILL_1__13656_ vdd gnd FILL
XFILL_2__9869_ vdd gnd FILL
XFILL_0__7904_ vdd gnd FILL
XFILL_0__12297_ vdd gnd FILL
XFILL_1__10868_ vdd gnd FILL
X_9231_ _9231_/A _9231_/Y vdd gnd INVX1
XFILL_0__11248_ vdd gnd FILL
XFILL_0__14036_ vdd gnd FILL
XFILL_1__13587_ vdd gnd FILL
XFILL_0__7835_ vdd gnd FILL
XFILL_1__10799_ vdd gnd FILL
X_9162_ _9162_/A _9162_/B _9162_/C _9162_/Y vdd gnd AOI21X1
XFILL_0__11179_ vdd gnd FILL
X_8113_ _8113_/A _8113_/B _8113_/S _8113_/Y vdd gnd MUX2X1
XFILL_0__7766_ vdd gnd FILL
X_9093_ _9093_/A _9093_/B _9093_/C _9093_/Y vdd gnd OAI21X1
XFILL_0__9505_ vdd gnd FILL
XFILL_1__12469_ vdd gnd FILL
X_8044_ _8044_/A _8044_/B _8044_/C _8044_/Y vdd gnd OAI21X1
XFILL_0__7697_ vdd gnd FILL
XFILL_0__9436_ vdd gnd FILL
XFILL_1__14139_ vdd gnd FILL
XFILL_0__9367_ vdd gnd FILL
XFILL_1__8160_ vdd gnd FILL
X_9995_ _9995_/A _9995_/B _9995_/Y vdd gnd OR2X2
XFILL_1__7111_ vdd gnd FILL
XFILL_0__8318_ vdd gnd FILL
XFILL_0__9298_ vdd gnd FILL
X_8946_ _8946_/A _8946_/B _8946_/C _8946_/Y vdd gnd AOI21X1
XFILL_1__8091_ vdd gnd FILL
XFILL_0__8249_ vdd gnd FILL
X_8877_ _8877_/D _8877_/CLK _8877_/Q vdd gnd DFFPOSX1
X_7828_ _7828_/A _7828_/B _7828_/C _7828_/Y vdd gnd OAI21X1
XFILL_1__8993_ vdd gnd FILL
X_7759_ _7759_/A _7759_/B _7759_/Y vdd gnd NAND2X1
X_11360_ _11360_/A _11360_/B _11360_/Y vdd gnd NAND2X1
X_9429_ _9429_/A _9429_/B _9429_/Y vdd gnd NAND2X1
XFILL_1__7875_ vdd gnd FILL
X_10311_ _10311_/A _10311_/B _10311_/Y vdd gnd OR2X2
XFILL_1__9614_ vdd gnd FILL
X_11291_ _11291_/A _11291_/B _11291_/Y vdd gnd NOR2X1
X_13030_ _13030_/A _13030_/B _13030_/Y vdd gnd NAND2X1
X_10242_ _10242_/A _10242_/B _10242_/Y vdd gnd NAND2X1
XFILL_1__9545_ vdd gnd FILL
X_10173_ _10173_/A _10173_/B _10173_/C _10173_/Y vdd gnd OAI21X1
XFILL_1__9476_ vdd gnd FILL
XFILL_1__8427_ vdd gnd FILL
X_13932_ _13932_/A _13932_/B _13932_/C _13932_/Y vdd gnd OAI21X1
XFILL_1__8358_ vdd gnd FILL
X_13863_ _13863_/A _13863_/B _13863_/Y vdd gnd AND2X2
XFILL_1__7309_ vdd gnd FILL
XFILL_1__8289_ vdd gnd FILL
XFILL_1_BUFX2_insert300 vdd gnd FILL
X_12814_ _12814_/A _12814_/B _12814_/C _12814_/Y vdd gnd OAI21X1
XFILL_1_BUFX2_insert311 vdd gnd FILL
X_13794_ _13794_/A _13794_/Y vdd gnd INVX1
XFILL_1_BUFX2_insert322 vdd gnd FILL
XFILL_0__10550_ vdd gnd FILL
XFILL_1_BUFX2_insert333 vdd gnd FILL
XFILL_1_BUFX2_insert344 vdd gnd FILL
X_12745_ _12745_/A _12745_/B _12745_/C _12745_/Y vdd gnd AOI21X1
XFILL_1_BUFX2_insert355 vdd gnd FILL
XFILL_2__11110_ vdd gnd FILL
XFILL_1_BUFX2_insert366 vdd gnd FILL
XFILL_1__11840_ vdd gnd FILL
XFILL_1_BUFX2_insert377 vdd gnd FILL
XFILL_0__10481_ vdd gnd FILL
X_12676_ _12676_/A _12676_/B _12676_/C _12676_/Y vdd gnd OAI21X1
XFILL_2__11041_ vdd gnd FILL
XFILL_0__12220_ vdd gnd FILL
XFILL_1__11771_ vdd gnd FILL
X_14415_ _14415_/A _14415_/Y vdd gnd INVX1
X_11627_ _11627_/D _11627_/CLK _11627_/Q vdd gnd DFFPOSX1
XFILL_1__13510_ vdd gnd FILL
XFILL_0__12151_ vdd gnd FILL
XFILL_1__14490_ vdd gnd FILL
X_14346_ _14346_/A _14346_/B _14346_/C _14346_/Y vdd gnd NAND3X1
X_11558_ _11558_/A _11558_/B _11558_/Y vdd gnd NAND2X1
XFILL_0__11102_ vdd gnd FILL
XFILL_1__10653_ vdd gnd FILL
XFILL_0__12082_ vdd gnd FILL
X_10509_ _10509_/A _10509_/Y vdd gnd INVX1
X_14277_ _14277_/A _14277_/B _14277_/Y vdd gnd NOR2X1
XFILL_2__8605_ vdd gnd FILL
X_11489_ _11489_/A _11489_/B _11489_/C _11489_/D _11489_/Y vdd gnd AOI22X1
XFILL_0__11033_ vdd gnd FILL
XFILL_2__11943_ vdd gnd FILL
XFILL_1__13372_ vdd gnd FILL
XFILL_0__7620_ vdd gnd FILL
XFILL_1__10584_ vdd gnd FILL
X_13228_ _13228_/A _13228_/B _13228_/C _13228_/Y vdd gnd AOI21X1
XFILL_2__8536_ vdd gnd FILL
XFILL_2__14662_ vdd gnd FILL
XFILL_1__12323_ vdd gnd FILL
XFILL_2__11874_ vdd gnd FILL
X_13159_ _13159_/A _13159_/Y vdd gnd INVX1
XFILL_0__7551_ vdd gnd FILL
XFILL_2__13613_ vdd gnd FILL
XFILL_2__8467_ vdd gnd FILL
XFILL_2__14593_ vdd gnd FILL
XFILL_1__12254_ vdd gnd FILL
XFILL_0__12984_ vdd gnd FILL
XFILL_0__7482_ vdd gnd FILL
XFILL_2__13544_ vdd gnd FILL
XFILL_1__11205_ vdd gnd FILL
XFILL_0__14723_ vdd gnd FILL
XFILL_2__8398_ vdd gnd FILL
XFILL_0__9221_ vdd gnd FILL
XFILL_0__11935_ vdd gnd FILL
XFILL_1__12185_ vdd gnd FILL
XFILL_1__11136_ vdd gnd FILL
XFILL_0__14654_ vdd gnd FILL
XFILL_2__10687_ vdd gnd FILL
XFILL_0__9152_ vdd gnd FILL
XFILL256650x86550 vdd gnd FILL
XFILL_0__11866_ vdd gnd FILL
X_8800_ _8800_/A _8800_/B _8800_/Y vdd gnd NAND2X1
X_9780_ _9780_/D _9780_/CLK _9780_/Q vdd gnd DFFPOSX1
XFILL_1__11067_ vdd gnd FILL
XFILL_0__13605_ vdd gnd FILL
XFILL_0__8103_ vdd gnd FILL
XFILL_0__10817_ vdd gnd FILL
XFILL_0__14585_ vdd gnd FILL
XFILL_0__9083_ vdd gnd FILL
XFILL_2__9019_ vdd gnd FILL
X_8731_ _8731_/A _8731_/B _8731_/Y vdd gnd NAND2X1
XFILL_0__11797_ vdd gnd FILL
XFILL_1__10018_ vdd gnd FILL
XFILL_0__13536_ vdd gnd FILL
XFILL_0__8034_ vdd gnd FILL
X_8662_ _8662_/A _8662_/B _8662_/C _8662_/Y vdd gnd AOI21X1
XFILL_2__11308_ vdd gnd FILL
XFILL_1__14826_ vdd gnd FILL
XFILL_0__10679_ vdd gnd FILL
X_7613_ _7613_/A _7613_/B _7613_/Y vdd gnd NAND2X1
X_8593_ _8593_/A _8593_/B _8593_/C _8593_/Y vdd gnd OAI21X1
XFILL_2__11239_ vdd gnd FILL
XFILL_1__14757_ vdd gnd FILL
XFILL_0__12418_ vdd gnd FILL
XFILL_1__11969_ vdd gnd FILL
XFILL_0__13398_ vdd gnd FILL
X_7544_ _7544_/A _7544_/B _7544_/C _7544_/Y vdd gnd OAI21X1
XFILL_0__9985_ vdd gnd FILL
XFILL_1__13708_ vdd gnd FILL
XFILL_1__14688_ vdd gnd FILL
XFILL_0__12349_ vdd gnd FILL
XFILL_0__8936_ vdd gnd FILL
X_7475_ _7475_/A _7475_/B _7475_/S _7475_/Y vdd gnd MUX2X1
XFILL_1__13639_ vdd gnd FILL
X_9214_ _9214_/A _9214_/B _9214_/Y vdd gnd AND2X2
XFILL_1__7660_ vdd gnd FILL
XFILL_0__14019_ vdd gnd FILL
XFILL_0__7818_ vdd gnd FILL
X_9145_ _9145_/A _9145_/B _9145_/C _9145_/Y vdd gnd OAI21X1
XFILL_1__7591_ vdd gnd FILL
XFILL_0__8798_ vdd gnd FILL
XFILL_1__9330_ vdd gnd FILL
XFILL_0__7749_ vdd gnd FILL
X_9076_ _9076_/A _9076_/Y vdd gnd INVX2
XFILL_1__9261_ vdd gnd FILL
X_8027_ _8027_/A _8027_/B _8027_/C _8027_/D _8027_/Y vdd gnd AOI22X1
XFILL_0__9419_ vdd gnd FILL
XFILL_1__8212_ vdd gnd FILL
XFILL_1__9192_ vdd gnd FILL
XFILL_1__8143_ vdd gnd FILL
X_9978_ _9978_/A _9978_/B _9978_/C _9978_/Y vdd gnd OAI21X1
X_10860_ _10860_/A _10860_/B _10860_/Y vdd gnd NAND2X1
X_8929_ _8929_/A _8929_/B _8929_/Y vdd gnd AND2X2
XFILL_1__8074_ vdd gnd FILL
X_10791_ _10791_/A _10791_/B _10791_/Y vdd gnd NAND2X1
X_12530_ _12530_/A _12530_/B _12530_/C _12530_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert307 vdd gnd FILL
XFILL_0_BUFX2_insert318 vdd gnd FILL
XFILL_0_BUFX2_insert329 vdd gnd FILL
X_12461_ _12461_/A _12461_/B _12461_/C _12461_/Y vdd gnd OAI21X1
XFILL_1__8976_ vdd gnd FILL
X_14200_ _14200_/D _14200_/CLK _14200_/Q vdd gnd DFFPOSX1
X_11412_ _11412_/A _11412_/Y vdd gnd INVX1
X_12392_ _12392_/A _12392_/B _12392_/Y vdd gnd NAND2X1
X_14131_ _14131_/A _14131_/B _14131_/Y vdd gnd NAND2X1
X_11343_ _11343_/A _11343_/B _11343_/C _11343_/Y vdd gnd NAND3X1
XFILL_1__7858_ vdd gnd FILL
X_14062_ _14062_/A _14062_/B _14062_/Y vdd gnd NAND2X1
X_11274_ _11274_/A _11274_/B _11274_/C _11274_/Y vdd gnd NOR3X1
XFILL_1__7789_ vdd gnd FILL
X_13013_ _13013_/A _13013_/B _13013_/C _13013_/Y vdd gnd OAI21X1
X_10225_ _10225_/A _10225_/B _10225_/Y vdd gnd NAND2X1
XFILL_1__9528_ vdd gnd FILL
X_10156_ _10156_/A _10156_/B _10156_/C _10156_/Y vdd gnd OAI21X1
XFILL_1__9459_ vdd gnd FILL
XFILL_2__7203_ vdd gnd FILL
X_10087_ _10087_/A _10087_/B _10087_/Y vdd gnd NOR2X1
XFILL_0__11720_ vdd gnd FILL
X_13915_ _13915_/A _13915_/Y vdd gnd INVX1
XFILL_2__7134_ vdd gnd FILL
X_14895_ _14895_/D _14895_/CLK _14895_/Q vdd gnd DFFPOSX1
XFILL_2__13260_ vdd gnd FILL
XFILL_1__13990_ vdd gnd FILL
X_13846_ _13846_/A _13846_/B _13846_/C _13846_/Y vdd gnd OAI21X1
XFILL_2__13191_ vdd gnd FILL
XFILL_1__12941_ vdd gnd FILL
XFILL_0__10602_ vdd gnd FILL
XFILL256650x18150 vdd gnd FILL
XFILL_0__14370_ vdd gnd FILL
XFILL_0__11582_ vdd gnd FILL
XFILL_1_BUFX2_insert130 vdd gnd FILL
XFILL_1_BUFX2_insert141 vdd gnd FILL
X_13777_ _13777_/A _13777_/B _13777_/C _13777_/Y vdd gnd NAND3X1
X_10989_ _10989_/A _10989_/Y vdd gnd INVX1
XFILL_1_BUFX2_insert152 vdd gnd FILL
XFILL_0__10533_ vdd gnd FILL
XFILL_1_BUFX2_insert163 vdd gnd FILL
XFILL_0__13321_ vdd gnd FILL
XFILL_1_BUFX2_insert174 vdd gnd FILL
XFILL_1__12872_ vdd gnd FILL
X_12728_ _12728_/A _12728_/B _12728_/S _12728_/Y vdd gnd MUX2X1
XFILL_1_BUFX2_insert185 vdd gnd FILL
XFILL_1__14611_ vdd gnd FILL
XFILL_1_BUFX2_insert196 vdd gnd FILL
XFILL_1__11823_ vdd gnd FILL
XFILL_0__10464_ vdd gnd FILL
XFILL_0__13252_ vdd gnd FILL
X_12659_ _12659_/A _12659_/B _12659_/Y vdd gnd NAND2X1
XFILL_2__11024_ vdd gnd FILL
XFILL_0__12203_ vdd gnd FILL
XFILL_0__13183_ vdd gnd FILL
XFILL_1__11754_ vdd gnd FILL
XFILL_0__10395_ vdd gnd FILL
XFILL256050x216150 vdd gnd FILL
XFILL_0__12134_ vdd gnd FILL
XFILL_1__14473_ vdd gnd FILL
XFILL_0__8721_ vdd gnd FILL
X_14329_ _14329_/A _14329_/Y vdd gnd INVX1
X_7260_ _7260_/A _7260_/B _7260_/Y vdd gnd NAND2X1
XFILL_1__13424_ vdd gnd FILL
XFILL_1__10636_ vdd gnd FILL
XFILL_0__12065_ vdd gnd FILL
XFILL_0__8652_ vdd gnd FILL
X_7191_ _7191_/A _7191_/B _7191_/S _7191_/Y vdd gnd MUX2X1
XFILL_0__11016_ vdd gnd FILL
XFILL_1__13355_ vdd gnd FILL
XFILL_0__7603_ vdd gnd FILL
XFILL_1__10567_ vdd gnd FILL
XFILL_0__8583_ vdd gnd FILL
XFILL_1__12306_ vdd gnd FILL
XFILL_2__11857_ vdd gnd FILL
XFILL_1__13286_ vdd gnd FILL
XFILL_0__7534_ vdd gnd FILL
XFILL_1__10498_ vdd gnd FILL
XFILL_2__10808_ vdd gnd FILL
XFILL_1__12237_ vdd gnd FILL
XFILL_2__11788_ vdd gnd FILL
XFILL_0__12967_ vdd gnd FILL
X_9901_ _9901_/A _9901_/B _9901_/C _9901_/Y vdd gnd OAI21X1
XFILL_0__7465_ vdd gnd FILL
XFILL_2__13527_ vdd gnd FILL
XFILL_0__14706_ vdd gnd FILL
XFILL_0__9204_ vdd gnd FILL
XFILL_0__11918_ vdd gnd FILL
XFILL_1__12168_ vdd gnd FILL
XFILL_0__12898_ vdd gnd FILL
X_9832_ _9832_/D _9832_/CLK _9832_/Q vdd gnd DFFPOSX1
XFILL_0__7396_ vdd gnd FILL
XFILL_1__11119_ vdd gnd FILL
XFILL_0__14637_ vdd gnd FILL
XFILL_0__9135_ vdd gnd FILL
XFILL_0__11849_ vdd gnd FILL
XFILL_1__12099_ vdd gnd FILL
X_9763_ _9763_/A _9763_/B _9763_/C _9763_/Y vdd gnd OAI21X1
XFILL_2__13389_ vdd gnd FILL
XFILL_0__14568_ vdd gnd FILL
XFILL_0__9066_ vdd gnd FILL
X_8714_ _8714_/A _8714_/B _8714_/Y vdd gnd NAND2X1
X_9694_ _9694_/A _9694_/B _9694_/Y vdd gnd NAND2X1
XFILL_0__13519_ vdd gnd FILL
XFILL_0__8017_ vdd gnd FILL
XFILL_0__14499_ vdd gnd FILL
X_8645_ _8645_/A _8645_/B _8645_/Y vdd gnd NOR2X1
XFILL_1__14809_ vdd gnd FILL
XFILL_1__8830_ vdd gnd FILL
X_8576_ _8576_/A _8576_/B _8576_/C _8576_/Y vdd gnd OAI21X1
X_7527_ _7527_/A _7527_/B _7527_/Y vdd gnd NAND2X1
XFILL_1__8761_ vdd gnd FILL
XFILL_0__9968_ vdd gnd FILL
XFILL_1__7712_ vdd gnd FILL
X_7458_ _7458_/A _7458_/B _7458_/Y vdd gnd NOR2X1
XFILL_1__8692_ vdd gnd FILL
XFILL_0__9899_ vdd gnd FILL
XFILL_1__7643_ vdd gnd FILL
X_7389_ _7389_/A _7389_/B _7389_/Y vdd gnd AND2X2
X_9128_ _9128_/A _9128_/Y vdd gnd INVX1
XFILL_1__7574_ vdd gnd FILL
X_10010_ _10010_/A _10010_/B _10010_/Y vdd gnd NAND2X1
XFILL_1__9313_ vdd gnd FILL
X_9059_ _9059_/A _9059_/B _9059_/S _9059_/Y vdd gnd MUX2X1
XFILL_1__9244_ vdd gnd FILL
X_11961_ _11961_/A _11961_/B _11961_/C _11961_/Y vdd gnd NAND3X1
XFILL_1__9175_ vdd gnd FILL
X_10912_ _10912_/A _10912_/B _10912_/Y vdd gnd NAND2X1
X_13700_ _13700_/A _13700_/B _13700_/C _13700_/Y vdd gnd OAI21X1
X_14680_ _14680_/A _14680_/B _14680_/Y vdd gnd NAND2X1
XFILL_1__8126_ vdd gnd FILL
X_11892_ _11892_/A _11892_/B _11892_/Y vdd gnd NOR2X1
X_13631_ _13631_/A _13631_/Y vdd gnd INVX1
XFILL257550x46950 vdd gnd FILL
X_10843_ _10843_/A _10843_/B _10843_/S _10843_/Y vdd gnd MUX2X1
XFILL_1__8057_ vdd gnd FILL
X_13562_ _13562_/A _13562_/B _13562_/S _13562_/Y vdd gnd MUX2X1
X_10774_ _10774_/A _10774_/B _10774_/Y vdd gnd NOR2X1
XFILL_0_BUFX2_insert115 vdd gnd FILL
X_12513_ _12513_/A _12513_/B _12513_/C _12513_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert126 vdd gnd FILL
XFILL_0_BUFX2_insert137 vdd gnd FILL
X_13493_ _13493_/D _13493_/CLK _13493_/Q vdd gnd DFFPOSX1
XFILL_0_BUFX2_insert148 vdd gnd FILL
XFILL_0_BUFX2_insert159 vdd gnd FILL
X_12444_ _12444_/A _12444_/B _12444_/Y vdd gnd NAND2X1
XFILL_1__8959_ vdd gnd FILL
XFILL_0__10180_ vdd gnd FILL
X_12375_ _12375_/A _12375_/B _12375_/Y vdd gnd NAND2X1
XFILL_1__11470_ vdd gnd FILL
X_14114_ _14114_/A _14114_/B _14114_/Y vdd gnd NAND2X1
X_11326_ _11326_/A _11326_/B _11326_/C _11326_/Y vdd gnd AOI21X1
XFILL_1_CLKBUF1_insert384 vdd gnd FILL
XFILL_2__9422_ vdd gnd FILL
XFILL_1__10421_ vdd gnd FILL
XFILL_2__12760_ vdd gnd FILL
X_14045_ _14045_/A _14045_/B _14045_/C _14045_/Y vdd gnd NAND3X1
X_11257_ _11257_/A _11257_/B _11257_/C _11257_/Y vdd gnd NAND3X1
XFILL_2__9353_ vdd gnd FILL
XFILL_1__13140_ vdd gnd FILL
XFILL_2__12691_ vdd gnd FILL
XFILL_1__10352_ vdd gnd FILL
X_10208_ _10208_/A _10208_/B _10208_/Y vdd gnd NAND2X1
XFILL_0__13870_ vdd gnd FILL
XFILL_2__14430_ vdd gnd FILL
X_11188_ _11188_/A _11188_/B _11188_/Y vdd gnd NAND2X1
XFILL_2__9284_ vdd gnd FILL
XFILL_1__10283_ vdd gnd FILL
XFILL_0__12821_ vdd gnd FILL
XFILL_1__13071_ vdd gnd FILL
X_10139_ _10139_/A _10139_/Y vdd gnd INVX1
XFILL_2__14361_ vdd gnd FILL
XFILL_1__12022_ vdd gnd FILL
XFILL_2__11573_ vdd gnd FILL
XFILL_0__12752_ vdd gnd FILL
XFILL_0__7250_ vdd gnd FILL
XFILL_2__14292_ vdd gnd FILL
XFILL_0__11703_ vdd gnd FILL
XFILL_0__12683_ vdd gnd FILL
XFILL_2__7117_ vdd gnd FILL
XFILL_0__7181_ vdd gnd FILL
X_14878_ _14878_/D _14878_/CLK _14878_/Q vdd gnd DFFPOSX1
XFILL_2__13243_ vdd gnd FILL
XFILL_0__14422_ vdd gnd FILL
XFILL_1__13973_ vdd gnd FILL
X_13829_ _13829_/A _13829_/B _13829_/C _13829_/Y vdd gnd OAI21X1
XFILL_2__13174_ vdd gnd FILL
XFILL_1__12924_ vdd gnd FILL
XFILL_0__14353_ vdd gnd FILL
XFILL_0__11565_ vdd gnd FILL
XFILL_0__13304_ vdd gnd FILL
XFILL_0__10516_ vdd gnd FILL
XFILL_1__12855_ vdd gnd FILL
XFILL_0__14284_ vdd gnd FILL
X_8430_ _8430_/A _8430_/B _8430_/C _8430_/Y vdd gnd OAI21X1
XFILL_0__11496_ vdd gnd FILL
XFILL_1__11806_ vdd gnd FILL
XFILL_0__13235_ vdd gnd FILL
XFILL_0__10447_ vdd gnd FILL
XFILL_1__12786_ vdd gnd FILL
X_8361_ _8361_/A _8361_/B _8361_/C _8361_/Y vdd gnd OAI21X1
XFILL_1__11737_ vdd gnd FILL
XFILL_0__13166_ vdd gnd FILL
XFILL_0__10378_ vdd gnd FILL
X_7312_ _7312_/A _7312_/B _7312_/C _7312_/Y vdd gnd NAND3X1
XFILL_0__9753_ vdd gnd FILL
X_8292_ _8292_/A _8292_/B _8292_/C _8292_/Y vdd gnd AOI21X1
XFILL_1__14456_ vdd gnd FILL
XFILL_0__12117_ vdd gnd FILL
XFILL_0__8704_ vdd gnd FILL
XFILL_0__13097_ vdd gnd FILL
XFILL_0__9684_ vdd gnd FILL
X_7243_ _7243_/A _7243_/B _7243_/Y vdd gnd NOR2X1
XFILL_1__13407_ vdd gnd FILL
XFILL_1__10619_ vdd gnd FILL
XFILL_0__12048_ vdd gnd FILL
XFILL_1__14387_ vdd gnd FILL
XFILL_0__8635_ vdd gnd FILL
XFILL_1__11599_ vdd gnd FILL
X_7174_ _7174_/A _7174_/B _7174_/C _7174_/Y vdd gnd OAI21X1
XFILL_1__13338_ vdd gnd FILL
XFILL_0__8566_ vdd gnd FILL
XFILL_1__13269_ vdd gnd FILL
XFILL_0__7517_ vdd gnd FILL
XFILL_0__13999_ vdd gnd FILL
XFILL_1__7290_ vdd gnd FILL
XFILL_0__8497_ vdd gnd FILL
XFILL_0__7448_ vdd gnd FILL
X_9815_ _9815_/D _9815_/CLK _9815_/Q vdd gnd DFFPOSX1
XFILL_0__7379_ vdd gnd FILL
XFILL_0__9118_ vdd gnd FILL
X_9746_ _9746_/A _9746_/B _9746_/C _9746_/Y vdd gnd OAI21X1
XFILL_0__9049_ vdd gnd FILL
XBUFX2_insert209 BUFX2_insert209/A BUFX2_insert209/Y vdd gnd BUFX2
XFILL_1__9931_ vdd gnd FILL
X_9677_ _9677_/A _9677_/B _9677_/Y vdd gnd NAND2X1
X_8628_ _8628_/A _8628_/B _8628_/Y vdd gnd NOR2X1
XFILL_1__9862_ vdd gnd FILL
X_10490_ _10490_/A _10490_/B _10490_/Y vdd gnd NAND2X1
XFILL_1__8813_ vdd gnd FILL
X_8559_ _8559_/A _8559_/Y vdd gnd INVX1
XFILL_1__8744_ vdd gnd FILL
X_12160_ _12160_/A _12160_/B _12160_/Y vdd gnd NOR2X1
XFILL_1__8675_ vdd gnd FILL
X_11111_ _11111_/A _11111_/B _11111_/C _11111_/Y vdd gnd OAI21X1
XFILL257550x21750 vdd gnd FILL
X_12091_ _12091_/A _12091_/B _12091_/C _12091_/Y vdd gnd OAI21X1
XFILL_1__7626_ vdd gnd FILL
X_11042_ _11042_/A _11042_/B _11042_/C _11042_/Y vdd gnd OAI21X1
XFILL_1__7557_ vdd gnd FILL
XFILL_1__7488_ vdd gnd FILL
X_14801_ _14801_/A _14801_/B _14801_/Y vdd gnd NOR2X1
XFILL_1__9227_ vdd gnd FILL
X_12993_ _12993_/A _12993_/B _12993_/C _12993_/Y vdd gnd OAI21X1
X_14732_ _14732_/A _14732_/B _14732_/C _14732_/Y vdd gnd OAI21X1
XFILL_1__9158_ vdd gnd FILL
X_11944_ _11944_/A _11944_/B _11944_/C _11944_/Y vdd gnd NAND3X1
XFILL_1__8109_ vdd gnd FILL
X_14663_ _14663_/A _14663_/B _14663_/Y vdd gnd OR2X2
X_11875_ _11875_/A _11875_/B _11875_/C _11875_/Y vdd gnd OAI21X1
XFILL_1__9089_ vdd gnd FILL
XFILL_2__9971_ vdd gnd FILL
XFILL_1__10970_ vdd gnd FILL
X_13614_ _13614_/A _13614_/B _13614_/C _13614_/Y vdd gnd OAI21X1
X_10826_ _10826_/A _10826_/Y vdd gnd INVX1
X_14594_ _14594_/A _14594_/Y vdd gnd INVX2
XFILL_0__11350_ vdd gnd FILL
X_13545_ _13545_/A _13545_/Y vdd gnd INVX1
X_10757_ _10757_/D _10757_/CLK _10757_/Q vdd gnd DFFPOSX1
XFILL_0__10301_ vdd gnd FILL
XFILL_1__12640_ vdd gnd FILL
XFILL_0__11281_ vdd gnd FILL
X_13476_ _13476_/D _13476_/CLK _13476_/Q vdd gnd DFFPOSX1
X_10688_ _10688_/D _10688_/CLK _10688_/Q vdd gnd DFFPOSX1
XFILL_2__13930_ vdd gnd FILL
XFILL_0__10232_ vdd gnd FILL
XFILL_0__13020_ vdd gnd FILL
XFILL_2__8784_ vdd gnd FILL
X_12427_ _12427_/A _12427_/B _12427_/Y vdd gnd NAND2X1
XFILL_1__14310_ vdd gnd FILL
XFILL_1__11522_ vdd gnd FILL
XFILL_2__13861_ vdd gnd FILL
XFILL_0__10163_ vdd gnd FILL
X_12358_ _12358_/A _12358_/B _12358_/C _12358_/Y vdd gnd AOI21X1
XFILL_1__14241_ vdd gnd FILL
XFILL_2__12812_ vdd gnd FILL
XFILL_1__11453_ vdd gnd FILL
XFILL_2__13792_ vdd gnd FILL
XFILL_0__10094_ vdd gnd FILL
X_11309_ _11309_/A _11309_/B _11309_/Y vdd gnd NAND2X1
XFILL_2__9405_ vdd gnd FILL
X_12289_ _12289_/A _12289_/B _12289_/C _12289_/Y vdd gnd OAI21X1
XFILL_1__10404_ vdd gnd FILL
XFILL_2__12743_ vdd gnd FILL
XFILL_0__13922_ vdd gnd FILL
XFILL_0__8420_ vdd gnd FILL
XFILL_1__11384_ vdd gnd FILL
X_14028_ _14028_/A _14028_/B _14028_/C _14028_/Y vdd gnd OAI21X1
XFILL_1__13123_ vdd gnd FILL
XFILL_2__9336_ vdd gnd FILL
XFILL_1__10335_ vdd gnd FILL
XFILL_2__12674_ vdd gnd FILL
XFILL_0__13853_ vdd gnd FILL
XFILL_0__8351_ vdd gnd FILL
XFILL_2__14413_ vdd gnd FILL
XFILL_2__9267_ vdd gnd FILL
XFILL_0__12804_ vdd gnd FILL
XFILL_1__13054_ vdd gnd FILL
XFILL_0__7302_ vdd gnd FILL
XFILL_1__10266_ vdd gnd FILL
XFILL_0__13784_ vdd gnd FILL
XFILL_0__10996_ vdd gnd FILL
X_7930_ _7930_/D _7930_/CLK _7930_/Q vdd gnd DFFPOSX1
XFILL_0__8282_ vdd gnd FILL
XFILL_1__12005_ vdd gnd FILL
XFILL_2__14344_ vdd gnd FILL
XFILL_2__9198_ vdd gnd FILL
XFILL_2__11556_ vdd gnd FILL
XFILL_0__12735_ vdd gnd FILL
XFILL_1__10197_ vdd gnd FILL
XFILL_0__7233_ vdd gnd FILL
X_7861_ _7861_/A _7861_/B _7861_/C _7861_/Y vdd gnd OAI21X1
XFILL_2__14275_ vdd gnd FILL
XFILL_2__11487_ vdd gnd FILL
X_9600_ _9600_/A _9600_/B _9600_/Y vdd gnd OR2X2
XFILL_0__12666_ vdd gnd FILL
XFILL_0__7164_ vdd gnd FILL
X_7792_ _7792_/A _7792_/B _7792_/C _7792_/Y vdd gnd AOI21X1
XFILL_0__14405_ vdd gnd FILL
XFILL_1__13956_ vdd gnd FILL
X_9531_ _9531_/A _9531_/B _9531_/C _9531_/Y vdd gnd OAI21X1
XFILL_0__7095_ vdd gnd FILL
XFILL_1__12907_ vdd gnd FILL
XFILL_0__14336_ vdd gnd FILL
XFILL_1__13887_ vdd gnd FILL
XFILL_0__11548_ vdd gnd FILL
X_9462_ _9462_/A _9462_/B _9462_/C _9462_/Y vdd gnd OAI21X1
XFILL_2__12108_ vdd gnd FILL
XFILL_1__12838_ vdd gnd FILL
XFILL_0__14267_ vdd gnd FILL
X_8413_ _8413_/A _8413_/B _8413_/C _8413_/Y vdd gnd OAI21X1
XFILL_0__11479_ vdd gnd FILL
X_9393_ _9393_/A _9393_/B _9393_/C _9393_/Y vdd gnd NAND3X1
XFILL_2__12039_ vdd gnd FILL
XFILL_0__13218_ vdd gnd FILL
XFILL_1__12769_ vdd gnd FILL
X_8344_ _8344_/A _8344_/B _8344_/Y vdd gnd NAND2X1
XFILL_0__7997_ vdd gnd FILL
XFILL_0__13149_ vdd gnd FILL
XFILL_0__9736_ vdd gnd FILL
X_8275_ _8275_/A _8275_/Y vdd gnd INVX1
XFILL_1__14439_ vdd gnd FILL
X_7226_ _7226_/A _7226_/B _7226_/C _7226_/Y vdd gnd OAI21X1
XFILL_1__8460_ vdd gnd FILL
XFILL_0__9667_ vdd gnd FILL
XFILL_1__7411_ vdd gnd FILL
XFILL_0__8618_ vdd gnd FILL
X_7157_ _7157_/A _7157_/Y vdd gnd INVX8
XFILL_1__8391_ vdd gnd FILL
XFILL_0__9598_ vdd gnd FILL
XFILL_1__7342_ vdd gnd FILL
XFILL_0__8549_ vdd gnd FILL
X_7088_ _7088_/A _7088_/B _7088_/C _7088_/Y vdd gnd OAI21X1
XFILL_1__7273_ vdd gnd FILL
XFILL_1__9012_ vdd gnd FILL
X_11660_ _11660_/D _11660_/CLK _11660_/Q vdd gnd DFFPOSX1
X_9729_ _9729_/A _9729_/B _9729_/C _9729_/Y vdd gnd OAI21X1
X_10611_ _10611_/A _10611_/Y vdd gnd INVX1
XFILL256950x169350 vdd gnd FILL
XFILL_1__9914_ vdd gnd FILL
X_11591_ _11591_/A _11591_/B _11591_/C _11591_/Y vdd gnd OAI21X1
X_13330_ _13330_/A _13330_/B _13330_/Y vdd gnd AND2X2
X_10542_ _10542_/A _10542_/B _10542_/Y vdd gnd NAND2X1
XFILL_1__9845_ vdd gnd FILL
X_13261_ _13261_/A _13261_/B _13261_/Y vdd gnd NOR2X1
X_10473_ _10473_/A _10473_/B _10473_/Y vdd gnd OR2X2
X_12212_ _12212_/A _12212_/B _12212_/C _12212_/Y vdd gnd NAND3X1
X_13192_ _13192_/A _13192_/Y vdd gnd INVX1
XFILL_2__7520_ vdd gnd FILL
XFILL_1__8727_ vdd gnd FILL
X_12143_ _12143_/A _12143_/B _12143_/C _12143_/Y vdd gnd NAND3X1
XFILL_2__7451_ vdd gnd FILL
XFILL_1__8658_ vdd gnd FILL
X_12074_ _12074_/A _12074_/B _12074_/C _12074_/Y vdd gnd OAI21X1
XFILL_1__7609_ vdd gnd FILL
XFILL257250x68550 vdd gnd FILL
XFILL_2__7382_ vdd gnd FILL
XFILL_1__8589_ vdd gnd FILL
X_11025_ _11025_/A _11025_/B _11025_/C _11025_/Y vdd gnd NAND3X1
XFILL_1__10120_ vdd gnd FILL
XFILL_0__10850_ vdd gnd FILL
XFILL_2__9052_ vdd gnd FILL
XFILL_2__11410_ vdd gnd FILL
XFILL_1__10051_ vdd gnd FILL
XFILL_0__10781_ vdd gnd FILL
X_12976_ _12976_/A _12976_/B _12976_/Y vdd gnd NOR2X1
XFILL_2__11341_ vdd gnd FILL
XFILL_0__12520_ vdd gnd FILL
X_14715_ _14715_/A _14715_/B _14715_/C _14715_/Y vdd gnd OAI21X1
X_11927_ _11927_/A _11927_/B _11927_/C _11927_/Y vdd gnd OAI21X1
XFILL_1__13810_ vdd gnd FILL
XFILL_2__11272_ vdd gnd FILL
XFILL_1__14790_ vdd gnd FILL
XFILL_0__12451_ vdd gnd FILL
X_14646_ _14646_/A _14646_/B _14646_/C _14646_/Y vdd gnd OAI21X1
X_11858_ _11858_/A _11858_/B _11858_/Y vdd gnd NAND2X1
XFILL_0__11402_ vdd gnd FILL
XFILL_1__13741_ vdd gnd FILL
XFILL_1__10953_ vdd gnd FILL
XFILL_0__12382_ vdd gnd FILL
X_10809_ _10809_/A _10809_/B _10809_/Y vdd gnd NAND2X1
X_14577_ _14577_/A _14577_/B _14577_/C _14577_/Y vdd gnd AOI21X1
X_11789_ _11789_/A _11789_/B _11789_/C _11789_/D _11789_/Y vdd gnd OAI22X1
XFILL_0__14121_ vdd gnd FILL
XFILL_1__13672_ vdd gnd FILL
XFILL_2__9885_ vdd gnd FILL
XFILL_0__11333_ vdd gnd FILL
XFILL_1__10884_ vdd gnd FILL
X_13528_ _13528_/A _13528_/Y vdd gnd INVX1
XFILL_1__12623_ vdd gnd FILL
XFILL_0__14052_ vdd gnd FILL
XFILL_0__11264_ vdd gnd FILL
XFILL_0__7851_ vdd gnd FILL
X_13459_ _13459_/D _13459_/CLK _13459_/Q vdd gnd DFFPOSX1
XFILL_2__13913_ vdd gnd FILL
XFILL_0__13003_ vdd gnd FILL
XFILL_0__10215_ vdd gnd FILL
XFILL_2__8767_ vdd gnd FILL
XFILL_0__11195_ vdd gnd FILL
XFILL_0__7782_ vdd gnd FILL
XFILL_2__7718_ vdd gnd FILL
XFILL_1__11505_ vdd gnd FILL
XFILL_0__10146_ vdd gnd FILL
XFILL_2__13844_ vdd gnd FILL
XFILL_1__12485_ vdd gnd FILL
XFILL_2__8698_ vdd gnd FILL
XFILL_0__9521_ vdd gnd FILL
X_8060_ _8060_/A _8060_/B _8060_/C _8060_/Y vdd gnd OAI21X1
XFILL_1__14224_ vdd gnd FILL
XFILL_1__11436_ vdd gnd FILL
XFILL_0__10077_ vdd gnd FILL
XFILL_2__13775_ vdd gnd FILL
XFILL_0__9452_ vdd gnd FILL
XFILL_2__12726_ vdd gnd FILL
XFILL_1__14155_ vdd gnd FILL
XFILL_0__13905_ vdd gnd FILL
XFILL_1__11367_ vdd gnd FILL
XFILL257550x219750 vdd gnd FILL
XFILL_0__8403_ vdd gnd FILL
XFILL_0__9383_ vdd gnd FILL
XFILL_1__13106_ vdd gnd FILL
XFILL_2__9319_ vdd gnd FILL
XFILL_2__12657_ vdd gnd FILL
XFILL_1__10318_ vdd gnd FILL
XFILL_1__14086_ vdd gnd FILL
XFILL_0__13836_ vdd gnd FILL
XFILL_1__11298_ vdd gnd FILL
XFILL_0__8334_ vdd gnd FILL
X_8962_ _8962_/A _8962_/Y vdd gnd INVX1
XFILL_1__13037_ vdd gnd FILL
XFILL_2__11608_ vdd gnd FILL
XFILL_1__10249_ vdd gnd FILL
XFILL_0__13767_ vdd gnd FILL
XFILL_0__10979_ vdd gnd FILL
X_7913_ _7913_/A _7913_/B _7913_/C _7913_/Y vdd gnd OAI21X1
XFILL_0__8265_ vdd gnd FILL
X_8893_ _8893_/D _8893_/CLK _8893_/Q vdd gnd DFFPOSX1
XFILL_2__11539_ vdd gnd FILL
XFILL_0__12718_ vdd gnd FILL
XFILL_0__7216_ vdd gnd FILL
XFILL_0__13698_ vdd gnd FILL
X_7844_ _7844_/A _7844_/B _7844_/C _7844_/Y vdd gnd OAI21X1
XFILL_0__8196_ vdd gnd FILL
XFILL_0__12649_ vdd gnd FILL
XFILL_0__7147_ vdd gnd FILL
XFILL_0_CLKBUF1_insert107 vdd gnd FILL
X_7775_ _7775_/A _7775_/B _7775_/Y vdd gnd NAND2X1
XFILL_1__13939_ vdd gnd FILL
X_9514_ _9514_/A _9514_/B _9514_/C _9514_/Y vdd gnd NAND3X1
XFILL_0__7078_ vdd gnd FILL
XFILL_0__14319_ vdd gnd FILL
X_9445_ _9445_/A _9445_/B _9445_/Y vdd gnd NAND2X1
XFILL_1__7891_ vdd gnd FILL
XFILL_1__9630_ vdd gnd FILL
X_9376_ _9376_/A _9376_/B _9376_/C _9376_/D _9376_/Y vdd gnd AOI22X1
X_8327_ _8327_/A _8327_/Y vdd gnd INVX1
XFILL_1__9561_ vdd gnd FILL
XFILL_0__9719_ vdd gnd FILL
XFILL_1__8512_ vdd gnd FILL
X_8258_ _8258_/A _8258_/B _8258_/C _8258_/Y vdd gnd NAND3X1
XFILL_1__9492_ vdd gnd FILL
X_7209_ _7209_/A _7209_/B _7209_/S _7209_/Y vdd gnd MUX2X1
XFILL_1__8443_ vdd gnd FILL
X_8189_ _8189_/A _8189_/B _8189_/C _8189_/Y vdd gnd OAI21X1
XFILL256950x144150 vdd gnd FILL
XFILL257550x129750 vdd gnd FILL
XFILL_1__8374_ vdd gnd FILL
XFILL_1__7325_ vdd gnd FILL
X_12830_ _12830_/A _12830_/Y vdd gnd INVX1
XFILL_1__7256_ vdd gnd FILL
X_12761_ _12761_/A _12761_/B _12761_/Y vdd gnd NOR2X1
XFILL_1__7187_ vdd gnd FILL
X_14500_ _14500_/D _14500_/CLK _14500_/Q vdd gnd DFFPOSX1
XFILL257550x172950 vdd gnd FILL
X_11712_ _11712_/A _11712_/B _11712_/C _11712_/Y vdd gnd OAI21X1
X_12692_ _12692_/A _12692_/B _12692_/C _12692_/Y vdd gnd OAI21X1
X_14431_ _14431_/A _14431_/B _14431_/C _14431_/Y vdd gnd NAND3X1
X_11643_ _11643_/D _11643_/CLK _11643_/Q vdd gnd DFFPOSX1
XFILL257250x43350 vdd gnd FILL
X_14362_ _14362_/A _14362_/B _14362_/C _14362_/Y vdd gnd OAI21X1
X_11574_ _11574_/A _11574_/B _11574_/Y vdd gnd NAND2X1
XFILL_2__9670_ vdd gnd FILL
X_10525_ _10525_/A _10525_/B _10525_/Y vdd gnd NAND2X1
X_13313_ _13313_/A _13313_/B _13313_/C _13313_/Y vdd gnd AOI21X1
X_14293_ _14293_/A _14293_/B _14293_/Y vdd gnd NAND2X1
X_13244_ _13244_/A _13244_/B _13244_/S _13244_/Y vdd gnd MUX2X1
X_10456_ _10456_/A _10456_/B _10456_/C _10456_/Y vdd gnd OAI21X1
XFILL_0__10000_ vdd gnd FILL
XFILL_2__10910_ vdd gnd FILL
XFILL_1__9759_ vdd gnd FILL
X_13175_ _13175_/A _13175_/B _13175_/C _13175_/D _13175_/Y vdd gnd OAI22X1
X_10387_ _10387_/A _10387_/B _10387_/Y vdd gnd NOR2X1
XFILL_2__7503_ vdd gnd FILL
XFILL_2__10841_ vdd gnd FILL
XFILL_1__12270_ vdd gnd FILL
X_12126_ _12126_/A _12126_/B _12126_/C _12126_/Y vdd gnd OAI21X1
XFILL_2__7434_ vdd gnd FILL
XFILL_1__11221_ vdd gnd FILL
XFILL_2__13560_ vdd gnd FILL
XFILL_2__10772_ vdd gnd FILL
XFILL_0__11951_ vdd gnd FILL
X_12057_ _12057_/A _12057_/B _12057_/C _12057_/Y vdd gnd OAI21X1
XFILL_2__7365_ vdd gnd FILL
XFILL_0_CLKBUF1_insert31 vdd gnd FILL
XFILL_0__10902_ vdd gnd FILL
XFILL_1__11152_ vdd gnd FILL
X_11008_ _11008_/A _11008_/B _11008_/C _11008_/Y vdd gnd NAND3X1
XFILL_0__14670_ vdd gnd FILL
XFILL_0_CLKBUF1_insert42 vdd gnd FILL
XFILL_0__11882_ vdd gnd FILL
XFILL_0_CLKBUF1_insert53 vdd gnd FILL
XFILL_0_CLKBUF1_insert64 vdd gnd FILL
XFILL_1__10103_ vdd gnd FILL
XFILL_0_CLKBUF1_insert75 vdd gnd FILL
XFILL_2__7296_ vdd gnd FILL
XFILL_0__13621_ vdd gnd FILL
XFILL_1__11083_ vdd gnd FILL
XFILL_0_CLKBUF1_insert86 vdd gnd FILL
XFILL_0__10833_ vdd gnd FILL
XFILL_0_CLKBUF1_insert97 vdd gnd FILL
XFILL_1__14911_ vdd gnd FILL
XFILL_1__10034_ vdd gnd FILL
XFILL_0__13552_ vdd gnd FILL
XFILL_0__8050_ vdd gnd FILL
XFILL_2_BUFX2_insert382 vdd gnd FILL
X_12959_ _12959_/A _12959_/B _12959_/Y vdd gnd NAND2X1
XFILL_0__12503_ vdd gnd FILL
XFILL_1__14842_ vdd gnd FILL
XFILL_1__14773_ vdd gnd FILL
XFILL_0__12434_ vdd gnd FILL
XFILL_1__11985_ vdd gnd FILL
X_14629_ _14629_/A _14629_/B _14629_/Y vdd gnd NOR2X1
X_7560_ _7560_/A _7560_/B _7560_/Y vdd gnd NOR2X1
XFILL_2__10206_ vdd gnd FILL
XFILL_2__11186_ vdd gnd FILL
XFILL_1__10936_ vdd gnd FILL
XFILL_1__13724_ vdd gnd FILL
XFILL_0__12365_ vdd gnd FILL
XFILL_0__8952_ vdd gnd FILL
X_7491_ _7491_/A _7491_/B _7491_/C _7491_/Y vdd gnd OAI21X1
XFILL_2__10137_ vdd gnd FILL
XFILL_0__14104_ vdd gnd FILL
XBUFX2_insert370 BUFX2_insert370/A BUFX2_insert370/Y vdd gnd BUFX2
XFILL_0__11316_ vdd gnd FILL
XFILL_1__13655_ vdd gnd FILL
XBUFX2_insert381 BUFX2_insert381/A BUFX2_insert381/Y vdd gnd BUFX2
XFILL_1__10867_ vdd gnd FILL
X_9230_ _9230_/A _9230_/B _9230_/C _9230_/Y vdd gnd NAND3X1
XFILL_0__7903_ vdd gnd FILL
XFILL_0__12296_ vdd gnd FILL
XFILL_0__14035_ vdd gnd FILL
XFILL_0__11247_ vdd gnd FILL
XFILL_1__13586_ vdd gnd FILL
XFILL_1__10798_ vdd gnd FILL
XFILL_0__7834_ vdd gnd FILL
X_9161_ _9161_/A _9161_/B _9161_/Y vdd gnd NAND2X1
X_8112_ _8112_/A _8112_/B _8112_/S _8112_/Y vdd gnd MUX2X1
XFILL_0__11178_ vdd gnd FILL
X_9092_ _9092_/A _9092_/B _9092_/C _9092_/D _9092_/Y vdd gnd AOI22X1
XFILL_0__7765_ vdd gnd FILL
XFILL_2__13827_ vdd gnd FILL
XFILL_0__10129_ vdd gnd FILL
XFILL_1__12468_ vdd gnd FILL
XFILL_0__9504_ vdd gnd FILL
X_8043_ _8043_/A _8043_/B _8043_/C _8043_/Y vdd gnd OAI21X1
XFILL_0__7696_ vdd gnd FILL
XFILL_1__11419_ vdd gnd FILL
XFILL_2__13758_ vdd gnd FILL
XFILL_1__12399_ vdd gnd FILL
XFILL_0__9435_ vdd gnd FILL
XFILL_1__14138_ vdd gnd FILL
XFILL_0__14868_ vdd gnd FILL
XFILL_2__13689_ vdd gnd FILL
XFILL_0__9366_ vdd gnd FILL
X_9994_ _9994_/A _9994_/Y vdd gnd INVX1
XFILL_1__14069_ vdd gnd FILL
XFILL_0__13819_ vdd gnd FILL
XFILL_1__7110_ vdd gnd FILL
XFILL_0__14799_ vdd gnd FILL
XFILL_0__8317_ vdd gnd FILL
XFILL_0__9297_ vdd gnd FILL
XFILL_1__8090_ vdd gnd FILL
X_8945_ _8945_/A _8945_/B _8945_/C _8945_/Y vdd gnd OAI21X1
XFILL_0__8248_ vdd gnd FILL
X_8876_ _8876_/D _8876_/CLK _8876_/Q vdd gnd DFFPOSX1
X_7827_ _7827_/A _7827_/B _7827_/C _7827_/Y vdd gnd OAI21X1
XFILL_0__8179_ vdd gnd FILL
X_7758_ _7758_/A _7758_/B _7758_/Y vdd gnd NOR2X1
XFILL_1__8992_ vdd gnd FILL
XFILL257550x104550 vdd gnd FILL
X_7689_ _7689_/A _7689_/B _7689_/Y vdd gnd NAND2X1
X_9428_ _9428_/A _9428_/B _9428_/C _9428_/Y vdd gnd OAI21X1
XFILL_1__7874_ vdd gnd FILL
X_10310_ _10310_/A _10310_/B _10310_/C _10310_/Y vdd gnd OAI21X1
XFILL_1__9613_ vdd gnd FILL
X_11290_ _11290_/A _11290_/B _11290_/C _11290_/Y vdd gnd OAI21X1
X_9359_ _9359_/A _9359_/B _9359_/C _9359_/Y vdd gnd OAI21X1
X_10241_ _10241_/A _10241_/B _10241_/C _10241_/Y vdd gnd OAI21X1
XFILL_1__9544_ vdd gnd FILL
X_10172_ _10172_/A _10172_/B _10172_/Y vdd gnd NAND2X1
XFILL_1__9475_ vdd gnd FILL
XFILL_1__8426_ vdd gnd FILL
X_13931_ _13931_/A _13931_/B _13931_/Y vdd gnd OR2X2
XFILL_2__7150_ vdd gnd FILL
XFILL_1__8357_ vdd gnd FILL
X_13862_ _13862_/A _13862_/B _13862_/Y vdd gnd NAND2X1
XFILL_1__7308_ vdd gnd FILL
XFILL_2__7081_ vdd gnd FILL
XFILL_1__8288_ vdd gnd FILL
X_12813_ _12813_/A _12813_/B _12813_/C _12813_/Y vdd gnd AOI21X1
XFILL_1_BUFX2_insert301 vdd gnd FILL
XFILL_1__7239_ vdd gnd FILL
XFILL_1_BUFX2_insert312 vdd gnd FILL
X_13793_ _13793_/A _13793_/B _13793_/C _13793_/Y vdd gnd NOR3X1
XFILL_1_BUFX2_insert323 vdd gnd FILL
XFILL_1_BUFX2_insert334 vdd gnd FILL
XFILL_1_BUFX2_insert345 vdd gnd FILL
X_12744_ _12744_/A _12744_/B _12744_/Y vdd gnd NAND2X1
XFILL_1_BUFX2_insert356 vdd gnd FILL
XFILL_1_BUFX2_insert367 vdd gnd FILL
XFILL_0__10480_ vdd gnd FILL
XFILL_1_BUFX2_insert378 vdd gnd FILL
X_12675_ _12675_/A _12675_/B _12675_/Y vdd gnd NAND2X1
XFILL_1__11770_ vdd gnd FILL
X_14414_ _14414_/A _14414_/B _14414_/C _14414_/Y vdd gnd NAND3X1
X_11626_ _11626_/D _11626_/CLK _11626_/Q vdd gnd DFFPOSX1
XFILL_2__9722_ vdd gnd FILL
XFILL_0__12150_ vdd gnd FILL
X_14345_ _14345_/A _14345_/B _14345_/Y vdd gnd NAND2X1
X_11557_ _11557_/A _11557_/B _11557_/C _11557_/Y vdd gnd OAI21X1
XFILL_2__9653_ vdd gnd FILL
XFILL_0__11101_ vdd gnd FILL
XFILL_1__10652_ vdd gnd FILL
XFILL_0__12081_ vdd gnd FILL
XFILL_2__12991_ vdd gnd FILL
X_10508_ _10508_/A _10508_/B _10508_/Y vdd gnd NAND2X1
X_14276_ _14276_/A _14276_/B _14276_/C _14276_/Y vdd gnd OAI21X1
X_11488_ _11488_/A _11488_/B _11488_/C _11488_/Y vdd gnd AOI21X1
XFILL_0__11032_ vdd gnd FILL
XFILL_2__9584_ vdd gnd FILL
XFILL_1__13371_ vdd gnd FILL
XFILL_1__10583_ vdd gnd FILL
X_10439_ _10439_/A _10439_/B _10439_/Y vdd gnd AND2X2
X_13227_ _13227_/A _13227_/B _13227_/Y vdd gnd NOR2X1
XFILL_1__12322_ vdd gnd FILL
XFILL_0__7550_ vdd gnd FILL
X_13158_ _13158_/A _13158_/B _13158_/C _13158_/Y vdd gnd AOI21X1
XFILL_1__12253_ vdd gnd FILL
XFILL_2__10824_ vdd gnd FILL
X_12109_ _12109_/A _12109_/B _12109_/C _12109_/Y vdd gnd OAI21X1
XFILL_0__12983_ vdd gnd FILL
X_13089_ _13089_/A _13089_/B _13089_/C _13089_/Y vdd gnd OAI21X1
XFILL_0__7481_ vdd gnd FILL
XFILL_2__7417_ vdd gnd FILL
XFILL_1__11204_ vdd gnd FILL
XFILL_0__14722_ vdd gnd FILL
XFILL_0__11934_ vdd gnd FILL
XFILL_1__12184_ vdd gnd FILL
XFILL_0__9220_ vdd gnd FILL
XFILL_2__7348_ vdd gnd FILL
XFILL_1__11135_ vdd gnd FILL
XFILL_0__14653_ vdd gnd FILL
XFILL_0__9151_ vdd gnd FILL
XFILL_0__11865_ vdd gnd FILL
XFILL_2__12425_ vdd gnd FILL
XFILL_0__13604_ vdd gnd FILL
XFILL_2__7279_ vdd gnd FILL
XFILL_0__8102_ vdd gnd FILL
XFILL_0__10816_ vdd gnd FILL
XFILL_1__11066_ vdd gnd FILL
XFILL_0__14584_ vdd gnd FILL
XFILL_0__9082_ vdd gnd FILL
X_8730_ _8730_/A _8730_/B _8730_/Y vdd gnd NOR2X1
XFILL_0__11796_ vdd gnd FILL
XFILL_1__10017_ vdd gnd FILL
XFILL_2__12356_ vdd gnd FILL
XFILL_0__13535_ vdd gnd FILL
XFILL_0__8033_ vdd gnd FILL
X_8661_ _8661_/A _8661_/Y vdd gnd INVX1
XFILL_1__14825_ vdd gnd FILL
X_7612_ _7612_/A _7612_/B _7612_/C _7612_/Y vdd gnd NAND3X1
XFILL_0__10678_ vdd gnd FILL
X_8592_ _8592_/A _8592_/B _8592_/Y vdd gnd NOR2X1
XFILL_0__12417_ vdd gnd FILL
XFILL_1__14756_ vdd gnd FILL
XFILL_1__11968_ vdd gnd FILL
XFILL_0__13397_ vdd gnd FILL
X_7543_ _7543_/A _7543_/B _7543_/Y vdd gnd OR2X2
XFILL_0__9984_ vdd gnd FILL
XFILL_1__10919_ vdd gnd FILL
XFILL_1__13707_ vdd gnd FILL
XFILL_0__12348_ vdd gnd FILL
XFILL_1__14687_ vdd gnd FILL
XFILL_1__11899_ vdd gnd FILL
XFILL_0__8935_ vdd gnd FILL
X_7474_ _7474_/A _7474_/B _7474_/S _7474_/Y vdd gnd MUX2X1
XFILL_1__13638_ vdd gnd FILL
X_9213_ _9213_/A _9213_/B _9213_/C _9213_/Y vdd gnd NAND3X1
XFILL_0__12279_ vdd gnd FILL
XFILL_0__14018_ vdd gnd FILL
XFILL_1__13569_ vdd gnd FILL
X_9144_ _9144_/A _9144_/B _9144_/C _9144_/Y vdd gnd OAI21X1
XFILL_0__7817_ vdd gnd FILL
XFILL_1__7590_ vdd gnd FILL
XFILL_0__8797_ vdd gnd FILL
X_9075_ _9075_/A _9075_/B _9075_/C _9075_/Y vdd gnd AOI21X1
XFILL_0__7748_ vdd gnd FILL
X_8026_ _8026_/A _8026_/B _8026_/C _8026_/Y vdd gnd OAI21X1
XFILL_1__9260_ vdd gnd FILL
XFILL_0__7679_ vdd gnd FILL
XFILL_0__9418_ vdd gnd FILL
XFILL_1__8211_ vdd gnd FILL
XFILL_1__9191_ vdd gnd FILL
XFILL_1__8142_ vdd gnd FILL
XFILL_0__9349_ vdd gnd FILL
X_9977_ _9977_/A _9977_/B _9977_/Y vdd gnd NAND2X1
XFILL_1__8073_ vdd gnd FILL
X_8928_ _8928_/A _8928_/Y vdd gnd INVX2
X_10790_ _10790_/A _10790_/B _10790_/C _10790_/D _10790_/Y vdd gnd AOI22X1
X_8859_ _8859_/D _8859_/CLK _8859_/Q vdd gnd DFFPOSX1
XFILL_0_BUFX2_insert308 vdd gnd FILL
XFILL_0_BUFX2_insert319 vdd gnd FILL
X_12460_ _12460_/A _12460_/B _12460_/Y vdd gnd OR2X2
XFILL_1__8975_ vdd gnd FILL
X_11411_ _11411_/A _11411_/B _11411_/Y vdd gnd NAND2X1
X_12391_ _12391_/A _12391_/B _12391_/C _12391_/Y vdd gnd OAI21X1
X_11342_ _11342_/A _11342_/B _11342_/Y vdd gnd OR2X2
X_14130_ _14130_/A _14130_/B _14130_/C _14130_/Y vdd gnd OAI21X1
XFILL_1__7857_ vdd gnd FILL
X_14061_ _14061_/A _14061_/B _14061_/C _14061_/Y vdd gnd NAND3X1
X_11273_ _11273_/A _11273_/B _11273_/C _11273_/Y vdd gnd NAND3X1
XFILL_1__7788_ vdd gnd FILL
X_10224_ _10224_/A _10224_/B _10224_/Y vdd gnd NAND2X1
X_13012_ _13012_/A _13012_/B _13012_/S _13012_/Y vdd gnd MUX2X1
XFILL_1__9527_ vdd gnd FILL
X_10155_ _10155_/A _10155_/Y vdd gnd INVX1
XFILL_1__9458_ vdd gnd FILL
X_10086_ _10086_/A _10086_/B _10086_/C _10086_/Y vdd gnd AOI21X1
XFILL_1__8409_ vdd gnd FILL
XFILL_1__9389_ vdd gnd FILL
X_13914_ _13914_/A _13914_/B _13914_/C _13914_/Y vdd gnd NAND3X1
X_14894_ _14894_/D _14894_/CLK _14894_/Q vdd gnd DFFPOSX1
XFILL_2__12210_ vdd gnd FILL
X_13845_ _13845_/A _13845_/B _13845_/C _13845_/Y vdd gnd OAI21X1
XFILL_0__10601_ vdd gnd FILL
XFILL_1__12940_ vdd gnd FILL
XFILL_1_BUFX2_insert120 vdd gnd FILL
XFILL_0__11581_ vdd gnd FILL
XFILL_1_BUFX2_insert131 vdd gnd FILL
XFILL_1_BUFX2_insert142 vdd gnd FILL
XFILL_2__12141_ vdd gnd FILL
X_13776_ _13776_/A _13776_/B _13776_/C _13776_/Y vdd gnd NAND3X1
X_10988_ _10988_/A _10988_/B _10988_/C _10988_/Y vdd gnd AOI21X1
XFILL_0__13320_ vdd gnd FILL
XFILL_0__10532_ vdd gnd FILL
XFILL_1_BUFX2_insert153 vdd gnd FILL
XFILL_1__12871_ vdd gnd FILL
XFILL_1_BUFX2_insert164 vdd gnd FILL
XFILL_1_BUFX2_insert175 vdd gnd FILL
X_12727_ _12727_/A _12727_/B _12727_/S _12727_/Y vdd gnd MUX2X1
XFILL_1_BUFX2_insert186 vdd gnd FILL
XFILL_1__14610_ vdd gnd FILL
XFILL_1_BUFX2_insert197 vdd gnd FILL
XFILL_1__11822_ vdd gnd FILL
XFILL_2__12072_ vdd gnd FILL
XFILL_0__13251_ vdd gnd FILL
XFILL_0__10463_ vdd gnd FILL
X_12658_ _12658_/A _12658_/B _12658_/C _12658_/D _12658_/Y vdd gnd AOI22X1
XFILL_0__12202_ vdd gnd FILL
XFILL_1__11753_ vdd gnd FILL
XFILL_0__13182_ vdd gnd FILL
XFILL_0__10394_ vdd gnd FILL
X_11609_ _11609_/A _11609_/B _11609_/C _11609_/Y vdd gnd OAI21X1
XFILL_2__9705_ vdd gnd FILL
X_12589_ _12589_/D _12589_/CLK _12589_/Q vdd gnd DFFPOSX1
XFILL_1__14472_ vdd gnd FILL
XFILL_0__12133_ vdd gnd FILL
XFILL_0__8720_ vdd gnd FILL
X_14328_ _14328_/A _14328_/B _14328_/C _14328_/Y vdd gnd NAND3X1
XFILL_2__9636_ vdd gnd FILL
XFILL_1__13423_ vdd gnd FILL
XFILL_1__10635_ vdd gnd FILL
XFILL_0__12064_ vdd gnd FILL
XFILL_2__12974_ vdd gnd FILL
XFILL_0__8651_ vdd gnd FILL
X_14259_ _14259_/A _14259_/B _14259_/C _14259_/Y vdd gnd OAI21X1
X_7190_ _7190_/A _7190_/B _7190_/S _7190_/Y vdd gnd MUX2X1
XFILL_2__14713_ vdd gnd FILL
XFILL_0__11015_ vdd gnd FILL
XFILL_2__9567_ vdd gnd FILL
XFILL_1__13354_ vdd gnd FILL
XFILL_1__10566_ vdd gnd FILL
XFILL_0__7602_ vdd gnd FILL
XFILL_0__8582_ vdd gnd FILL
XFILL_1__12305_ vdd gnd FILL
XFILL_2__9498_ vdd gnd FILL
XFILL_1__13285_ vdd gnd FILL
XFILL_1__10497_ vdd gnd FILL
XFILL_0__7533_ vdd gnd FILL
XFILL_1__12236_ vdd gnd FILL
XFILL_0__12966_ vdd gnd FILL
X_9900_ _9900_/A _9900_/B _9900_/C _9900_/D _9900_/Y vdd gnd AOI22X1
XFILL_0__7464_ vdd gnd FILL
XFILL_0__14705_ vdd gnd FILL
XFILL_0__11917_ vdd gnd FILL
XFILL_1__12167_ vdd gnd FILL
XFILL_0__9203_ vdd gnd FILL
XFILL_0__12897_ vdd gnd FILL
XFILL_0__7395_ vdd gnd FILL
X_9831_ _9831_/D _9831_/CLK _9831_/Q vdd gnd DFFPOSX1
XFILL_1__11118_ vdd gnd FILL
XFILL_0__14636_ vdd gnd FILL
XFILL_0__11848_ vdd gnd FILL
XFILL_1__12098_ vdd gnd FILL
XFILL_0__9134_ vdd gnd FILL
X_9762_ _9762_/A _9762_/B _9762_/Y vdd gnd NAND2X1
XFILL_2__12408_ vdd gnd FILL
XFILL_1__11049_ vdd gnd FILL
XFILL_0__14567_ vdd gnd FILL
XFILL_0__11779_ vdd gnd FILL
XFILL_0__9065_ vdd gnd FILL
X_8713_ _8713_/A _8713_/B _8713_/Y vdd gnd NAND2X1
X_9693_ _9693_/A _9693_/B _9693_/C _9693_/Y vdd gnd OAI21X1
XFILL_2__12339_ vdd gnd FILL
XFILL_0__13518_ vdd gnd FILL
XFILL_0__8016_ vdd gnd FILL
XFILL_0__14498_ vdd gnd FILL
X_8644_ _8644_/A _8644_/B _8644_/C _8644_/D _8644_/Y vdd gnd OAI22X1
XFILL_1__14808_ vdd gnd FILL
X_8575_ _8575_/A _8575_/B _8575_/Y vdd gnd AND2X2
XFILL_2__14009_ vdd gnd FILL
XFILL_1__14739_ vdd gnd FILL
X_7526_ _7526_/A _7526_/B _7526_/Y vdd gnd NAND2X1
XFILL_0__9967_ vdd gnd FILL
XFILL_1__8760_ vdd gnd FILL
XFILL_1__7711_ vdd gnd FILL
X_7457_ _7457_/A _7457_/B _7457_/Y vdd gnd NAND2X1
XFILL_0__9898_ vdd gnd FILL
XFILL_1__8691_ vdd gnd FILL
XFILL_1__7642_ vdd gnd FILL
X_7388_ _7388_/A _7388_/B _7388_/C _7388_/Y vdd gnd NAND3X1
X_9127_ _9127_/A _9127_/B _9127_/C _9127_/Y vdd gnd OAI21X1
XFILL_1__7573_ vdd gnd FILL
XFILL_1__9312_ vdd gnd FILL
X_9058_ _9058_/A _9058_/B _9058_/S _9058_/Y vdd gnd MUX2X1
X_8009_ _8009_/A _8009_/B _8009_/C _8009_/D _8009_/Y vdd gnd AOI22X1
XFILL_1__9243_ vdd gnd FILL
X_11960_ _11960_/A _11960_/B _11960_/Y vdd gnd NAND2X1
XFILL_1__9174_ vdd gnd FILL
X_10911_ _10911_/A _10911_/B _10911_/C _10911_/Y vdd gnd AOI21X1
XFILL_1__8125_ vdd gnd FILL
X_11891_ _11891_/A _11891_/B _11891_/C _11891_/Y vdd gnd NAND3X1
X_13630_ _13630_/A _13630_/B _13630_/Y vdd gnd NAND2X1
X_10842_ _10842_/A _10842_/B _10842_/C _10842_/Y vdd gnd OAI21X1
XFILL_1__8056_ vdd gnd FILL
X_13561_ _13561_/A _13561_/B _13561_/S _13561_/Y vdd gnd MUX2X1
X_10773_ _10773_/A _10773_/Y vdd gnd INVX4
X_12512_ _12512_/A _12512_/B _12512_/Y vdd gnd NAND2X1
XFILL_0_BUFX2_insert116 vdd gnd FILL
XFILL_0_BUFX2_insert127 vdd gnd FILL
XFILL_0_BUFX2_insert138 vdd gnd FILL
XFILL_2__7820_ vdd gnd FILL
X_13492_ _13492_/D _13492_/CLK _13492_/Q vdd gnd DFFPOSX1
XFILL_0_BUFX2_insert149 vdd gnd FILL
X_12443_ _12443_/A _12443_/B _12443_/Y vdd gnd NAND2X1
XFILL_1__8958_ vdd gnd FILL
XFILL_2__7751_ vdd gnd FILL
XFILL_1__7909_ vdd gnd FILL
X_12374_ _12374_/A _12374_/B _12374_/Y vdd gnd OR2X2
XFILL_2__7682_ vdd gnd FILL
X_14113_ _14113_/A _14113_/B _14113_/Y vdd gnd NAND2X1
X_11325_ _11325_/A _11325_/B _11325_/Y vdd gnd NAND2X1
XFILL_1_CLKBUF1_insert385 vdd gnd FILL
XFILL_1__10420_ vdd gnd FILL
X_14044_ _14044_/A _14044_/B _14044_/C _14044_/Y vdd gnd AOI21X1
X_11256_ _11256_/A _11256_/B _11256_/Y vdd gnd NOR2X1
XFILL_2__11710_ vdd gnd FILL
XFILL_1__10351_ vdd gnd FILL
X_10207_ _10207_/A _10207_/Y vdd gnd INVX1
X_11187_ _11187_/A _11187_/B _11187_/C _11187_/Y vdd gnd OAI21X1
XFILL_2__8303_ vdd gnd FILL
XFILL_0__12820_ vdd gnd FILL
XFILL_1__13070_ vdd gnd FILL
XFILL_1__10282_ vdd gnd FILL
X_10138_ _10138_/A _10138_/B _10138_/Y vdd gnd AND2X2
XFILL_1__12021_ vdd gnd FILL
XFILL_2__8234_ vdd gnd FILL
XFILL_0__12751_ vdd gnd FILL
X_10069_ _10069_/A _10069_/B _10069_/C _10069_/Y vdd gnd OAI21X1
XFILL_2__10523_ vdd gnd FILL
XFILL_2__8165_ vdd gnd FILL
XFILL_0__11702_ vdd gnd FILL
XFILL_0__12682_ vdd gnd FILL
XFILL_0__7180_ vdd gnd FILL
X_14877_ _14877_/D _14877_/CLK _14877_/Q vdd gnd DFFPOSX1
XFILL_0__14421_ vdd gnd FILL
XFILL_1__13972_ vdd gnd FILL
X_13828_ _13828_/A _13828_/B _13828_/C _13828_/Y vdd gnd OAI21X1
XFILL_0__14352_ vdd gnd FILL
XFILL_1__12923_ vdd gnd FILL
XFILL_0__11564_ vdd gnd FILL
X_13759_ _13759_/A _13759_/B _13759_/C _13759_/Y vdd gnd OAI21X1
XFILL_2__12124_ vdd gnd FILL
XFILL_0__13303_ vdd gnd FILL
XFILL_0__10515_ vdd gnd FILL
XFILL_0__14283_ vdd gnd FILL
XFILL_1__12854_ vdd gnd FILL
XFILL_0__11495_ vdd gnd FILL
XFILL_2__12055_ vdd gnd FILL
XFILL_1__11805_ vdd gnd FILL
XFILL_0__13234_ vdd gnd FILL
XFILL_0__10446_ vdd gnd FILL
XFILL_2__8998_ vdd gnd FILL
XFILL_1__12785_ vdd gnd FILL
X_8360_ _8360_/A _8360_/B _8360_/Y vdd gnd NAND2X1
XFILL_0__13165_ vdd gnd FILL
XFILL_1__11736_ vdd gnd FILL
XFILL_0__10377_ vdd gnd FILL
X_7311_ _7311_/A _7311_/B _7311_/Y vdd gnd NAND2X1
XFILL_0__9752_ vdd gnd FILL
X_8291_ _8291_/A _8291_/Y vdd gnd INVX1
XFILL_0__12116_ vdd gnd FILL
XFILL_1__14455_ vdd gnd FILL
XFILL_0__13096_ vdd gnd FILL
XFILL_0__8703_ vdd gnd FILL
X_7242_ _7242_/A _7242_/B _7242_/Y vdd gnd NOR2X1
XFILL_0__9683_ vdd gnd FILL
XFILL_1__10618_ vdd gnd FILL
XFILL_1__13406_ vdd gnd FILL
XFILL_1__14386_ vdd gnd FILL
XFILL_0__12047_ vdd gnd FILL
XFILL_2__12957_ vdd gnd FILL
XFILL_1__11598_ vdd gnd FILL
XFILL_0__8634_ vdd gnd FILL
X_7173_ _7173_/A _7173_/B _7173_/Y vdd gnd NAND2X1
XFILL_2__11908_ vdd gnd FILL
XFILL_1__10549_ vdd gnd FILL
XFILL_1__13337_ vdd gnd FILL
XFILL_2__12888_ vdd gnd FILL
XFILL_0__8565_ vdd gnd FILL
XFILL_2__14627_ vdd gnd FILL
XFILL_1__13268_ vdd gnd FILL
XCLKBUF1_insert384 CLKBUF1_insert384/A CLKBUF1_insert384/Y vdd gnd CLKBUF1
XFILL_0__7516_ vdd gnd FILL
XFILL_0__13998_ vdd gnd FILL
XFILL_0__8496_ vdd gnd FILL
XFILL_1__12219_ vdd gnd FILL
XFILL_2__14558_ vdd gnd FILL
XFILL_1__13199_ vdd gnd FILL
XFILL_0__12949_ vdd gnd FILL
XFILL_0__7447_ vdd gnd FILL
X_9814_ _9814_/D _9814_/CLK _9814_/Q vdd gnd DFFPOSX1
XFILL_0__7378_ vdd gnd FILL
XFILL_0__14619_ vdd gnd FILL
XFILL_0__9117_ vdd gnd FILL
X_9745_ _9745_/A _9745_/Y vdd gnd INVX1
XFILL_0__9048_ vdd gnd FILL
XFILL_1__9930_ vdd gnd FILL
X_9676_ _9676_/A _9676_/B _9676_/C _9676_/Y vdd gnd OAI21X1
XFILL_1__9861_ vdd gnd FILL
X_8627_ _8627_/A _8627_/B _8627_/Y vdd gnd NAND2X1
XFILL_1__8812_ vdd gnd FILL
X_8558_ _8558_/A _8558_/B _8558_/C _8558_/Y vdd gnd OAI21X1
X_7509_ _7509_/A _7509_/Y vdd gnd INVX1
XFILL_1__8743_ vdd gnd FILL
X_8489_ _8489_/A _8489_/Y vdd gnd INVX1
XFILL_1__8674_ vdd gnd FILL
X_11110_ _11110_/A _11110_/B _11110_/C _11110_/Y vdd gnd OAI21X1
X_12090_ _12090_/A _12090_/B _12090_/Y vdd gnd NAND2X1
XFILL_1__7625_ vdd gnd FILL
X_11041_ _11041_/A _11041_/B _11041_/C _11041_/Y vdd gnd OAI21X1
XFILL_1__7556_ vdd gnd FILL
XFILL_1__7487_ vdd gnd FILL
X_14800_ _14800_/A _14800_/B _14800_/C _14800_/Y vdd gnd OAI21X1
XFILL_1__9226_ vdd gnd FILL
XFILL257250x183750 vdd gnd FILL
X_12992_ _12992_/A _12992_/B _12992_/C _12992_/Y vdd gnd OAI21X1
X_14731_ _14731_/A _14731_/B _14731_/C _14731_/Y vdd gnd AOI21X1
X_11943_ _11943_/A _11943_/B _11943_/Y vdd gnd AND2X2
XFILL_1__9157_ vdd gnd FILL
X_14662_ _14662_/A _14662_/B _14662_/Y vdd gnd NAND2X1
XFILL_1__8108_ vdd gnd FILL
X_11874_ _11874_/A _11874_/B _11874_/C _11874_/Y vdd gnd AOI21X1
XFILL_1__9088_ vdd gnd FILL
X_13613_ _13613_/A _13613_/B _13613_/Y vdd gnd AND2X2
X_10825_ _10825_/A _10825_/B _10825_/C _10825_/Y vdd gnd OAI21X1
X_14593_ _14593_/A _14593_/Y vdd gnd INVX8
XFILL_2__8921_ vdd gnd FILL
XFILL_1__8039_ vdd gnd FILL
XFILL_2__10170_ vdd gnd FILL
X_13544_ _13544_/A _13544_/Y vdd gnd INVX1
X_10756_ _10756_/D _10756_/CLK _10756_/Q vdd gnd DFFPOSX1
XFILL_0__10300_ vdd gnd FILL
XFILL_0__11280_ vdd gnd FILL
XFILL_2__7803_ vdd gnd FILL
X_13475_ _13475_/D _13475_/CLK _13475_/Q vdd gnd DFFPOSX1
X_10687_ _10687_/A _10687_/B _10687_/C _10687_/Y vdd gnd OAI21X1
XFILL_0__10231_ vdd gnd FILL
X_12426_ _12426_/A _12426_/B _12426_/Y vdd gnd NOR2X1
XFILL_2__7734_ vdd gnd FILL
XFILL_1__11521_ vdd gnd FILL
XFILL_0__10162_ vdd gnd FILL
X_12357_ _12357_/A _12357_/Y vdd gnd INVX1
XFILL_1__14240_ vdd gnd FILL
XFILL_2__7665_ vdd gnd FILL
XFILL_1__11452_ vdd gnd FILL
XFILL_0__10093_ vdd gnd FILL
X_11308_ _11308_/A _11308_/B _11308_/C _11308_/Y vdd gnd NAND3X1
XFILL_1__10403_ vdd gnd FILL
XFILL_2_BUFX2_insert3 vdd gnd FILL
X_12288_ _12288_/A _12288_/B _12288_/Y vdd gnd NOR2X1
XFILL_2__7596_ vdd gnd FILL
XFILL_1__11383_ vdd gnd FILL
XFILL_0__13921_ vdd gnd FILL
X_14027_ _14027_/A _14027_/B _14027_/Y vdd gnd NAND2X1
X_11239_ _11239_/A _11239_/B _11239_/Y vdd gnd OR2X2
XFILL_1__13122_ vdd gnd FILL
XFILL_1__10334_ vdd gnd FILL
XFILL_0__13852_ vdd gnd FILL
XFILL_0__8350_ vdd gnd FILL
XFILL_1__13053_ vdd gnd FILL
XFILL_1__10265_ vdd gnd FILL
XFILL_0__12803_ vdd gnd FILL
XFILL_0__7301_ vdd gnd FILL
XFILL_0__13783_ vdd gnd FILL
XFILL_0__10995_ vdd gnd FILL
XFILL_1__12004_ vdd gnd FILL
XFILL_0__8281_ vdd gnd FILL
XFILL_2__8217_ vdd gnd FILL
XFILL_0__12734_ vdd gnd FILL
XFILL_1__10196_ vdd gnd FILL
XFILL_0__7232_ vdd gnd FILL
X_7860_ _7860_/A _7860_/B _7860_/Y vdd gnd NAND2X1
XFILL_2__10506_ vdd gnd FILL
XFILL_2__8148_ vdd gnd FILL
XFILL_0__12665_ vdd gnd FILL
XFILL_0__7163_ vdd gnd FILL
X_7791_ _7791_/A _7791_/B _7791_/Y vdd gnd OR2X2
XFILL_2__10437_ vdd gnd FILL
XFILL_0__14404_ vdd gnd FILL
XFILL_2__8079_ vdd gnd FILL
XFILL_1__13955_ vdd gnd FILL
X_9530_ _9530_/A _9530_/B _9530_/Y vdd gnd AND2X2
XFILL_0__7094_ vdd gnd FILL
XFILL_1__12906_ vdd gnd FILL
XFILL_2__10368_ vdd gnd FILL
XFILL_0__14335_ vdd gnd FILL
XFILL_0__11547_ vdd gnd FILL
XFILL_1__13886_ vdd gnd FILL
X_9461_ _9461_/A _9461_/B _9461_/Y vdd gnd NAND2X1
XFILL_2__10299_ vdd gnd FILL
XFILL_0__14266_ vdd gnd FILL
XFILL_1__12837_ vdd gnd FILL
XFILL_0__11478_ vdd gnd FILL
X_8412_ _8412_/A _8412_/B _8412_/Y vdd gnd NAND2X1
X_9392_ _9392_/A _9392_/B _9392_/C _9392_/Y vdd gnd OAI21X1
XFILL_0__13217_ vdd gnd FILL
XFILL_0__10429_ vdd gnd FILL
XFILL_1__12768_ vdd gnd FILL
X_8343_ _8343_/A _8343_/Y vdd gnd INVX1
XFILL_0__7996_ vdd gnd FILL
XFILL_0__13148_ vdd gnd FILL
XFILL_1__11719_ vdd gnd FILL
XFILL_0__9735_ vdd gnd FILL
XFILL_1__12699_ vdd gnd FILL
X_8274_ _8274_/A _8274_/B _8274_/C _8274_/Y vdd gnd OAI21X1
XFILL_1__14438_ vdd gnd FILL
XFILL_0__13079_ vdd gnd FILL
XFILL_2__13989_ vdd gnd FILL
X_7225_ _7225_/A _7225_/Y vdd gnd INVX1
XFILL_0__9666_ vdd gnd FILL
XFILL_1__14369_ vdd gnd FILL
XFILL_1__7410_ vdd gnd FILL
XFILL_0__8617_ vdd gnd FILL
X_7156_ _7156_/A _7156_/B _7156_/C _7156_/Y vdd gnd OAI21X1
XFILL_0__9597_ vdd gnd FILL
XFILL_1__8390_ vdd gnd FILL
XFILL_1__7341_ vdd gnd FILL
XFILL_0__8548_ vdd gnd FILL
X_7087_ _7087_/A _7087_/Y vdd gnd INVX1
XFILL_1__7272_ vdd gnd FILL
XFILL_0__8479_ vdd gnd FILL
XFILL_1__9011_ vdd gnd FILL
XFILL257250x115350 vdd gnd FILL
X_7989_ _7989_/D _7989_/CLK _7989_/Q vdd gnd DFFPOSX1
X_9728_ _9728_/A _9728_/B _9728_/Y vdd gnd NAND2X1
X_10610_ _10610_/A _10610_/B _10610_/C _10610_/Y vdd gnd OAI21X1
XFILL_1__9913_ vdd gnd FILL
X_11590_ _11590_/A _11590_/Y vdd gnd INVX1
X_9659_ _9659_/A _9659_/B _9659_/Y vdd gnd OR2X2
X_10541_ _10541_/A _10541_/B _10541_/Y vdd gnd NOR2X1
XFILL_1__9844_ vdd gnd FILL
X_13260_ _13260_/A _13260_/Y vdd gnd INVX1
X_10472_ _10472_/A _10472_/B _10472_/Y vdd gnd OR2X2
X_12211_ _12211_/A _12211_/B _12211_/Y vdd gnd AND2X2
X_13191_ _13191_/A _13191_/Y vdd gnd INVX1
XFILL_1__8726_ vdd gnd FILL
X_12142_ _12142_/A _12142_/Y vdd gnd INVX1
XFILL_1__8657_ vdd gnd FILL
XFILL_1__7608_ vdd gnd FILL
X_12073_ _12073_/A _12073_/B _12073_/Y vdd gnd NAND2X1
XFILL_1__8588_ vdd gnd FILL
X_11024_ _11024_/A _11024_/Y vdd gnd INVX1
XFILL_1__7539_ vdd gnd FILL
XFILL_1__10050_ vdd gnd FILL
XFILL_0__10780_ vdd gnd FILL
XFILL_1__9209_ vdd gnd FILL
XFILL_2__8002_ vdd gnd FILL
X_12975_ _12975_/A _12975_/B _12975_/Y vdd gnd NAND2X1
X_14714_ _14714_/A _14714_/B _14714_/Y vdd gnd OR2X2
X_11926_ _11926_/A _11926_/Y vdd gnd INVX1
XFILL_0__12450_ vdd gnd FILL
X_14645_ _14645_/A _14645_/B _14645_/Y vdd gnd NAND2X1
XFILL_2__10222_ vdd gnd FILL
X_11857_ _11857_/A _11857_/Y vdd gnd INVX1
XFILL_2__13010_ vdd gnd FILL
XFILL_0__11401_ vdd gnd FILL
XFILL_1__13740_ vdd gnd FILL
XFILL_0__12381_ vdd gnd FILL
XFILL_1__10952_ vdd gnd FILL
X_10808_ _10808_/A _10808_/B _10808_/C _10808_/D _10808_/Y vdd gnd AOI22X1
X_14576_ _14576_/A _14576_/Y vdd gnd INVX1
XFILL_2__10153_ vdd gnd FILL
X_11788_ _11788_/A _11788_/B _11788_/C _11788_/Y vdd gnd NAND3X1
XFILL_0__14120_ vdd gnd FILL
XFILL_0__11332_ vdd gnd FILL
XFILL_1__13671_ vdd gnd FILL
XFILL_1__10883_ vdd gnd FILL
X_13527_ _13527_/A _13527_/B _13527_/Y vdd gnd NAND2X1
X_10739_ _10739_/D _10739_/CLK _10739_/Q vdd gnd DFFPOSX1
XFILL_1__12622_ vdd gnd FILL
XFILL_2__10084_ vdd gnd FILL
XFILL_0__14051_ vdd gnd FILL
XFILL_0__11263_ vdd gnd FILL
XFILL_0__7850_ vdd gnd FILL
X_13458_ _13458_/D _13458_/CLK _13458_/Q vdd gnd DFFPOSX1
XFILL_0__13002_ vdd gnd FILL
XFILL_0__10214_ vdd gnd FILL
X_12409_ _12409_/A _12409_/B _12409_/Y vdd gnd NAND2X1
XFILL_0__11194_ vdd gnd FILL
XFILL_0__7781_ vdd gnd FILL
X_13389_ _13389_/A _13389_/B _13389_/C _13389_/Y vdd gnd OAI21X1
XFILL_1__11504_ vdd gnd FILL
XFILL_0__10145_ vdd gnd FILL
XFILL_1__12484_ vdd gnd FILL
XFILL_0__9520_ vdd gnd FILL
XFILL_2__7648_ vdd gnd FILL
XFILL_1__14223_ vdd gnd FILL
XFILL_1__11435_ vdd gnd FILL
XFILL_2__10986_ vdd gnd FILL
XFILL_0__10076_ vdd gnd FILL
XFILL_0__9451_ vdd gnd FILL
XFILL_2__7579_ vdd gnd FILL
XFILL_1__11366_ vdd gnd FILL
XFILL_0__13904_ vdd gnd FILL
XFILL_1__14154_ vdd gnd FILL
XFILL_0__8402_ vdd gnd FILL
XFILL_0__9382_ vdd gnd FILL
XFILL_1__13105_ vdd gnd FILL
XFILL_1__10317_ vdd gnd FILL
XFILL_1__14085_ vdd gnd FILL
XFILL_0__13835_ vdd gnd FILL
XFILL_1__11297_ vdd gnd FILL
XFILL_0__8333_ vdd gnd FILL
X_8961_ _8961_/A _8961_/B _8961_/Y vdd gnd NAND2X1
XFILL_1__13036_ vdd gnd FILL
XFILL_1__10248_ vdd gnd FILL
XFILL_0__10978_ vdd gnd FILL
XFILL_0__13766_ vdd gnd FILL
X_7912_ _7912_/A _7912_/B _7912_/Y vdd gnd NAND2X1
XFILL_0__8264_ vdd gnd FILL
X_8892_ _8892_/D _8892_/CLK _8892_/Q vdd gnd DFFPOSX1
XFILL_1__10179_ vdd gnd FILL
XFILL_0__12717_ vdd gnd FILL
XFILL_0__7215_ vdd gnd FILL
XFILL_0__13697_ vdd gnd FILL
X_7843_ _7843_/A _7843_/Y vdd gnd INVX1
XFILL_0__8195_ vdd gnd FILL
XFILL_0__12648_ vdd gnd FILL
XFILL_0__7146_ vdd gnd FILL
XFILL_2__13208_ vdd gnd FILL
X_7774_ _7774_/A _7774_/B _7774_/Y vdd gnd OR2X2
XFILL_1__13938_ vdd gnd FILL
X_9513_ _9513_/A _9513_/B _9513_/Y vdd gnd OR2X2
XFILL_0__7077_ vdd gnd FILL
XFILL_2__13139_ vdd gnd FILL
XFILL_0__14318_ vdd gnd FILL
XFILL_1__13869_ vdd gnd FILL
X_9444_ _9444_/A _9444_/B _9444_/C _9444_/Y vdd gnd OAI21X1
XFILL_1__7890_ vdd gnd FILL
XFILL_0__14249_ vdd gnd FILL
X_9375_ _9375_/A _9375_/B _9375_/Y vdd gnd NAND2X1
XFILL_1__9560_ vdd gnd FILL
X_8326_ _8326_/A _8326_/B _8326_/Y vdd gnd NAND2X1
XFILL_0__9718_ vdd gnd FILL
XFILL_1__8511_ vdd gnd FILL
X_8257_ _8257_/A _8257_/B _8257_/C _8257_/Y vdd gnd OAI21X1
XFILL_1__9491_ vdd gnd FILL
X_7208_ _7208_/A _7208_/B _7208_/C _7208_/Y vdd gnd AOI21X1
XFILL_0__9649_ vdd gnd FILL
XFILL_1__8442_ vdd gnd FILL
X_8188_ _8188_/A _8188_/B _8188_/Y vdd gnd NAND2X1
X_7139_ _7139_/A _7139_/B _7139_/C _7139_/Y vdd gnd OAI21X1
XFILL_1__8373_ vdd gnd FILL
XFILL_1__7324_ vdd gnd FILL
XFILL_1__7255_ vdd gnd FILL
X_12760_ _12760_/A _12760_/B _12760_/Y vdd gnd OR2X2
XFILL_1__7186_ vdd gnd FILL
X_11711_ _11711_/A _11711_/B _11711_/Y vdd gnd NAND2X1
X_12691_ _12691_/A _12691_/Y vdd gnd INVX2
X_14430_ _14430_/A _14430_/B _14430_/Y vdd gnd NAND2X1
X_11642_ _11642_/D _11642_/CLK _11642_/Q vdd gnd DFFPOSX1
X_14361_ _14361_/A _14361_/B _14361_/C _14361_/Y vdd gnd NAND3X1
X_11573_ _11573_/A _11573_/B _11573_/C _11573_/Y vdd gnd OAI21X1
X_13312_ _13312_/A _13312_/B _13312_/Y vdd gnd OR2X2
X_10524_ _10524_/A _10524_/B _10524_/Y vdd gnd OR2X2
X_14292_ _14292_/A _14292_/B _14292_/Y vdd gnd NOR2X1
XFILL_2__8620_ vdd gnd FILL
X_13243_ _13243_/A _13243_/B _13243_/C _13243_/Y vdd gnd OAI21X1
X_10455_ _10455_/A _10455_/B _10455_/C _10455_/Y vdd gnd OAI21X1
XFILL_1__9758_ vdd gnd FILL
XFILL_2_CLKBUF1_insert39 vdd gnd FILL
XFILL_2__8551_ vdd gnd FILL
X_13174_ _13174_/A _13174_/B _13174_/C _13174_/Y vdd gnd OAI21X1
XFILL_1__8709_ vdd gnd FILL
X_10386_ _10386_/A _10386_/B _10386_/C _10386_/Y vdd gnd OAI21X1
XFILL_1__9689_ vdd gnd FILL
X_12125_ _12125_/A _12125_/B _12125_/Y vdd gnd NOR2X1
XFILL_1__11220_ vdd gnd FILL
XFILL_0__11950_ vdd gnd FILL
X_12056_ _12056_/A _12056_/B _12056_/Y vdd gnd NAND2X1
XFILL_2__12510_ vdd gnd FILL
XFILL_0__10901_ vdd gnd FILL
XFILL_1__11151_ vdd gnd FILL
XFILL_0_CLKBUF1_insert32 vdd gnd FILL
X_11007_ _11007_/A _11007_/B _11007_/Y vdd gnd NAND2X1
XFILL_0__11881_ vdd gnd FILL
XFILL_0_CLKBUF1_insert43 vdd gnd FILL
XFILL_1__10102_ vdd gnd FILL
XFILL_0_CLKBUF1_insert54 vdd gnd FILL
XFILL_0_CLKBUF1_insert65 vdd gnd FILL
XFILL_2__12441_ vdd gnd FILL
XFILL_1__11082_ vdd gnd FILL
XFILL_0_CLKBUF1_insert76 vdd gnd FILL
XFILL_0__13620_ vdd gnd FILL
XFILL_0__10832_ vdd gnd FILL
XFILL_0_CLKBUF1_insert87 vdd gnd FILL
XFILL_0_CLKBUF1_insert98 vdd gnd FILL
XFILL_1__10033_ vdd gnd FILL
XFILL_1__14910_ vdd gnd FILL
XFILL_0__13551_ vdd gnd FILL
XFILL_2_BUFX2_insert361 vdd gnd FILL
XFILL_2__12372_ vdd gnd FILL
XFILL_2_BUFX2_insert372 vdd gnd FILL
XFILL_2__14111_ vdd gnd FILL
X_12958_ _12958_/A _12958_/Y vdd gnd INVX1
XFILL_0__12502_ vdd gnd FILL
XFILL_1__14841_ vdd gnd FILL
X_11909_ _11909_/A _11909_/Y vdd gnd INVX1
XFILL_2__14042_ vdd gnd FILL
X_12889_ _12889_/A _12889_/B _12889_/C _12889_/Y vdd gnd OAI21X1
XFILL_0__12433_ vdd gnd FILL
XFILL_1__14772_ vdd gnd FILL
X_14628_ _14628_/A _14628_/B _14628_/Y vdd gnd NOR2X1
XFILL_1__11984_ vdd gnd FILL
XFILL_1__13723_ vdd gnd FILL
XFILL_0__12364_ vdd gnd FILL
XFILL_1__10935_ vdd gnd FILL
X_14559_ _14559_/A _14559_/Y vdd gnd INVX1
XFILL_0__8951_ vdd gnd FILL
X_7490_ _7490_/A _7490_/B _7490_/Y vdd gnd NAND2X1
XFILL_0__14103_ vdd gnd FILL
XBUFX2_insert360 BUFX2_insert360/A BUFX2_insert360/Y vdd gnd BUFX2
XFILL_0__11315_ vdd gnd FILL
XBUFX2_insert371 BUFX2_insert371/A BUFX2_insert371/Y vdd gnd BUFX2
XFILL_1__13654_ vdd gnd FILL
XFILL_0__7902_ vdd gnd FILL
XFILL_0__12295_ vdd gnd FILL
XFILL_1__10866_ vdd gnd FILL
XBUFX2_insert382 BUFX2_insert382/A BUFX2_insert382/Y vdd gnd BUFX2
XFILL_2__10067_ vdd gnd FILL
XFILL_0__14034_ vdd gnd FILL
XFILL_0__11246_ vdd gnd FILL
XFILL_1__13585_ vdd gnd FILL
XFILL_1__10797_ vdd gnd FILL
X_9160_ _9160_/A _9160_/B _9160_/C _9160_/Y vdd gnd NAND3X1
XFILL_0__7833_ vdd gnd FILL
X_8111_ _8111_/A _8111_/B _8111_/C _8111_/Y vdd gnd NAND3X1
XFILL_0__11177_ vdd gnd FILL
X_9091_ _9091_/A _9091_/B _9091_/Y vdd gnd NOR2X1
XFILL_0__7764_ vdd gnd FILL
XFILL_0__10128_ vdd gnd FILL
XFILL_0__9503_ vdd gnd FILL
XFILL_1__12467_ vdd gnd FILL
X_8042_ _8042_/A _8042_/B _8042_/Y vdd gnd NAND2X1
XFILL_0__7695_ vdd gnd FILL
XFILL_1__11418_ vdd gnd FILL
XFILL_0__10059_ vdd gnd FILL
XFILL_1__12398_ vdd gnd FILL
XFILL_0__9434_ vdd gnd FILL
XFILL_1__14137_ vdd gnd FILL
XFILL_1__11349_ vdd gnd FILL
XFILL_0__14867_ vdd gnd FILL
XFILL_0__9365_ vdd gnd FILL
X_9993_ _9993_/A _9993_/B _9993_/C _9993_/Y vdd gnd NAND3X1
XFILL_1__14068_ vdd gnd FILL
XFILL_0__13818_ vdd gnd FILL
XFILL_0__8316_ vdd gnd FILL
XFILL_0__14798_ vdd gnd FILL
XFILL_0__9296_ vdd gnd FILL
X_8944_ _8944_/A _8944_/Y vdd gnd INVX1
XFILL_1__13019_ vdd gnd FILL
XFILL_0__13749_ vdd gnd FILL
XFILL_0__8247_ vdd gnd FILL
XFILL_2__14309_ vdd gnd FILL
X_8875_ _8875_/D _8875_/CLK _8875_/Q vdd gnd DFFPOSX1
X_7826_ _7826_/A _7826_/B _7826_/Y vdd gnd AND2X2
XFILL_0__8178_ vdd gnd FILL
XFILL_0__7129_ vdd gnd FILL
XFILL_1__8991_ vdd gnd FILL
X_7757_ _7757_/A _7757_/Y vdd gnd INVX1
X_7688_ _7688_/A _7688_/B _7688_/Y vdd gnd NOR2X1
X_9427_ _9427_/A _9427_/Y vdd gnd INVX1
XFILL_1__7873_ vdd gnd FILL
XFILL_1__9612_ vdd gnd FILL
X_9358_ _9358_/A _9358_/B _9358_/Y vdd gnd NAND2X1
X_10240_ _10240_/A _10240_/B _10240_/Y vdd gnd NAND2X1
XFILL_1__9543_ vdd gnd FILL
X_8309_ _8309_/A _8309_/B _8309_/C _8309_/Y vdd gnd NAND3X1
X_9289_ _9289_/A _9289_/B _9289_/C _9289_/D _9289_/Y vdd gnd AOI22X1
X_10171_ _10171_/A _10171_/B _10171_/Y vdd gnd NAND2X1
XFILL_1__9474_ vdd gnd FILL
XFILL_1__8425_ vdd gnd FILL
X_13930_ _13930_/A _13930_/B _13930_/Y vdd gnd NAND2X1
XFILL_1__8356_ vdd gnd FILL
X_13861_ _13861_/A _13861_/B _13861_/S _13861_/Y vdd gnd MUX2X1
XFILL_1__7307_ vdd gnd FILL
XFILL_1__8287_ vdd gnd FILL
X_12812_ _12812_/A _12812_/B _12812_/Y vdd gnd NAND2X1
XFILL_1__7238_ vdd gnd FILL
X_13792_ _13792_/A _13792_/Y vdd gnd INVX1
XFILL_1_BUFX2_insert302 vdd gnd FILL
XFILL_1_BUFX2_insert313 vdd gnd FILL
XFILL_1_BUFX2_insert324 vdd gnd FILL
XFILL_1_BUFX2_insert335 vdd gnd FILL
X_12743_ _12743_/A _12743_/B _12743_/C _12743_/Y vdd gnd OAI21X1
XFILL_1_BUFX2_insert346 vdd gnd FILL
XFILL_1__7169_ vdd gnd FILL
XFILL_1_BUFX2_insert357 vdd gnd FILL
XFILL_1_BUFX2_insert368 vdd gnd FILL
XFILL_1_BUFX2_insert379 vdd gnd FILL
X_12674_ _12674_/A _12674_/Y vdd gnd INVX1
X_14413_ _14413_/A _14413_/B _14413_/C _14413_/Y vdd gnd NAND3X1
X_11625_ _11625_/D _11625_/CLK _11625_/Q vdd gnd DFFPOSX1
X_14344_ _14344_/A _14344_/B _14344_/C _14344_/Y vdd gnd NAND3X1
X_11556_ _11556_/A _11556_/B _11556_/Y vdd gnd NAND2X1
XFILL_0__11100_ vdd gnd FILL
XFILL_1__10651_ vdd gnd FILL
XFILL_0__12080_ vdd gnd FILL
X_10507_ _10507_/A _10507_/B _10507_/Y vdd gnd NOR2X1
XFILL_2__8603_ vdd gnd FILL
X_14275_ _14275_/A _14275_/B _14275_/Y vdd gnd NAND2X1
X_11487_ _11487_/A _11487_/B _11487_/Y vdd gnd OR2X2
XFILL_0__11031_ vdd gnd FILL
XFILL_2__11941_ vdd gnd FILL
XFILL_1__10582_ vdd gnd FILL
XFILL_1__13370_ vdd gnd FILL
X_13226_ _13226_/A _13226_/Y vdd gnd INVX1
X_10438_ _10438_/A _10438_/B _10438_/C _10438_/Y vdd gnd NAND3X1
XFILL_2__8534_ vdd gnd FILL
XFILL_2__14660_ vdd gnd FILL
XFILL_1__12321_ vdd gnd FILL
XFILL_2__11872_ vdd gnd FILL
XFILL256650x21750 vdd gnd FILL
X_13157_ _13157_/A _13157_/B _13157_/Y vdd gnd NOR2X1
XFILL_2__13611_ vdd gnd FILL
X_10369_ _10369_/A _10369_/B _10369_/Y vdd gnd NAND2X1
XFILL_2__8465_ vdd gnd FILL
XFILL_1__12252_ vdd gnd FILL
XFILL_2__14591_ vdd gnd FILL
X_12108_ _12108_/A _12108_/B _12108_/Y vdd gnd NAND2X1
XFILL_0__12982_ vdd gnd FILL
X_13088_ _13088_/A _13088_/Y vdd gnd INVX1
XFILL_0__7480_ vdd gnd FILL
XFILL_1__11203_ vdd gnd FILL
XFILL_0__14721_ vdd gnd FILL
XFILL_2__8396_ vdd gnd FILL
XFILL_1__12183_ vdd gnd FILL
XFILL_0__11933_ vdd gnd FILL
X_12039_ _12039_/A _12039_/Y vdd gnd INVX1
XFILL_1__11134_ vdd gnd FILL
XFILL_0__14652_ vdd gnd FILL
XFILL_2__10685_ vdd gnd FILL
XFILL_0__11864_ vdd gnd FILL
XFILL_0__9150_ vdd gnd FILL
XFILL_0__13603_ vdd gnd FILL
XFILL_1__11065_ vdd gnd FILL
XFILL_0__8101_ vdd gnd FILL
XFILL_0__10815_ vdd gnd FILL
XFILL_0__14583_ vdd gnd FILL
XFILL_0__11795_ vdd gnd FILL
XFILL_0__9081_ vdd gnd FILL
XFILL_2__9017_ vdd gnd FILL
XFILL_1__10016_ vdd gnd FILL
XFILL_2_BUFX2_insert191 vdd gnd FILL
XFILL_0__13534_ vdd gnd FILL
XFILL_0__8032_ vdd gnd FILL
X_8660_ _8660_/A _8660_/B _8660_/Y vdd gnd NAND2X1
XFILL_2__11306_ vdd gnd FILL
XFILL_1__14824_ vdd gnd FILL
XFILL_2__12286_ vdd gnd FILL
XFILL_0__10677_ vdd gnd FILL
X_7611_ _7611_/A _7611_/B _7611_/Y vdd gnd NAND2X1
XFILL_2__14025_ vdd gnd FILL
X_8591_ _8591_/A _8591_/B _8591_/Y vdd gnd AND2X2
XFILL_2__11237_ vdd gnd FILL
XFILL_1__14755_ vdd gnd FILL
XFILL_0__12416_ vdd gnd FILL
XFILL_1__11967_ vdd gnd FILL
XFILL_0__13396_ vdd gnd FILL
X_7542_ _7542_/A _7542_/B _7542_/C _7542_/Y vdd gnd NAND3X1
XFILL_0__9983_ vdd gnd FILL
XFILL_2__9919_ vdd gnd FILL
XFILL_1__13706_ vdd gnd FILL
XFILL_0__12347_ vdd gnd FILL
XFILL_1__10918_ vdd gnd FILL
XFILL_1__14686_ vdd gnd FILL
XFILL_0__8934_ vdd gnd FILL
XFILL_1__11898_ vdd gnd FILL
X_7473_ _7473_/A _7473_/B _7473_/C _7473_/Y vdd gnd NAND3X1
XBUFX2_insert190 BUFX2_insert190/A BUFX2_insert190/Y vdd gnd BUFX2
XFILL_1__13637_ vdd gnd FILL
XFILL_0__12278_ vdd gnd FILL
XFILL_1__10849_ vdd gnd FILL
X_9212_ _9212_/A _9212_/B _9212_/C _9212_/Y vdd gnd OAI21X1
XFILL_0__11229_ vdd gnd FILL
XFILL_0__14017_ vdd gnd FILL
XFILL_1__13568_ vdd gnd FILL
XFILL_0__7816_ vdd gnd FILL
X_9143_ _9143_/A _9143_/B _9143_/Y vdd gnd AND2X2
XFILL_0__8796_ vdd gnd FILL
XFILL_2__14858_ vdd gnd FILL
XFILL_1__12519_ vdd gnd FILL
X_9074_ _9074_/A _9074_/B _9074_/C _9074_/Y vdd gnd OAI21X1
XFILL_0__7747_ vdd gnd FILL
XFILL_2__14789_ vdd gnd FILL
X_8025_ _8025_/A _8025_/B _8025_/C _8025_/Y vdd gnd OAI21X1
XFILL_0__7678_ vdd gnd FILL
XFILL_0__14919_ vdd gnd FILL
XFILL_0__9417_ vdd gnd FILL
XFILL_1__8210_ vdd gnd FILL
XFILL_1__9190_ vdd gnd FILL
XFILL_0__9348_ vdd gnd FILL
XFILL_1__8141_ vdd gnd FILL
X_9976_ _9976_/A _9976_/Y vdd gnd INVX1
XFILL_0__9279_ vdd gnd FILL
X_8927_ _8927_/A _8927_/B _8927_/C _8927_/Y vdd gnd OAI21X1
XFILL_1__8072_ vdd gnd FILL
X_8858_ _8858_/D _8858_/CLK _8858_/Q vdd gnd DFFPOSX1
X_7809_ _7809_/A _7809_/B _7809_/C _7809_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert309 vdd gnd FILL
X_8789_ _8789_/A _8789_/B _8789_/C _8789_/Y vdd gnd OAI21X1
XFILL_1__8974_ vdd gnd FILL
X_11410_ _11410_/A _11410_/B _11410_/Y vdd gnd OR2X2
X_12390_ _12390_/A _12390_/B _12390_/Y vdd gnd NAND2X1
X_11341_ _11341_/A _11341_/B _11341_/Y vdd gnd NAND2X1
XFILL_1__7856_ vdd gnd FILL
X_14060_ _14060_/A _14060_/B _14060_/Y vdd gnd OR2X2
X_11272_ _11272_/A _11272_/B _11272_/C _11272_/Y vdd gnd OAI21X1
XFILL_1__7787_ vdd gnd FILL
X_13011_ _13011_/A _13011_/B _13011_/S _13011_/Y vdd gnd MUX2X1
X_10223_ _10223_/A _10223_/B _10223_/Y vdd gnd NAND2X1
XFILL_1__9526_ vdd gnd FILL
X_10154_ _10154_/A _10154_/B _10154_/C _10154_/Y vdd gnd NAND3X1
XFILL_1__9457_ vdd gnd FILL
XFILL_2__8250_ vdd gnd FILL
XFILL_1__8408_ vdd gnd FILL
X_10085_ _10085_/A _10085_/B _10085_/Y vdd gnd NAND2X1
XFILL_1__9388_ vdd gnd FILL
XFILL_2__8181_ vdd gnd FILL
X_13913_ _13913_/A _13913_/B _13913_/C _13913_/Y vdd gnd OAI21X1
X_14893_ _14893_/D _14893_/CLK _14893_/Q vdd gnd DFFPOSX1
XFILL_1__8339_ vdd gnd FILL
XFILL_2__10470_ vdd gnd FILL
X_13844_ _13844_/A _13844_/B _13844_/C _13844_/Y vdd gnd AOI21X1
XFILL_0__10600_ vdd gnd FILL
XFILL_1_BUFX2_insert110 vdd gnd FILL
XFILL_0__11580_ vdd gnd FILL
XFILL_1_BUFX2_insert121 vdd gnd FILL
X_13775_ _13775_/A _13775_/B _13775_/C _13775_/Y vdd gnd OAI21X1
X_10987_ _10987_/A _10987_/B _10987_/C _10987_/Y vdd gnd NAND3X1
XFILL_1_BUFX2_insert132 vdd gnd FILL
XFILL_0__10531_ vdd gnd FILL
XFILL_1_BUFX2_insert143 vdd gnd FILL
XFILL_1_BUFX2_insert154 vdd gnd FILL
XFILL_1__12870_ vdd gnd FILL
XFILL_1_BUFX2_insert165 vdd gnd FILL
X_12726_ _12726_/A _12726_/B _12726_/S _12726_/Y vdd gnd MUX2X1
XFILL_1_BUFX2_insert176 vdd gnd FILL
XFILL_1_BUFX2_insert187 vdd gnd FILL
XFILL_1__11821_ vdd gnd FILL
XFILL_0__13250_ vdd gnd FILL
XFILL_1_BUFX2_insert198 vdd gnd FILL
XFILL_0__10462_ vdd gnd FILL
X_12657_ _12657_/A _12657_/B _12657_/C _12657_/Y vdd gnd OAI21X1
XFILL_2__11022_ vdd gnd FILL
XFILL_0__12201_ vdd gnd FILL
XFILL_0__13181_ vdd gnd FILL
XFILL_1__11752_ vdd gnd FILL
XFILL_0__10393_ vdd gnd FILL
X_11608_ _11608_/A _11608_/B _11608_/Y vdd gnd NAND2X1
X_12588_ _12588_/D _12588_/CLK _12588_/Q vdd gnd DFFPOSX1
XFILL_0__12132_ vdd gnd FILL
XFILL_2__7896_ vdd gnd FILL
XFILL_1__14471_ vdd gnd FILL
X_14327_ _14327_/A _14327_/B _14327_/C _14327_/Y vdd gnd NAND3X1
X_11539_ _11539_/A _11539_/Y vdd gnd INVX1
XFILL_1__13422_ vdd gnd FILL
XFILL_1__10634_ vdd gnd FILL
XFILL_0__12063_ vdd gnd FILL
XFILL_0__8650_ vdd gnd FILL
X_14258_ _14258_/A _14258_/Y vdd gnd INVX1
XFILL_0__11014_ vdd gnd FILL
XFILL_2__11924_ vdd gnd FILL
XFILL_1__13353_ vdd gnd FILL
X_13209_ _13209_/A _13209_/B _13209_/Y vdd gnd NOR2X1
XFILL_0__7601_ vdd gnd FILL
XFILL_1__10565_ vdd gnd FILL
XFILL_0__8581_ vdd gnd FILL
XFILL_2__8517_ vdd gnd FILL
X_14189_ _14189_/D _14189_/CLK _14189_/Q vdd gnd DFFPOSX1
XFILL_2__14643_ vdd gnd FILL
XFILL_1__12304_ vdd gnd FILL
XFILL_2__11855_ vdd gnd FILL
XFILL_1__10496_ vdd gnd FILL
XFILL_1__13284_ vdd gnd FILL
XFILL_0__7532_ vdd gnd FILL
XFILL_2__8448_ vdd gnd FILL
XFILL_2__14574_ vdd gnd FILL
XFILL_1__12235_ vdd gnd FILL
XFILL_2__11786_ vdd gnd FILL
XFILL_0__12965_ vdd gnd FILL
XFILL_0__7463_ vdd gnd FILL
XFILL_2__13525_ vdd gnd FILL
XFILL_0__14704_ vdd gnd FILL
XFILL_2__8379_ vdd gnd FILL
XFILL_0__9202_ vdd gnd FILL
XFILL_0__11916_ vdd gnd FILL
XFILL_1__12166_ vdd gnd FILL
X_9830_ _9830_/D _9830_/CLK _9830_/Q vdd gnd DFFPOSX1
XFILL_0__12896_ vdd gnd FILL
XFILL_0__7394_ vdd gnd FILL
XFILL_1__11117_ vdd gnd FILL
XFILL_0__14635_ vdd gnd FILL
XFILL_2__10668_ vdd gnd FILL
XFILL_1__12097_ vdd gnd FILL
XFILL_0__9133_ vdd gnd FILL
XFILL_0__11847_ vdd gnd FILL
X_9761_ _9761_/A _9761_/B _9761_/C _9761_/Y vdd gnd OAI21X1
XFILL_1__11048_ vdd gnd FILL
XFILL_0__14566_ vdd gnd FILL
XFILL_2__10599_ vdd gnd FILL
XFILL_0__9064_ vdd gnd FILL
XFILL_0__11778_ vdd gnd FILL
X_8712_ _8712_/A _8712_/Y vdd gnd INVX1
X_9692_ _9692_/A _9692_/B _9692_/C _9692_/Y vdd gnd OAI21X1
XFILL_0__13517_ vdd gnd FILL
XFILL_0__8015_ vdd gnd FILL
XFILL_0__14497_ vdd gnd FILL
X_8643_ _8643_/A _8643_/B _8643_/Y vdd gnd NAND2X1
XFILL_1__14807_ vdd gnd FILL
XFILL_1__12999_ vdd gnd FILL
X_8574_ _8574_/A _8574_/B _8574_/Y vdd gnd NAND2X1
XFILL_1__14738_ vdd gnd FILL
XFILL_0__13379_ vdd gnd FILL
X_7525_ _7525_/A _7525_/B _7525_/Y vdd gnd OR2X2
XFILL_0__9966_ vdd gnd FILL
XFILL_1__14669_ vdd gnd FILL
XFILL_1__7710_ vdd gnd FILL
XFILL_0__9897_ vdd gnd FILL
X_7456_ _7456_/A _7456_/B _7456_/C _7456_/Y vdd gnd OAI21X1
XFILL_1__8690_ vdd gnd FILL
XFILL_1__7641_ vdd gnd FILL
X_7387_ _7387_/A _7387_/B _7387_/C _7387_/Y vdd gnd OAI21X1
X_9126_ _9126_/A _9126_/B _9126_/C _9126_/D _9126_/Y vdd gnd AOI22X1
XFILL_1__7572_ vdd gnd FILL
XFILL_0__8779_ vdd gnd FILL
XFILL_1__9311_ vdd gnd FILL
X_9057_ _9057_/A _9057_/B _9057_/S _9057_/Y vdd gnd MUX2X1
XFILL_1__9242_ vdd gnd FILL
X_8008_ _8008_/A _8008_/B _8008_/Y vdd gnd NOR2X1
XFILL_1__9173_ vdd gnd FILL
X_10910_ _10910_/A _10910_/B _10910_/C _10910_/Y vdd gnd AOI21X1
XFILL_1__8124_ vdd gnd FILL
X_11890_ _11890_/A _11890_/B _11890_/C _11890_/Y vdd gnd OAI21X1
X_9959_ _9959_/A _9959_/B _9959_/C _9959_/Y vdd gnd NAND3X1
X_10841_ _10841_/A _10841_/B _10841_/Y vdd gnd NAND2X1
XFILL_1__8055_ vdd gnd FILL
X_13560_ _13560_/A _13560_/B _13560_/C _13560_/Y vdd gnd OAI21X1
X_10772_ _10772_/A _10772_/B _10772_/Y vdd gnd NOR2X1
X_12511_ _12511_/A _12511_/B _12511_/C _12511_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert117 vdd gnd FILL
X_13491_ _13491_/D _13491_/CLK _13491_/Q vdd gnd DFFPOSX1
XFILL_0_BUFX2_insert128 vdd gnd FILL
XFILL_0_BUFX2_insert139 vdd gnd FILL
X_12442_ _12442_/A _12442_/Y vdd gnd INVX1
XFILL_1__8957_ vdd gnd FILL
X_12373_ _12373_/A _12373_/B _12373_/Y vdd gnd NAND2X1
XFILL_1__7908_ vdd gnd FILL
X_14112_ _14112_/A _14112_/B _14112_/C _14112_/Y vdd gnd OAI21X1
X_11324_ _11324_/A _11324_/B _11324_/C _11324_/Y vdd gnd OAI21X1
XFILL_1__7839_ vdd gnd FILL
XFILL_1_CLKBUF1_insert386 vdd gnd FILL
X_14043_ _14043_/A _14043_/B _14043_/Y vdd gnd NAND2X1
X_11255_ _11255_/A _11255_/B _11255_/C _11255_/Y vdd gnd NAND3X1
XFILL_1__10350_ vdd gnd FILL
X_10206_ _10206_/A _10206_/B _10206_/Y vdd gnd NAND2X1
X_11186_ _11186_/A _11186_/B _11186_/Y vdd gnd NAND2X1
XFILL_1__9509_ vdd gnd FILL
XFILL_1__10281_ vdd gnd FILL
X_10137_ _10137_/A _10137_/B _10137_/C _10137_/Y vdd gnd NAND3X1
XFILL_1__12020_ vdd gnd FILL
XFILL_0__12750_ vdd gnd FILL
X_10068_ _10068_/A _10068_/B _10068_/C _10068_/Y vdd gnd OAI21X1
XFILL_2__13310_ vdd gnd FILL
XFILL_2__14290_ vdd gnd FILL
XFILL_0__11701_ vdd gnd FILL
XFILL_0__12681_ vdd gnd FILL
XFILL_2__7115_ vdd gnd FILL
X_14876_ _14876_/D _14876_/CLK _14876_/Q vdd gnd DFFPOSX1
XFILL_2__13241_ vdd gnd FILL
XFILL_2__10453_ vdd gnd FILL
XFILL_0__14420_ vdd gnd FILL
XFILL_2__8095_ vdd gnd FILL
XFILL_1__13971_ vdd gnd FILL
X_13827_ _13827_/A _13827_/B _13827_/C _13827_/Y vdd gnd NAND3X1
XFILL_2__13172_ vdd gnd FILL
XFILL_1__12922_ vdd gnd FILL
XFILL_2__10384_ vdd gnd FILL
XFILL_0__14351_ vdd gnd FILL
XFILL_0__11563_ vdd gnd FILL
X_13758_ _13758_/A _13758_/B _13758_/Y vdd gnd NOR2X1
XFILL_0__10514_ vdd gnd FILL
XFILL_0__13302_ vdd gnd FILL
XFILL_1__12853_ vdd gnd FILL
X_12709_ _12709_/A _12709_/Y vdd gnd INVX1
XFILL_0__14282_ vdd gnd FILL
XFILL_0__11494_ vdd gnd FILL
XFILL256350x43350 vdd gnd FILL
X_13689_ _13689_/A _13689_/B _13689_/Y vdd gnd NAND2X1
XFILL_1__11804_ vdd gnd FILL
XFILL_0__10445_ vdd gnd FILL
XFILL_0__13233_ vdd gnd FILL
XFILL_1__12784_ vdd gnd FILL
XFILL_2__11005_ vdd gnd FILL
XFILL_0__13164_ vdd gnd FILL
XFILL_1__11735_ vdd gnd FILL
XFILL_0__10376_ vdd gnd FILL
X_7310_ _7310_/A _7310_/B _7310_/C _7310_/Y vdd gnd NAND3X1
XFILL_0__9751_ vdd gnd FILL
XFILL256950x219750 vdd gnd FILL
X_8290_ _8290_/A _8290_/B _8290_/Y vdd gnd AND2X2
XFILL_0__12115_ vdd gnd FILL
XFILL_1__14454_ vdd gnd FILL
XFILL_0__13095_ vdd gnd FILL
XFILL_0__8702_ vdd gnd FILL
X_7241_ _7241_/A _7241_/B _7241_/C _7241_/Y vdd gnd OAI21X1
XFILL_0__9682_ vdd gnd FILL
XFILL_1__13405_ vdd gnd FILL
XFILL_1__10617_ vdd gnd FILL
XFILL_0__12046_ vdd gnd FILL
XFILL_1__14385_ vdd gnd FILL
XFILL_0__8633_ vdd gnd FILL
XFILL_1__11597_ vdd gnd FILL
X_7172_ _7172_/A _7172_/Y vdd gnd INVX1
XFILL_1__13336_ vdd gnd FILL
XFILL_1__10548_ vdd gnd FILL
XFILL_0__8564_ vdd gnd FILL
XFILL_2__11838_ vdd gnd FILL
XFILL_1__13267_ vdd gnd FILL
XFILL_0__7515_ vdd gnd FILL
XFILL_1__10479_ vdd gnd FILL
XCLKBUF1_insert385 CLKBUF1_insert385/A CLKBUF1_insert385/Y vdd gnd CLKBUF1
XFILL_0__13997_ vdd gnd FILL
XFILL_0__8495_ vdd gnd FILL
XFILL_1__12218_ vdd gnd FILL
XFILL_2__11769_ vdd gnd FILL
XFILL_0__12948_ vdd gnd FILL
XFILL_1__13198_ vdd gnd FILL
XFILL_0__7446_ vdd gnd FILL
XFILL_2__13508_ vdd gnd FILL
XFILL_1__12149_ vdd gnd FILL
X_9813_ _9813_/D _9813_/CLK _9813_/Q vdd gnd DFFPOSX1
XFILL_0__12879_ vdd gnd FILL
XFILL_0__7377_ vdd gnd FILL
XFILL_0__14618_ vdd gnd FILL
XFILL_0__9116_ vdd gnd FILL
X_9744_ _9744_/A _9744_/B _9744_/C _9744_/Y vdd gnd OAI21X1
XFILL_0__9047_ vdd gnd FILL
X_9675_ _9675_/A _9675_/B _9675_/C _9675_/Y vdd gnd OAI21X1
XFILL_1__9860_ vdd gnd FILL
X_8626_ _8626_/A _8626_/B _8626_/C _8626_/Y vdd gnd OAI21X1
XFILL_1__8811_ vdd gnd FILL
X_8557_ _8557_/A _8557_/B _8557_/C _8557_/Y vdd gnd AOI21X1
X_7508_ _7508_/A _7508_/B _7508_/C _7508_/Y vdd gnd OAI21X1
XFILL_1__8742_ vdd gnd FILL
XFILL_0__9949_ vdd gnd FILL
X_8488_ _8488_/A _8488_/B _8488_/C _8488_/Y vdd gnd AOI21X1
X_7439_ _7439_/A _7439_/B _7439_/Y vdd gnd NOR2X1
XFILL_1__8673_ vdd gnd FILL
XFILL_1__7624_ vdd gnd FILL
X_11040_ _11040_/A _11040_/B _11040_/Y vdd gnd NOR2X1
X_9109_ _9109_/A _9109_/B _9109_/C _9109_/Y vdd gnd OAI21X1
XFILL_1__7555_ vdd gnd FILL
XFILL_1__7486_ vdd gnd FILL
XFILL_1__9225_ vdd gnd FILL
X_12991_ _12991_/A _12991_/B _12991_/C _12991_/Y vdd gnd OAI21X1
XFILL257250x28950 vdd gnd FILL
X_14730_ _14730_/A _14730_/B _14730_/Y vdd gnd OR2X2
X_11942_ _11942_/A _11942_/B _11942_/C _11942_/Y vdd gnd AOI21X1
XFILL_1__9156_ vdd gnd FILL
X_14661_ _14661_/A _14661_/B _14661_/C _14661_/Y vdd gnd AOI21X1
XFILL_1__8107_ vdd gnd FILL
X_11873_ _11873_/A _11873_/B _11873_/Y vdd gnd NAND2X1
XFILL_1__9087_ vdd gnd FILL
X_13612_ _13612_/A _13612_/B _13612_/C _13612_/Y vdd gnd NAND3X1
X_10824_ _10824_/A _10824_/B _10824_/C _10824_/D _10824_/Y vdd gnd AOI22X1
X_14592_ _14592_/A _14592_/B _14592_/C _14592_/Y vdd gnd OAI21X1
XFILL_1__8038_ vdd gnd FILL
X_13543_ _13543_/A _13543_/B _13543_/C _13543_/Y vdd gnd OAI21X1
X_10755_ _10755_/D _10755_/CLK _10755_/Q vdd gnd DFFPOSX1
X_13474_ _13474_/D _13474_/CLK _13474_/Q vdd gnd DFFPOSX1
X_10686_ _10686_/A _10686_/B _10686_/Y vdd gnd NAND2X1
XFILL_0__10230_ vdd gnd FILL
XFILL_2__8782_ vdd gnd FILL
XFILL_1__9989_ vdd gnd FILL
X_12425_ _12425_/A _12425_/B _12425_/C _12425_/Y vdd gnd OAI21X1
XFILL_1__11520_ vdd gnd FILL
XFILL_0__10161_ vdd gnd FILL
X_12356_ _12356_/A _12356_/B _12356_/Y vdd gnd NAND2X1
XFILL_2__12810_ vdd gnd FILL
XFILL_1__11451_ vdd gnd FILL
XFILL_0__10092_ vdd gnd FILL
X_11307_ _11307_/A _11307_/B _11307_/Y vdd gnd NAND2X1
XFILL_2__9403_ vdd gnd FILL
X_12287_ _12287_/A _12287_/B _12287_/Y vdd gnd AND2X2
XFILL_1__10402_ vdd gnd FILL
XFILL_2__12741_ vdd gnd FILL
XFILL_0__13920_ vdd gnd FILL
XFILL_1__11382_ vdd gnd FILL
X_14026_ _14026_/A _14026_/B _14026_/C _14026_/Y vdd gnd NAND3X1
X_11238_ _11238_/A _11238_/B _11238_/C _11238_/Y vdd gnd NAND3X1
XFILL_2__9334_ vdd gnd FILL
XFILL_1__13121_ vdd gnd FILL
XFILL_1__10333_ vdd gnd FILL
XFILL_0__13851_ vdd gnd FILL
XFILL_2__14411_ vdd gnd FILL
X_11169_ _11169_/A _11169_/B _11169_/C _11169_/Y vdd gnd NAND3X1
XFILL_1__10264_ vdd gnd FILL
XFILL_0__12802_ vdd gnd FILL
XFILL_1__13052_ vdd gnd FILL
XFILL_0__7300_ vdd gnd FILL
XFILL_0__13782_ vdd gnd FILL
XFILL_0__10994_ vdd gnd FILL
XFILL_0__8280_ vdd gnd FILL
XFILL_1__12003_ vdd gnd FILL
XFILL_2__14342_ vdd gnd FILL
XFILL_1__10195_ vdd gnd FILL
XFILL_0__12733_ vdd gnd FILL
XFILL_0__7231_ vdd gnd FILL
XFILL_2__14273_ vdd gnd FILL
XFILL_0__12664_ vdd gnd FILL
XFILL_0__7162_ vdd gnd FILL
X_14859_ _14859_/A _14859_/B _14859_/C _14859_/Y vdd gnd AOI21X1
XFILL_2__13224_ vdd gnd FILL
X_7790_ _7790_/A _7790_/B _7790_/Y vdd gnd NAND2X1
XFILL_0__14403_ vdd gnd FILL
XFILL_1__13954_ vdd gnd FILL
XFILL_0__7093_ vdd gnd FILL
XFILL_2__13155_ vdd gnd FILL
XFILL_1__12905_ vdd gnd FILL
XFILL_0__14334_ vdd gnd FILL
XFILL_1__13885_ vdd gnd FILL
XFILL_0__11546_ vdd gnd FILL
X_9460_ _9460_/A _9460_/B _9460_/C _9460_/Y vdd gnd NAND3X1
XFILL_2__13086_ vdd gnd FILL
XFILL_1__12836_ vdd gnd FILL
XFILL_0__14265_ vdd gnd FILL
XFILL_0__11477_ vdd gnd FILL
X_8411_ _8411_/A _8411_/B _8411_/Y vdd gnd NAND2X1
X_9391_ _9391_/A _9391_/B _9391_/Y vdd gnd OR2X2
XFILL_0__13216_ vdd gnd FILL
XFILL_0__10428_ vdd gnd FILL
XFILL_1__12767_ vdd gnd FILL
X_8342_ _8342_/A _8342_/B _8342_/Y vdd gnd NAND2X1
XFILL_1__11718_ vdd gnd FILL
XFILL_0__13147_ vdd gnd FILL
XFILL_0__10359_ vdd gnd FILL
XFILL_1__12698_ vdd gnd FILL
XFILL_0__9734_ vdd gnd FILL
X_8273_ _8273_/A _8273_/B _8273_/C _8273_/Y vdd gnd OAI21X1
XFILL_1__14437_ vdd gnd FILL
XFILL_0__13078_ vdd gnd FILL
X_7224_ _7224_/A _7224_/B _7224_/Y vdd gnd NOR2X1
XFILL_0__9665_ vdd gnd FILL
XFILL_0__12029_ vdd gnd FILL
XFILL_1__14368_ vdd gnd FILL
XFILL_0__8616_ vdd gnd FILL
X_7155_ _7155_/A _7155_/B _7155_/C _7155_/Y vdd gnd OAI21X1
XFILL_0__9596_ vdd gnd FILL
XFILL_1__13319_ vdd gnd FILL
XFILL_1__14299_ vdd gnd FILL
XFILL_1__7340_ vdd gnd FILL
XFILL_0__8547_ vdd gnd FILL
X_7086_ _7086_/A _7086_/B _7086_/C _7086_/Y vdd gnd OAI21X1
XFILL_1__7271_ vdd gnd FILL
XFILL_0__8478_ vdd gnd FILL
XFILL_1__9010_ vdd gnd FILL
XFILL256950x104550 vdd gnd FILL
XFILL_0__7429_ vdd gnd FILL
X_7988_ _7988_/D _7988_/CLK _7988_/Q vdd gnd DFFPOSX1
X_9727_ _9727_/A _9727_/B _9727_/C _9727_/Y vdd gnd OAI21X1
XFILL_1__9912_ vdd gnd FILL
X_9658_ _9658_/A _9658_/B _9658_/C _9658_/Y vdd gnd AOI21X1
X_10540_ _10540_/A _10540_/B _10540_/C _10540_/Y vdd gnd OAI21X1
X_8609_ _8609_/A _8609_/B _8609_/C _8609_/Y vdd gnd OAI21X1
X_9589_ _9589_/A _9589_/B _9589_/Y vdd gnd OR2X2
X_10471_ _10471_/A _10471_/B _10471_/Y vdd gnd AND2X2
X_12210_ _12210_/A _12210_/B _12210_/Y vdd gnd AND2X2
X_13190_ _13190_/A _13190_/B _13190_/C _13190_/Y vdd gnd OAI21X1
XFILL_1__8725_ vdd gnd FILL
X_12141_ _12141_/A _12141_/B _12141_/C _12141_/Y vdd gnd AOI21X1
XFILL_1__8656_ vdd gnd FILL
XFILL_1__7607_ vdd gnd FILL
X_12072_ _12072_/A _12072_/B _12072_/Y vdd gnd NAND2X1
XFILL_1__8587_ vdd gnd FILL
X_11023_ _11023_/A _11023_/B _11023_/C _11023_/Y vdd gnd AOI21X1
XFILL_1__7538_ vdd gnd FILL
XFILL_2__9050_ vdd gnd FILL
XFILL_1__7469_ vdd gnd FILL
XFILL_1__9208_ vdd gnd FILL
X_12974_ _12974_/A _12974_/B _12974_/C _12974_/Y vdd gnd OAI21X1
X_14713_ _14713_/A _14713_/Y vdd gnd INVX1
XFILL_1__9139_ vdd gnd FILL
X_11925_ _11925_/A _11925_/B _11925_/C _11925_/Y vdd gnd NAND3X1
XFILL_2__11270_ vdd gnd FILL
X_14644_ _14644_/A _14644_/B _14644_/Y vdd gnd NAND2X1
X_11856_ _11856_/A _11856_/B _11856_/C _11856_/Y vdd gnd NAND3X1
XFILL_2__9952_ vdd gnd FILL
XFILL_0__11400_ vdd gnd FILL
XFILL_0__12380_ vdd gnd FILL
XFILL_1__10951_ vdd gnd FILL
X_10807_ _10807_/A _10807_/B _10807_/C _10807_/Y vdd gnd OAI21X1
X_14575_ _14575_/A _14575_/B _14575_/C _14575_/Y vdd gnd OAI21X1
X_11787_ _11787_/A _11787_/B _11787_/C _11787_/Y vdd gnd NAND3X1
XFILL_0__11331_ vdd gnd FILL
XFILL_2__9883_ vdd gnd FILL
XFILL_1__13670_ vdd gnd FILL
XFILL_1__10882_ vdd gnd FILL
X_10738_ _10738_/D _10738_/CLK _10738_/Q vdd gnd DFFPOSX1
X_13526_ _13526_/A _13526_/B _13526_/C _13526_/D _13526_/Y vdd gnd AOI22X1
XFILL_1__12621_ vdd gnd FILL
XFILL_2__8834_ vdd gnd FILL
XFILL_0__14050_ vdd gnd FILL
XFILL_0__11262_ vdd gnd FILL
X_13457_ _13457_/D _13457_/CLK _13457_/Q vdd gnd DFFPOSX1
X_10669_ _10669_/A _10669_/Y vdd gnd INVX1
XFILL_2__13911_ vdd gnd FILL
XFILL_0__10213_ vdd gnd FILL
XFILL_0__13001_ vdd gnd FILL
XFILL_2__8765_ vdd gnd FILL
X_12408_ _12408_/A _12408_/Y vdd gnd INVX1
XFILL_0__11193_ vdd gnd FILL
XFILL_0__7780_ vdd gnd FILL
X_13388_ _13388_/A _13388_/B _13388_/Y vdd gnd NAND2X1
XFILL_1__11503_ vdd gnd FILL
XFILL_2__13842_ vdd gnd FILL
XFILL_0__10144_ vdd gnd FILL
XFILL_2__8696_ vdd gnd FILL
XFILL_1__12483_ vdd gnd FILL
X_12339_ _12339_/A _12339_/B _12339_/Y vdd gnd NAND2X1
XFILL_1__14222_ vdd gnd FILL
XFILL_1__11434_ vdd gnd FILL
XFILL_2__13773_ vdd gnd FILL
XFILL_0__10075_ vdd gnd FILL
XFILL_0__9450_ vdd gnd FILL
XFILL_2__12724_ vdd gnd FILL
XFILL_0__13903_ vdd gnd FILL
XFILL_1__14153_ vdd gnd FILL
XFILL_0__8401_ vdd gnd FILL
XFILL_1__11365_ vdd gnd FILL
X_14009_ _14009_/A _14009_/B _14009_/Y vdd gnd NOR2X1
XFILL_0__9381_ vdd gnd FILL
XFILL_1__13104_ vdd gnd FILL
XFILL_2__9317_ vdd gnd FILL
XFILL_2__12655_ vdd gnd FILL
XFILL_1__10316_ vdd gnd FILL
XFILL_1__14084_ vdd gnd FILL
XFILL_0__13834_ vdd gnd FILL
XFILL_0__8332_ vdd gnd FILL
XFILL_1__11296_ vdd gnd FILL
X_8960_ _8960_/A _8960_/B _8960_/C _8960_/D _8960_/Y vdd gnd AOI22X1
XFILL_2__11606_ vdd gnd FILL
XFILL_2__9248_ vdd gnd FILL
XFILL_1__13035_ vdd gnd FILL
XFILL_1__10247_ vdd gnd FILL
XFILL_0__13765_ vdd gnd FILL
XFILL_0__10977_ vdd gnd FILL
X_7911_ _7911_/A _7911_/B _7911_/C _7911_/Y vdd gnd OAI21X1
XFILL_0__8263_ vdd gnd FILL
XFILL_2__14325_ vdd gnd FILL
XFILL_2__9179_ vdd gnd FILL
X_8891_ _8891_/D _8891_/CLK _8891_/Q vdd gnd DFFPOSX1
XFILL_2__11537_ vdd gnd FILL
XFILL_0__12716_ vdd gnd FILL
XFILL_0__7214_ vdd gnd FILL
XFILL_1__10178_ vdd gnd FILL
XFILL_0__13696_ vdd gnd FILL
X_7842_ _7842_/A _7842_/B _7842_/C _7842_/Y vdd gnd OAI21X1
XFILL_0__8194_ vdd gnd FILL
XFILL_2__14256_ vdd gnd FILL
XFILL_2__11468_ vdd gnd FILL
XFILL_0__12647_ vdd gnd FILL
XFILL_0__7145_ vdd gnd FILL
X_7773_ _7773_/A _7773_/B _7773_/Y vdd gnd NAND2X1
XFILL_1__13937_ vdd gnd FILL
XFILL_2__11399_ vdd gnd FILL
X_9512_ _9512_/A _9512_/B _9512_/Y vdd gnd NAND2X1
XFILL_0__7076_ vdd gnd FILL
XFILL_0__14317_ vdd gnd FILL
XFILL_1__13868_ vdd gnd FILL
XFILL_0__11529_ vdd gnd FILL
X_9443_ _9443_/A _9443_/B _9443_/Y vdd gnd NOR2X1
XFILL_1__12819_ vdd gnd FILL
XFILL_2__13069_ vdd gnd FILL
XFILL_0__14248_ vdd gnd FILL
XFILL_1__13799_ vdd gnd FILL
X_9374_ _9374_/A _9374_/B _9374_/Y vdd gnd NAND2X1
X_8325_ _8325_/A _8325_/B _8325_/C _8325_/Y vdd gnd OAI21X1
XFILL_1__8510_ vdd gnd FILL
XFILL_0__9717_ vdd gnd FILL
XFILL_1__9490_ vdd gnd FILL
X_8256_ _8256_/A _8256_/Y vdd gnd INVX1
X_7207_ _7207_/A _7207_/B _7207_/Y vdd gnd NAND2X1
XFILL_1__8441_ vdd gnd FILL
XFILL_0__9648_ vdd gnd FILL
X_8187_ _8187_/A _8187_/B _8187_/C _8187_/Y vdd gnd OAI21X1
X_7138_ _7138_/A _7138_/B _7138_/Y vdd gnd NAND2X1
XFILL_0__9579_ vdd gnd FILL
XFILL_1__8372_ vdd gnd FILL
XFILL_1__7323_ vdd gnd FILL
XFILL_1__7254_ vdd gnd FILL
XFILL_1__7185_ vdd gnd FILL
X_11710_ _11710_/A _11710_/Y vdd gnd INVX1
X_12690_ _12690_/A _12690_/B _12690_/C _12690_/Y vdd gnd OAI21X1
X_11641_ _11641_/D _11641_/CLK _11641_/Q vdd gnd DFFPOSX1
X_14360_ _14360_/A _14360_/B _14360_/C _14360_/Y vdd gnd OAI21X1
X_11572_ _11572_/A _11572_/B _11572_/Y vdd gnd NAND2X1
X_13311_ _13311_/A _13311_/B _13311_/Y vdd gnd NAND2X1
X_10523_ _10523_/A _10523_/B _10523_/C _10523_/Y vdd gnd OAI21X1
X_14291_ _14291_/A _14291_/B _14291_/C _14291_/D _14291_/Y vdd gnd AOI22X1
X_13242_ _13242_/A _13242_/B _13242_/C _13242_/Y vdd gnd OAI21X1
X_10454_ _10454_/A _10454_/B _10454_/Y vdd gnd AND2X2
XFILL_2_CLKBUF1_insert29 vdd gnd FILL
XFILL_1__9757_ vdd gnd FILL
X_13173_ _13173_/A _13173_/B _13173_/Y vdd gnd OR2X2
XFILL_2__7501_ vdd gnd FILL
X_10385_ _10385_/A _10385_/B _10385_/Y vdd gnd NAND2X1
XFILL_1__8708_ vdd gnd FILL
XFILL_2__8481_ vdd gnd FILL
XFILL_1__9688_ vdd gnd FILL
X_12124_ _12124_/A _12124_/B _12124_/Y vdd gnd AND2X2
XFILL_2__7432_ vdd gnd FILL
XFILL_1__8639_ vdd gnd FILL
X_12055_ _12055_/A _12055_/Y vdd gnd INVX1
XFILL_0__10900_ vdd gnd FILL
XFILL_1__11150_ vdd gnd FILL
X_11006_ _11006_/A _11006_/B _11006_/C _11006_/Y vdd gnd NAND3X1
XFILL257550x97350 vdd gnd FILL
XFILL_0__11880_ vdd gnd FILL
XFILL_0_CLKBUF1_insert33 vdd gnd FILL
XFILL_2__9102_ vdd gnd FILL
XFILL_0_CLKBUF1_insert44 vdd gnd FILL
XFILL_1__10101_ vdd gnd FILL
XFILL_0_CLKBUF1_insert55 vdd gnd FILL
XFILL_0_CLKBUF1_insert66 vdd gnd FILL
XFILL_1__11081_ vdd gnd FILL
XFILL_0__10831_ vdd gnd FILL
XFILL_0_CLKBUF1_insert77 vdd gnd FILL
XFILL_2__9033_ vdd gnd FILL
XFILL_0_CLKBUF1_insert88 vdd gnd FILL
XFILL_0_CLKBUF1_insert99 vdd gnd FILL
XFILL_1__10032_ vdd gnd FILL
XFILL_2_BUFX2_insert351 vdd gnd FILL
XFILL_0__13550_ vdd gnd FILL
XFILL_2__11322_ vdd gnd FILL
X_12957_ _12957_/A _12957_/B _12957_/Y vdd gnd NAND2X1
XFILL_1__14840_ vdd gnd FILL
XFILL_0__12501_ vdd gnd FILL
X_11908_ _11908_/A _11908_/B _11908_/C _11908_/Y vdd gnd NOR3X1
XFILL_2__11253_ vdd gnd FILL
X_12888_ _12888_/A _12888_/Y vdd gnd INVX1
XFILL_1__14771_ vdd gnd FILL
XFILL_0__12432_ vdd gnd FILL
XFILL_1__11983_ vdd gnd FILL
X_14627_ _14627_/A _14627_/B _14627_/Y vdd gnd AND2X2
X_11839_ _11839_/A _11839_/B _11839_/Y vdd gnd NAND2X1
XFILL_2__9935_ vdd gnd FILL
XFILL_1__13722_ vdd gnd FILL
XFILL_2__11184_ vdd gnd FILL
XFILL_1__10934_ vdd gnd FILL
XFILL_0__12363_ vdd gnd FILL
XFILL_0__8950_ vdd gnd FILL
X_14558_ _14558_/A _14558_/Y vdd gnd INVX1
XFILL_0__14102_ vdd gnd FILL
XBUFX2_insert350 BUFX2_insert350/A BUFX2_insert350/Y vdd gnd BUFX2
XFILL_2__9866_ vdd gnd FILL
XFILL_0__11314_ vdd gnd FILL
XFILL_1__13653_ vdd gnd FILL
XBUFX2_insert361 BUFX2_insert361/A BUFX2_insert361/Y vdd gnd BUFX2
XFILL_1__10865_ vdd gnd FILL
XBUFX2_insert372 BUFX2_insert372/A BUFX2_insert372/Y vdd gnd BUFX2
XFILL_0__7901_ vdd gnd FILL
XFILL_0__12294_ vdd gnd FILL
X_13509_ _13509_/A _13509_/B _13509_/Y vdd gnd NOR2X1
XBUFX2_insert383 BUFX2_insert383/A BUFX2_insert383/Y vdd gnd BUFX2
XFILL_2__8817_ vdd gnd FILL
X_14489_ _14489_/A _14489_/B _14489_/C _14489_/Y vdd gnd OAI21X1
XFILL_0__14033_ vdd gnd FILL
XFILL_1__13584_ vdd gnd FILL
XFILL_0__11245_ vdd gnd FILL
XFILL_0__7832_ vdd gnd FILL
XFILL_1__10796_ vdd gnd FILL
XFILL_2__8748_ vdd gnd FILL
XFILL_1__12535_ vdd gnd FILL
XFILL_0__11176_ vdd gnd FILL
X_8110_ _8110_/A _8110_/B _8110_/S _8110_/Y vdd gnd MUX2X1
XFILL_0__7763_ vdd gnd FILL
X_9090_ _9090_/A _9090_/B _9090_/Y vdd gnd NOR2X1
XFILL_0__10127_ vdd gnd FILL
XFILL_2__13825_ vdd gnd FILL
XFILL_1__12466_ vdd gnd FILL
XFILL_2__8679_ vdd gnd FILL
XFILL_0__9502_ vdd gnd FILL
X_8041_ _8041_/A _8041_/Y vdd gnd INVX1
XFILL_0__7694_ vdd gnd FILL
XFILL_1__11417_ vdd gnd FILL
XFILL_0__10058_ vdd gnd FILL
XFILL_2__13756_ vdd gnd FILL
XFILL_0__9433_ vdd gnd FILL
XFILL_1__12397_ vdd gnd FILL
XFILL_2__12707_ vdd gnd FILL
XFILL_1__14136_ vdd gnd FILL
XFILL_1__11348_ vdd gnd FILL
XFILL_2__13687_ vdd gnd FILL
XFILL_0__14866_ vdd gnd FILL
XFILL_0__9364_ vdd gnd FILL
X_9992_ _9992_/A _9992_/B _9992_/C _9992_/Y vdd gnd AOI21X1
XFILL_2__12638_ vdd gnd FILL
XFILL_1__14067_ vdd gnd FILL
XFILL_0__13817_ vdd gnd FILL
XFILL_0__8315_ vdd gnd FILL
XFILL_1__11279_ vdd gnd FILL
XFILL_0__14797_ vdd gnd FILL
XFILL_0__9295_ vdd gnd FILL
X_8943_ _8943_/A _8943_/B _8943_/Y vdd gnd NAND2X1
XFILL_1__13018_ vdd gnd FILL
XFILL_0__13748_ vdd gnd FILL
XFILL_0__8246_ vdd gnd FILL
X_8874_ _8874_/D _8874_/CLK _8874_/Q vdd gnd DFFPOSX1
XFILL_0__13679_ vdd gnd FILL
X_7825_ _7825_/A _7825_/B _7825_/Y vdd gnd NAND2X1
XFILL_0__8177_ vdd gnd FILL
XFILL_2__14239_ vdd gnd FILL
XFILL_0__7128_ vdd gnd FILL
X_7756_ _7756_/A _7756_/B _7756_/Y vdd gnd NAND2X1
XFILL_1__8990_ vdd gnd FILL
X_7687_ _7687_/A _7687_/Y vdd gnd INVX1
X_9426_ _9426_/A _9426_/B _9426_/C _9426_/Y vdd gnd NOR3X1
XFILL_1__7872_ vdd gnd FILL
XFILL_1__9611_ vdd gnd FILL
X_9357_ _9357_/A _9357_/Y vdd gnd INVX1
X_8308_ _8308_/A _8308_/B _8308_/C _8308_/Y vdd gnd OAI21X1
XFILL_1__9542_ vdd gnd FILL
X_9288_ _9288_/A _9288_/B _9288_/Y vdd gnd NOR2X1
X_10170_ _10170_/A _10170_/B _10170_/C _10170_/Y vdd gnd NAND3X1
XFILL_1__9473_ vdd gnd FILL
X_8239_ _8239_/A _8239_/B _8239_/Y vdd gnd NOR2X1
XFILL_1__8424_ vdd gnd FILL
XFILL_1__8355_ vdd gnd FILL
XFILL_1__7306_ vdd gnd FILL
X_13860_ _13860_/A _13860_/B _13860_/C _13860_/Y vdd gnd OAI21X1
XFILL_1__8286_ vdd gnd FILL
X_12811_ _12811_/A _12811_/B _12811_/C _12811_/Y vdd gnd OAI21X1
XFILL_1__7237_ vdd gnd FILL
X_13791_ _13791_/A _13791_/B _13791_/C _13791_/Y vdd gnd AOI21X1
XFILL_1_BUFX2_insert303 vdd gnd FILL
XFILL_1_BUFX2_insert314 vdd gnd FILL
X_12742_ _12742_/A _12742_/B _12742_/Y vdd gnd NAND2X1
XFILL_1_BUFX2_insert325 vdd gnd FILL
XFILL_1__7168_ vdd gnd FILL
XFILL_1_BUFX2_insert336 vdd gnd FILL
XFILL_1_BUFX2_insert347 vdd gnd FILL
XFILL_1_BUFX2_insert358 vdd gnd FILL
XFILL_1_BUFX2_insert369 vdd gnd FILL
X_12673_ _12673_/A _12673_/B _12673_/C _12673_/Y vdd gnd OAI21X1
XFILL_1__7099_ vdd gnd FILL
X_14412_ _14412_/A _14412_/B _14412_/Y vdd gnd NOR2X1
X_11624_ _11624_/D _11624_/CLK _11624_/Q vdd gnd DFFPOSX1
XFILL_2__9720_ vdd gnd FILL
XFILL257550x72150 vdd gnd FILL
X_14343_ _14343_/A _14343_/B _14343_/C _14343_/Y vdd gnd OAI21X1
X_11555_ _11555_/A _11555_/B _11555_/C _11555_/Y vdd gnd OAI21X1
XFILL_2__9651_ vdd gnd FILL
XFILL_1__10650_ vdd gnd FILL
X_10506_ _10506_/A _10506_/B _10506_/C _10506_/Y vdd gnd AOI21X1
X_14274_ _14274_/A _14274_/B _14274_/Y vdd gnd NAND2X1
X_11486_ _11486_/A _11486_/B _11486_/Y vdd gnd NAND2X1
XFILL_0__11030_ vdd gnd FILL
XFILL_1__10581_ vdd gnd FILL
X_13225_ _13225_/A _13225_/B _13225_/Y vdd gnd NAND2X1
X_10437_ _10437_/A _10437_/B _10437_/Y vdd gnd OR2X2
XFILL_1__12320_ vdd gnd FILL
X_13156_ _13156_/A _13156_/B _13156_/C _13156_/Y vdd gnd OAI21X1
X_10368_ _10368_/A _10368_/B _10368_/C _10368_/Y vdd gnd OAI21X1
XFILL_2__10822_ vdd gnd FILL
XFILL_1__12251_ vdd gnd FILL
X_12107_ _12107_/A _12107_/B _12107_/Y vdd gnd NAND2X1
XFILL_0__12981_ vdd gnd FILL
X_13087_ _13087_/A _13087_/B _13087_/C _13087_/D _13087_/Y vdd gnd AOI22X1
XFILL_2__7415_ vdd gnd FILL
X_10299_ _10299_/A _10299_/B _10299_/Y vdd gnd NAND2X1
XFILL_2__13541_ vdd gnd FILL
XFILL_1__11202_ vdd gnd FILL
XFILL_0__14720_ vdd gnd FILL
XFILL_0__11932_ vdd gnd FILL
XFILL_1__12182_ vdd gnd FILL
X_12038_ _12038_/A _12038_/B _12038_/Y vdd gnd NAND2X1
XFILL_2__7346_ vdd gnd FILL
XFILL_1__11133_ vdd gnd FILL
XFILL_0__14651_ vdd gnd FILL
XFILL_0__11863_ vdd gnd FILL
XFILL_2__7277_ vdd gnd FILL
XFILL_0__13602_ vdd gnd FILL
XFILL_0__8100_ vdd gnd FILL
XFILL_0__10814_ vdd gnd FILL
XFILL_1__11064_ vdd gnd FILL
XFILL_0__14582_ vdd gnd FILL
XFILL_0__9080_ vdd gnd FILL
XFILL_0__11794_ vdd gnd FILL
XFILL_2_BUFX2_insert170 vdd gnd FILL
XFILL_1__10015_ vdd gnd FILL
X_13989_ _13989_/A _13989_/B _13989_/Y vdd gnd NAND2X1
XFILL_0__13533_ vdd gnd FILL
XFILL_0__8031_ vdd gnd FILL
XFILL_1__14823_ vdd gnd FILL
X_7610_ _7610_/A _7610_/B _7610_/C _7610_/Y vdd gnd NAND3X1
XFILL_0__10676_ vdd gnd FILL
X_8590_ _8590_/A _8590_/B _8590_/C _8590_/Y vdd gnd NAND3X1
XFILL_1__14754_ vdd gnd FILL
XFILL_0__12415_ vdd gnd FILL
XFILL_1__11966_ vdd gnd FILL
XFILL_0__13395_ vdd gnd FILL
X_7541_ _7541_/A _7541_/B _7541_/C _7541_/Y vdd gnd OAI21X1
XFILL_0__9982_ vdd gnd FILL
XFILL_1__13705_ vdd gnd FILL
XFILL_2__11167_ vdd gnd FILL
XFILL_1__10917_ vdd gnd FILL
XFILL_1__14685_ vdd gnd FILL
XFILL_0__12346_ vdd gnd FILL
XFILL_1__11897_ vdd gnd FILL
XFILL_0__8933_ vdd gnd FILL
X_7472_ _7472_/A _7472_/B _7472_/C _7472_/Y vdd gnd OAI21X1
XFILL_1__13636_ vdd gnd FILL
XBUFX2_insert180 BUFX2_insert180/A BUFX2_insert180/Y vdd gnd BUFX2
XBUFX2_insert191 BUFX2_insert191/A BUFX2_insert191/Y vdd gnd BUFX2
XFILL_1__10848_ vdd gnd FILL
XFILL_2__11098_ vdd gnd FILL
X_9211_ _9211_/A _9211_/B _9211_/C _9211_/Y vdd gnd NAND3X1
XFILL_0__12277_ vdd gnd FILL
XFILL_0__14016_ vdd gnd FILL
XFILL_0__11228_ vdd gnd FILL
XFILL_1__13567_ vdd gnd FILL
XFILL_1__10779_ vdd gnd FILL
X_9142_ _9142_/A _9142_/B _9142_/Y vdd gnd NAND2X1
XFILL_0__7815_ vdd gnd FILL
XFILL_1__12518_ vdd gnd FILL
XFILL_0__8795_ vdd gnd FILL
XFILL_0__11159_ vdd gnd FILL
X_9073_ _9073_/A _9073_/Y vdd gnd INVX1
XFILL_0__7746_ vdd gnd FILL
XFILL_2__13808_ vdd gnd FILL
XFILL_1__12449_ vdd gnd FILL
X_8024_ _8024_/A _8024_/B _8024_/Y vdd gnd NAND2X1
XFILL_0__7677_ vdd gnd FILL
XFILL_2__13739_ vdd gnd FILL
XFILL_0__14918_ vdd gnd FILL
XFILL_0__9416_ vdd gnd FILL
XFILL_1__14119_ vdd gnd FILL
XFILL_0__14849_ vdd gnd FILL
XFILL_1__8140_ vdd gnd FILL
XFILL_0__9347_ vdd gnd FILL
X_9975_ _9975_/A _9975_/B _9975_/C _9975_/Y vdd gnd OAI21X1
XFILL_0__9278_ vdd gnd FILL
X_8926_ _8926_/A _8926_/B _8926_/Y vdd gnd NOR2X1
XFILL_1__8071_ vdd gnd FILL
XFILL_0__8229_ vdd gnd FILL
X_8857_ _8857_/D _8857_/CLK _8857_/Q vdd gnd DFFPOSX1
X_7808_ _7808_/A _7808_/B _7808_/Y vdd gnd NAND2X1
X_8788_ _8788_/A _8788_/B _8788_/Y vdd gnd NAND2X1
X_7739_ _7739_/A _7739_/B _7739_/C _7739_/Y vdd gnd OAI21X1
XFILL_1__8973_ vdd gnd FILL
X_11340_ _11340_/A _11340_/B _11340_/C _11340_/Y vdd gnd OAI21X1
X_9409_ _9409_/A _9409_/B _9409_/C _9409_/Y vdd gnd NAND3X1
XFILL_1__7855_ vdd gnd FILL
X_11271_ _11271_/A _11271_/B _11271_/Y vdd gnd NAND2X1
XFILL256650x183750 vdd gnd FILL
XFILL_1__7786_ vdd gnd FILL
X_13010_ _13010_/A _13010_/B _13010_/C _13010_/Y vdd gnd NAND3X1
X_10222_ _10222_/A _10222_/B _10222_/Y vdd gnd NOR2X1
XFILL_1__9525_ vdd gnd FILL
X_10153_ _10153_/A _10153_/B _10153_/C _10153_/Y vdd gnd OAI21X1
XFILL_1__9456_ vdd gnd FILL
XFILL_2__7200_ vdd gnd FILL
X_10084_ _10084_/A _10084_/B _10084_/C _10084_/Y vdd gnd NAND3X1
XFILL_1__8407_ vdd gnd FILL
XFILL_1__9387_ vdd gnd FILL
X_13912_ _13912_/A _13912_/B _13912_/C _13912_/Y vdd gnd AOI21X1
XFILL_2__7131_ vdd gnd FILL
X_14892_ _14892_/D _14892_/CLK _14892_/Q vdd gnd DFFPOSX1
XFILL_1__8338_ vdd gnd FILL
X_13843_ _13843_/A _13843_/B _13843_/C _13843_/Y vdd gnd NOR3X1
XFILL_1__8269_ vdd gnd FILL
XFILL_1_BUFX2_insert111 vdd gnd FILL
X_10986_ _10986_/A _10986_/B _10986_/C _10986_/Y vdd gnd OAI21X1
XFILL_1_BUFX2_insert122 vdd gnd FILL
X_13774_ _13774_/A _13774_/Y vdd gnd INVX1
XFILL_1_BUFX2_insert133 vdd gnd FILL
XFILL_0__10530_ vdd gnd FILL
XFILL_1_BUFX2_insert144 vdd gnd FILL
XFILL_1_BUFX2_insert155 vdd gnd FILL
X_12725_ _12725_/A _12725_/B _12725_/S _12725_/Y vdd gnd MUX2X1
XFILL_1_BUFX2_insert166 vdd gnd FILL
XFILL_1_BUFX2_insert177 vdd gnd FILL
XFILL_1__11820_ vdd gnd FILL
XFILL_2__12070_ vdd gnd FILL
XFILL_1_BUFX2_insert188 vdd gnd FILL
XFILL_0__10461_ vdd gnd FILL
XFILL_1_BUFX2_insert199 vdd gnd FILL
X_12656_ _12656_/A _12656_/B _12656_/C _12656_/Y vdd gnd OAI21X1
XFILL_0__12200_ vdd gnd FILL
XFILL_1__11751_ vdd gnd FILL
XFILL_0__13180_ vdd gnd FILL
XFILL_0__10392_ vdd gnd FILL
X_11607_ _11607_/A _11607_/B _11607_/C _11607_/Y vdd gnd OAI21X1
XFILL_2__9703_ vdd gnd FILL
X_12587_ _12587_/D _12587_/CLK _12587_/Q vdd gnd DFFPOSX1
XFILL_0__12131_ vdd gnd FILL
XFILL_1__14470_ vdd gnd FILL
X_14326_ _14326_/A _14326_/B _14326_/Y vdd gnd NOR2X1
X_11538_ _11538_/A _11538_/B _11538_/C _11538_/Y vdd gnd OAI21X1
XFILL_2__9634_ vdd gnd FILL
XFILL_1__13421_ vdd gnd FILL
XFILL_1__10633_ vdd gnd FILL
XFILL_0__12062_ vdd gnd FILL
XFILL_2__12972_ vdd gnd FILL
X_14257_ _14257_/A _14257_/Y vdd gnd INVX4
X_11469_ _11469_/A _11469_/B _11469_/Y vdd gnd NAND2X1
XFILL_0__11013_ vdd gnd FILL
XFILL_2__9565_ vdd gnd FILL
XFILL_1__13352_ vdd gnd FILL
XFILL_1__10564_ vdd gnd FILL
X_13208_ _13208_/A _13208_/B _13208_/Y vdd gnd AND2X2
XFILL_0__7600_ vdd gnd FILL
XFILL_0__8580_ vdd gnd FILL
XFILL_1__12303_ vdd gnd FILL
X_14188_ _14188_/D _14188_/CLK _14188_/Q vdd gnd DFFPOSX1
XFILL_2__9496_ vdd gnd FILL
XFILL_1__13283_ vdd gnd FILL
XFILL_0__7531_ vdd gnd FILL
XFILL_1__10495_ vdd gnd FILL
X_13139_ _13139_/A _13139_/B _13139_/Y vdd gnd NOR2X1
XFILL_1__12234_ vdd gnd FILL
XFILL_2__10805_ vdd gnd FILL
XFILL_0__12964_ vdd gnd FILL
XFILL_0__7462_ vdd gnd FILL
XFILL_0__14703_ vdd gnd FILL
XFILL_0__11915_ vdd gnd FILL
XFILL_1__12165_ vdd gnd FILL
XFILL_0__9201_ vdd gnd FILL
XFILL_0__12895_ vdd gnd FILL
XFILL_0__7393_ vdd gnd FILL
XFILL_2__7329_ vdd gnd FILL
XFILL_1__11116_ vdd gnd FILL
XFILL_0__14634_ vdd gnd FILL
XFILL_0__9132_ vdd gnd FILL
XFILL_0__11846_ vdd gnd FILL
XFILL_1__12096_ vdd gnd FILL
X_9760_ _9760_/A _9760_/B _9760_/Y vdd gnd NAND2X1
XFILL_2__12406_ vdd gnd FILL
XFILL_2__13386_ vdd gnd FILL
XFILL_1__11047_ vdd gnd FILL
XFILL_0__14565_ vdd gnd FILL
XFILL_0__9063_ vdd gnd FILL
X_8711_ _8711_/A _8711_/B _8711_/Y vdd gnd NOR2X1
XFILL_0__11777_ vdd gnd FILL
X_9691_ _9691_/A _9691_/Y vdd gnd INVX1
XFILL_0__13516_ vdd gnd FILL
XFILL_0__8014_ vdd gnd FILL
XFILL_0__14496_ vdd gnd FILL
X_8642_ _8642_/A _8642_/B _8642_/Y vdd gnd NAND2X1
XFILL_1__14806_ vdd gnd FILL
XFILL_0__10659_ vdd gnd FILL
XFILL_1__12998_ vdd gnd FILL
X_8573_ _8573_/A _8573_/B _8573_/Y vdd gnd NAND2X1
XFILL_1__14737_ vdd gnd FILL
XFILL_1__11949_ vdd gnd FILL
XFILL_0__13378_ vdd gnd FILL
X_7524_ _7524_/A _7524_/B _7524_/Y vdd gnd NAND2X1
XFILL_0__9965_ vdd gnd FILL
XFILL_0__12329_ vdd gnd FILL
XFILL_1__14668_ vdd gnd FILL
X_7455_ _7455_/A _7455_/B _7455_/C _7455_/Y vdd gnd OAI21X1
XFILL_0__9896_ vdd gnd FILL
XFILL_1__13619_ vdd gnd FILL
XFILL_1__14599_ vdd gnd FILL
XFILL_1__7640_ vdd gnd FILL
X_7386_ _7386_/A _7386_/B _7386_/C _7386_/Y vdd gnd NAND3X1
XFILL_2__14909_ vdd gnd FILL
X_9125_ _9125_/A _9125_/B _9125_/C _9125_/Y vdd gnd OAI21X1
XFILL_1__7571_ vdd gnd FILL
XFILL_0__8778_ vdd gnd FILL
XFILL_1__9310_ vdd gnd FILL
X_9056_ _9056_/A _9056_/B _9056_/C _9056_/Y vdd gnd AOI21X1
XFILL_0__7729_ vdd gnd FILL
X_8007_ _8007_/A _8007_/B _8007_/C _8007_/Y vdd gnd OAI21X1
XFILL_1__9241_ vdd gnd FILL
XFILL_1__9172_ vdd gnd FILL
XFILL_1__8123_ vdd gnd FILL
X_9958_ _9958_/A _9958_/B _9958_/S _9958_/Y vdd gnd MUX2X1
X_10840_ _10840_/A _10840_/Y vdd gnd INVX1
XFILL_1__8054_ vdd gnd FILL
X_8909_ _8909_/D _8909_/CLK _8909_/Q vdd gnd DFFPOSX1
X_9889_ _9889_/A _9889_/Y vdd gnd INVX1
X_10771_ _10771_/A _10771_/Y vdd gnd INVX2
X_12510_ _12510_/A _12510_/B _12510_/Y vdd gnd NAND2X1
X_13490_ _13490_/D _13490_/CLK _13490_/Q vdd gnd DFFPOSX1
XFILL_0_BUFX2_insert118 vdd gnd FILL
XFILL_0_BUFX2_insert129 vdd gnd FILL
X_12441_ _12441_/A _12441_/B _12441_/C _12441_/Y vdd gnd AOI21X1
XFILL_1__8956_ vdd gnd FILL
X_12372_ _12372_/A _12372_/B _12372_/Y vdd gnd OR2X2
XFILL_1__7907_ vdd gnd FILL
X_14111_ _14111_/A _14111_/B _14111_/C _14111_/Y vdd gnd OAI21X1
X_11323_ _11323_/A _11323_/B _11323_/C _11323_/Y vdd gnd NAND3X1
XFILL_1__7838_ vdd gnd FILL
XFILL_1_CLKBUF1_insert387 vdd gnd FILL
X_11254_ _11254_/A _11254_/Y vdd gnd INVX1
X_14042_ _14042_/A _14042_/B _14042_/C _14042_/Y vdd gnd OAI21X1
XFILL_2__9350_ vdd gnd FILL
XFILL_1__7769_ vdd gnd FILL
X_10205_ _10205_/A _10205_/B _10205_/Y vdd gnd NAND2X1
X_11185_ _11185_/A _11185_/B _11185_/C _11185_/Y vdd gnd OAI21X1
XFILL_1__9508_ vdd gnd FILL
XFILL_2__9281_ vdd gnd FILL
XFILL_1__10280_ vdd gnd FILL
X_10136_ _10136_/A _10136_/B _10136_/C _10136_/Y vdd gnd OAI21X1
XFILL_1__9439_ vdd gnd FILL
XFILL_2__11570_ vdd gnd FILL
X_10067_ _10067_/A _10067_/B _10067_/Y vdd gnd AND2X2
XFILL_0__11700_ vdd gnd FILL
XFILL_0__12680_ vdd gnd FILL
X_14875_ _14875_/D _14875_/CLK _14875_/Q vdd gnd DFFPOSX1
XFILL_1__13970_ vdd gnd FILL
X_13826_ _13826_/A _13826_/B _13826_/Y vdd gnd AND2X2
XFILL_1__12921_ vdd gnd FILL
XFILL_0__14350_ vdd gnd FILL
XFILL_0__11562_ vdd gnd FILL
XFILL_2__12122_ vdd gnd FILL
X_13757_ _13757_/A _13757_/Y vdd gnd INVX1
X_10969_ _10969_/A _10969_/B _10969_/Y vdd gnd AND2X2
XFILL_0__13301_ vdd gnd FILL
XFILL_0__10513_ vdd gnd FILL
XFILL_1__12852_ vdd gnd FILL
XFILL_0__14281_ vdd gnd FILL
XFILL_0__11493_ vdd gnd FILL
X_12708_ _12708_/A _12708_/Y vdd gnd INVX8
XFILL_2__12053_ vdd gnd FILL
XFILL_1__11803_ vdd gnd FILL
X_13688_ _13688_/A _13688_/B _13688_/C _13688_/Y vdd gnd OAI21X1
XFILL_0__13232_ vdd gnd FILL
XFILL_0__10444_ vdd gnd FILL
XFILL_1__12783_ vdd gnd FILL
X_12639_ _12639_/A _12639_/B _12639_/C _12639_/Y vdd gnd OAI21X1
XFILL_1__11734_ vdd gnd FILL
XFILL_0__13163_ vdd gnd FILL
XFILL_0__10375_ vdd gnd FILL
XFILL_0__9750_ vdd gnd FILL
XFILL_0__12114_ vdd gnd FILL
XFILL_1__14453_ vdd gnd FILL
X_14309_ _14309_/A _14309_/Y vdd gnd INVX1
XFILL_0__8701_ vdd gnd FILL
XFILL_0__13094_ vdd gnd FILL
X_7240_ _7240_/A _7240_/B _7240_/Y vdd gnd NAND2X1
XFILL_0__9681_ vdd gnd FILL
XFILL_2__9617_ vdd gnd FILL
XFILL_1__13404_ vdd gnd FILL
XFILL_1__10616_ vdd gnd FILL
XFILL_2__12955_ vdd gnd FILL
XFILL_1__14384_ vdd gnd FILL
XFILL_0__12045_ vdd gnd FILL
XFILL_1__11596_ vdd gnd FILL
XFILL_0__8632_ vdd gnd FILL
X_7171_ _7171_/A _7171_/Y vdd gnd INVX8
XFILL_2__9548_ vdd gnd FILL
XFILL_1__13335_ vdd gnd FILL
XFILL_1__10547_ vdd gnd FILL
XFILL_2__12886_ vdd gnd FILL
XFILL_0__8563_ vdd gnd FILL
XFILL_2__9479_ vdd gnd FILL
XFILL_1__13266_ vdd gnd FILL
XFILL_1__10478_ vdd gnd FILL
XFILL_0__7514_ vdd gnd FILL
XFILL_0__13996_ vdd gnd FILL
XFILL_0__8494_ vdd gnd FILL
XCLKBUF1_insert386 CLKBUF1_insert386/A CLKBUF1_insert386/Y vdd gnd CLKBUF1
XFILL_1__12217_ vdd gnd FILL
XFILL_0__12947_ vdd gnd FILL
XFILL_1__13197_ vdd gnd FILL
XFILL_0__7445_ vdd gnd FILL
XFILL_1__12148_ vdd gnd FILL
XFILL_2__14487_ vdd gnd FILL
XFILL_0__12878_ vdd gnd FILL
X_9812_ _9812_/D _9812_/CLK _9812_/Q vdd gnd DFFPOSX1
XFILL_0__7376_ vdd gnd FILL
XFILL_0__14617_ vdd gnd FILL
XFILL_1__12079_ vdd gnd FILL
XFILL_0__11829_ vdd gnd FILL
XFILL_0__9115_ vdd gnd FILL
X_9743_ _9743_/A _9743_/B _9743_/C _9743_/Y vdd gnd OAI21X1
XFILL_0__9046_ vdd gnd FILL
X_9674_ _9674_/A _9674_/B _9674_/Y vdd gnd AND2X2
XFILL_0__14479_ vdd gnd FILL
X_8625_ _8625_/A _8625_/B _8625_/Y vdd gnd OR2X2
XFILL_1__8810_ vdd gnd FILL
X_8556_ _8556_/A _8556_/B _8556_/Y vdd gnd NAND2X1
X_7507_ _7507_/A _7507_/B _7507_/C _7507_/Y vdd gnd OAI21X1
XFILL_0__9948_ vdd gnd FILL
XFILL_1__8741_ vdd gnd FILL
X_8487_ _8487_/A _8487_/B _8487_/Y vdd gnd NAND2X1
X_7438_ _7438_/A _7438_/B _7438_/Y vdd gnd NAND2X1
XFILL_0__9879_ vdd gnd FILL
XFILL_1__8672_ vdd gnd FILL
XFILL_1__7623_ vdd gnd FILL
X_7369_ _7369_/A _7369_/B _7369_/C _7369_/Y vdd gnd OAI21X1
X_9108_ _9108_/A _9108_/B _9108_/Y vdd gnd NAND2X1
XFILL_1__7554_ vdd gnd FILL
X_9039_ _9039_/A _9039_/B _9039_/S _9039_/Y vdd gnd MUX2X1
XFILL_1__7485_ vdd gnd FILL
XFILL_1__9224_ vdd gnd FILL
X_12990_ _12990_/A _12990_/B _12990_/Y vdd gnd NAND2X1
X_11941_ _11941_/A _11941_/Y vdd gnd INVX1
XFILL_1__9155_ vdd gnd FILL
X_14660_ _14660_/A _14660_/B _14660_/Y vdd gnd AND2X2
XFILL_1__8106_ vdd gnd FILL
X_11872_ _11872_/A _11872_/Y vdd gnd INVX1
XFILL_1__9086_ vdd gnd FILL
X_13611_ _13611_/A _13611_/Y vdd gnd INVX1
X_10823_ _10823_/A _10823_/B _10823_/C _10823_/Y vdd gnd OAI21X1
X_14591_ _14591_/A _14591_/B _14591_/Y vdd gnd NAND2X1
XFILL_1__8037_ vdd gnd FILL
X_13542_ _13542_/A _13542_/B _13542_/C _13542_/D _13542_/Y vdd gnd AOI22X1
X_10754_ _10754_/D _10754_/CLK _10754_/Q vdd gnd DFFPOSX1
XFILL_2__7801_ vdd gnd FILL
X_10685_ _10685_/A _10685_/B _10685_/C _10685_/Y vdd gnd OAI21X1
X_13473_ _13473_/D _13473_/CLK _13473_/Q vdd gnd DFFPOSX1
XFILL_1__9988_ vdd gnd FILL
X_12424_ _12424_/A _12424_/B _12424_/C _12424_/Y vdd gnd NAND3X1
XFILL_1__8939_ vdd gnd FILL
XFILL_2__7732_ vdd gnd FILL
XFILL_0__10160_ vdd gnd FILL
X_12355_ _12355_/A _12355_/B _12355_/Y vdd gnd NOR2X1
XFILL_2__7663_ vdd gnd FILL
XFILL_1__11450_ vdd gnd FILL
XFILL_0__10091_ vdd gnd FILL
X_11306_ _11306_/A _11306_/B _11306_/C _11306_/Y vdd gnd NAND3X1
X_12286_ _12286_/A _12286_/B _12286_/C _12286_/Y vdd gnd NAND3X1
XFILL_1__10401_ vdd gnd FILL
XFILL_2__7594_ vdd gnd FILL
XFILL_2_BUFX2_insert5 vdd gnd FILL
XFILL_1__11381_ vdd gnd FILL
X_11237_ _11237_/A _11237_/B _11237_/C _11237_/Y vdd gnd OAI21X1
X_14025_ _14025_/A _14025_/B _14025_/Y vdd gnd NAND2X1
XFILL_1__13120_ vdd gnd FILL
XFILL_1__10332_ vdd gnd FILL
XFILL_0__13850_ vdd gnd FILL
XFILL_2__12671_ vdd gnd FILL
X_11168_ _11168_/A _11168_/B _11168_/C _11168_/Y vdd gnd OAI21X1
XFILL_2__9264_ vdd gnd FILL
XFILL_0__12801_ vdd gnd FILL
XFILL_1__13051_ vdd gnd FILL
XFILL_1__10263_ vdd gnd FILL
X_10119_ _10119_/A _10119_/B _10119_/C _10119_/Y vdd gnd OAI21X1
XFILL_0__13781_ vdd gnd FILL
XFILL_0__10993_ vdd gnd FILL
XFILL_1__12002_ vdd gnd FILL
XFILL_2__8215_ vdd gnd FILL
X_11099_ _11099_/A _11099_/Y vdd gnd INVX1
XFILL_2__11553_ vdd gnd FILL
XFILL_2__9195_ vdd gnd FILL
XFILL_0__12732_ vdd gnd FILL
XFILL_1__10194_ vdd gnd FILL
XFILL_0__7230_ vdd gnd FILL
XFILL_2__10504_ vdd gnd FILL
XFILL_2__11484_ vdd gnd FILL
XFILL_0__12663_ vdd gnd FILL
XFILL_0__7161_ vdd gnd FILL
X_14858_ _14858_/A _14858_/B _14858_/C _14858_/Y vdd gnd OAI21X1
XFILL_0__14402_ vdd gnd FILL
XFILL_1__13953_ vdd gnd FILL
X_13809_ _13809_/A _13809_/B _13809_/C _13809_/Y vdd gnd OAI21X1
XFILL_0__7092_ vdd gnd FILL
X_14789_ _14789_/A _14789_/B _14789_/C _14789_/Y vdd gnd AOI21X1
XFILL_1__12904_ vdd gnd FILL
XFILL_0__14333_ vdd gnd FILL
XFILL_0__11545_ vdd gnd FILL
XFILL_1__13884_ vdd gnd FILL
XFILL_2__12105_ vdd gnd FILL
XFILL_0__14264_ vdd gnd FILL
XFILL_1__12835_ vdd gnd FILL
X_8410_ _8410_/A _8410_/B _8410_/C _8410_/Y vdd gnd AOI21X1
XFILL_0__11476_ vdd gnd FILL
X_9390_ _9390_/A _9390_/B _9390_/C _9390_/Y vdd gnd NAND3X1
XFILL_2__12036_ vdd gnd FILL
XFILL_0__13215_ vdd gnd FILL
XFILL_0__10427_ vdd gnd FILL
XFILL_2__8979_ vdd gnd FILL
XFILL_1__12766_ vdd gnd FILL
X_8341_ _8341_/A _8341_/B _8341_/C _8341_/D _8341_/Y vdd gnd AOI22X1
XFILL_1__11717_ vdd gnd FILL
XFILL_0__13146_ vdd gnd FILL
XFILL_0__10358_ vdd gnd FILL
XFILL_1__12697_ vdd gnd FILL
XFILL_0__9733_ vdd gnd FILL
X_8272_ _8272_/A _8272_/Y vdd gnd INVX1
XFILL_1__14436_ vdd gnd FILL
XFILL_2__13987_ vdd gnd FILL
XFILL_0__13077_ vdd gnd FILL
XFILL_0__10289_ vdd gnd FILL
X_7223_ _7223_/A _7223_/B _7223_/Y vdd gnd OR2X2
XFILL_0__9664_ vdd gnd FILL
XFILL_2__12938_ vdd gnd FILL
XFILL_1__14367_ vdd gnd FILL
XFILL_0__12028_ vdd gnd FILL
XFILL_1__11579_ vdd gnd FILL
XFILL_0__8615_ vdd gnd FILL
X_7154_ _7154_/A _7154_/Y vdd gnd INVX2
XFILL_0__9595_ vdd gnd FILL
XFILL_1__13318_ vdd gnd FILL
XFILL_1__14298_ vdd gnd FILL
XFILL_2__12869_ vdd gnd FILL
XFILL_0__8546_ vdd gnd FILL
XFILL_2__14608_ vdd gnd FILL
X_7085_ _7085_/A _7085_/B _7085_/C _7085_/D _7085_/Y vdd gnd AOI22X1
XFILL_1__13249_ vdd gnd FILL
XFILL_0__13979_ vdd gnd FILL
XFILL_1__7270_ vdd gnd FILL
XFILL_0__8477_ vdd gnd FILL
XFILL_0__7428_ vdd gnd FILL
XFILL_0__7359_ vdd gnd FILL
X_7987_ _7987_/D _7987_/CLK _7987_/Q vdd gnd DFFPOSX1
X_9726_ _9726_/A _9726_/B _9726_/Y vdd gnd NAND2X1
XFILL_0__9029_ vdd gnd FILL
XFILL_1__9911_ vdd gnd FILL
X_9657_ _9657_/A _9657_/B _9657_/C _9657_/Y vdd gnd OAI21X1
X_8608_ _8608_/A _8608_/B _8608_/C _8608_/Y vdd gnd OAI21X1
X_9588_ _9588_/A _9588_/B _9588_/C _9588_/Y vdd gnd OAI21X1
X_10470_ _10470_/A _10470_/B _10470_/C _10470_/Y vdd gnd OAI21X1
X_8539_ _8539_/A _8539_/B _8539_/Y vdd gnd NOR2X1
XFILL_1__8724_ vdd gnd FILL
X_12140_ _12140_/A _12140_/B _12140_/C _12140_/Y vdd gnd OAI21X1
XFILL_1__8655_ vdd gnd FILL
X_12071_ _12071_/A _12071_/B _12071_/Y vdd gnd NAND2X1
XFILL_1__7606_ vdd gnd FILL
XFILL_1__8586_ vdd gnd FILL
X_11022_ _11022_/A _11022_/B _11022_/C _11022_/Y vdd gnd OAI21X1
XFILL_1__7537_ vdd gnd FILL
XFILL_1__7468_ vdd gnd FILL
XFILL_1__9207_ vdd gnd FILL
XFILL_2__8000_ vdd gnd FILL
X_12973_ _12973_/A _12973_/B _12973_/Y vdd gnd NAND2X1
XFILL_1__7399_ vdd gnd FILL
X_14712_ _14712_/A _14712_/B _14712_/C _14712_/Y vdd gnd OAI21X1
X_11924_ _11924_/A _11924_/B _11924_/C _11924_/Y vdd gnd OAI21X1
XFILL_1__9138_ vdd gnd FILL
X_14643_ _14643_/A _14643_/B _14643_/Y vdd gnd NOR2X1
XFILL_2__10220_ vdd gnd FILL
X_11855_ _11855_/A _11855_/Y vdd gnd INVX1
XFILL_1__9069_ vdd gnd FILL
XFILL_1__10950_ vdd gnd FILL
X_10806_ _10806_/A _10806_/B _10806_/C _10806_/Y vdd gnd OAI21X1
X_14574_ _14574_/A _14574_/Y vdd gnd INVX1
XFILL_2__10151_ vdd gnd FILL
X_11786_ _11786_/A _11786_/B _11786_/C _11786_/Y vdd gnd NAND3X1
XFILL_0__11330_ vdd gnd FILL
XFILL_1__10881_ vdd gnd FILL
X_13525_ _13525_/A _13525_/B _13525_/C _13525_/Y vdd gnd OAI21X1
X_10737_ _10737_/D _10737_/CLK _10737_/Q vdd gnd DFFPOSX1
XFILL_1__12620_ vdd gnd FILL
XFILL_2__10082_ vdd gnd FILL
XFILL_0__11261_ vdd gnd FILL
X_13456_ _13456_/D _13456_/CLK _13456_/Q vdd gnd DFFPOSX1
X_10668_ _10668_/A _10668_/B _10668_/C _10668_/Y vdd gnd OAI21X1
XFILL_0__13000_ vdd gnd FILL
XFILL_0__10212_ vdd gnd FILL
X_12407_ _12407_/A _12407_/B _12407_/Y vdd gnd NOR2X1
XFILL_0__11192_ vdd gnd FILL
XFILL_2__7715_ vdd gnd FILL
X_10599_ _10599_/A _10599_/B _10599_/C _10599_/Y vdd gnd OAI21X1
XFILL_1__11502_ vdd gnd FILL
X_13387_ _13387_/A _13387_/B _13387_/C _13387_/Y vdd gnd OAI21X1
XFILL_0__10143_ vdd gnd FILL
XFILL_1__12482_ vdd gnd FILL
X_12338_ _12338_/A _12338_/B _12338_/Y vdd gnd NAND2X1
XFILL_1__14221_ vdd gnd FILL
XFILL_2__7646_ vdd gnd FILL
XFILL_1__11433_ vdd gnd FILL
XFILL_2__10984_ vdd gnd FILL
XFILL_0__10074_ vdd gnd FILL
X_12269_ _12269_/A _12269_/B _12269_/Y vdd gnd NAND2X1
XFILL_1__14152_ vdd gnd FILL
XFILL_2__7577_ vdd gnd FILL
XFILL_0__13902_ vdd gnd FILL
XFILL_1__11364_ vdd gnd FILL
X_14008_ _14008_/A _14008_/B _14008_/C _14008_/Y vdd gnd OAI21X1
XFILL_0__8400_ vdd gnd FILL
XFILL_1__13103_ vdd gnd FILL
XFILL_0__9380_ vdd gnd FILL
XFILL_1__10315_ vdd gnd FILL
XFILL_1__14083_ vdd gnd FILL
XFILL_0__13833_ vdd gnd FILL
XFILL_1__11295_ vdd gnd FILL
XFILL_0__8331_ vdd gnd FILL
XFILL_1__13034_ vdd gnd FILL
XFILL_1__10246_ vdd gnd FILL
XFILL_0__13764_ vdd gnd FILL
XFILL_0__10976_ vdd gnd FILL
X_7910_ _7910_/A _7910_/B _7910_/C _7910_/Y vdd gnd OAI21X1
XFILL_0__8262_ vdd gnd FILL
X_8890_ _8890_/D _8890_/CLK _8890_/Q vdd gnd DFFPOSX1
XFILL_0__12715_ vdd gnd FILL
XFILL_1__10177_ vdd gnd FILL
XFILL_0__13695_ vdd gnd FILL
XFILL_0__7213_ vdd gnd FILL
X_7841_ _7841_/A _7841_/B _7841_/C _7841_/Y vdd gnd OAI21X1
XFILL_0__8193_ vdd gnd FILL
XFILL_2__8129_ vdd gnd FILL
XFILL_0__12646_ vdd gnd FILL
XFILL_0__7144_ vdd gnd FILL
X_7772_ _7772_/A _7772_/B _7772_/Y vdd gnd NAND2X1
XFILL_2__10418_ vdd gnd FILL
XFILL_1__13936_ vdd gnd FILL
X_9511_ _9511_/A _9511_/B _9511_/C _9511_/Y vdd gnd OAI21X1
XFILL_0__7075_ vdd gnd FILL
XFILL_2__10349_ vdd gnd FILL
XFILL_0__14316_ vdd gnd FILL
XFILL_0__11528_ vdd gnd FILL
XFILL_1__13867_ vdd gnd FILL
X_9442_ _9442_/A _9442_/B _9442_/C _9442_/Y vdd gnd OAI21X1
XFILL_0__14247_ vdd gnd FILL
XFILL_1__12818_ vdd gnd FILL
XFILL_0__11459_ vdd gnd FILL
XFILL_1__13798_ vdd gnd FILL
X_9373_ _9373_/A _9373_/B _9373_/Y vdd gnd OR2X2
XFILL_0_BUFX2_insert290 vdd gnd FILL
XFILL_1__12749_ vdd gnd FILL
X_8324_ _8324_/A _8324_/B _8324_/Y vdd gnd NAND2X1
XFILL_0__13129_ vdd gnd FILL
XFILL_0__9716_ vdd gnd FILL
X_8255_ _8255_/A _8255_/B _8255_/Y vdd gnd NOR2X1
XFILL_1__14419_ vdd gnd FILL
X_7206_ _7206_/A _7206_/B _7206_/C _7206_/Y vdd gnd OAI21X1
XFILL_0__9647_ vdd gnd FILL
XFILL_1__8440_ vdd gnd FILL
X_8186_ _8186_/A _8186_/B _8186_/Y vdd gnd NAND2X1
X_7137_ _7137_/A _7137_/Y vdd gnd INVX1
XFILL_0__9578_ vdd gnd FILL
XFILL_1__8371_ vdd gnd FILL
XFILL_1__7322_ vdd gnd FILL
XFILL_0__8529_ vdd gnd FILL
XFILL_1__7253_ vdd gnd FILL
XFILL_1__7184_ vdd gnd FILL
X_11640_ _11640_/D _11640_/CLK _11640_/Q vdd gnd DFFPOSX1
X_9709_ _9709_/A _9709_/B _9709_/C _9709_/Y vdd gnd OAI21X1
X_11571_ _11571_/A _11571_/B _11571_/C _11571_/Y vdd gnd OAI21X1
X_13310_ _13310_/A _13310_/B _13310_/Y vdd gnd NAND2X1
X_10522_ _10522_/A _10522_/B _10522_/C _10522_/Y vdd gnd OAI21X1
X_14290_ _14290_/A _14290_/B _14290_/Y vdd gnd NOR2X1
X_10453_ _10453_/A _10453_/B _10453_/Y vdd gnd NOR2X1
X_13241_ _13241_/A _13241_/B _13241_/C _13241_/Y vdd gnd OAI21X1
XFILL_1__9756_ vdd gnd FILL
X_13172_ _13172_/A _13172_/Y vdd gnd INVX1
X_10384_ _10384_/A _10384_/B _10384_/C _10384_/Y vdd gnd NAND3X1
XFILL_1__8707_ vdd gnd FILL
XFILL_1__9687_ vdd gnd FILL
X_12123_ _12123_/A _12123_/B _12123_/Y vdd gnd NOR2X1
XFILL_1__8638_ vdd gnd FILL
X_12054_ _12054_/A _12054_/B _12054_/Y vdd gnd NAND2X1
XFILL_2__7362_ vdd gnd FILL
XFILL_1__8569_ vdd gnd FILL
X_11005_ _11005_/A _11005_/B _11005_/C _11005_/Y vdd gnd NAND3X1
XFILL_0_CLKBUF1_insert34 vdd gnd FILL
XFILL_1__10100_ vdd gnd FILL
XFILL_0_CLKBUF1_insert45 vdd gnd FILL
XFILL_1__11080_ vdd gnd FILL
XFILL_2__7293_ vdd gnd FILL
XFILL_0_CLKBUF1_insert56 vdd gnd FILL
XFILL_0__10830_ vdd gnd FILL
XFILL_0_CLKBUF1_insert67 vdd gnd FILL
XFILL_0_CLKBUF1_insert78 vdd gnd FILL
XFILL_0_CLKBUF1_insert89 vdd gnd FILL
XFILL_2_BUFX2_insert330 vdd gnd FILL
XFILL_1__10031_ vdd gnd FILL
XFILL_2__12370_ vdd gnd FILL
XFILL_2_BUFX2_insert341 vdd gnd FILL
XFILL_2_BUFX2_insert363 vdd gnd FILL
X_12956_ _12956_/A _12956_/Y vdd gnd INVX1
XFILL_0__12500_ vdd gnd FILL
X_11907_ _11907_/A _11907_/B _11907_/C _11907_/Y vdd gnd NAND3X1
X_12887_ _12887_/A _12887_/B _12887_/C _12887_/Y vdd gnd OAI21X1
XFILL_0__12431_ vdd gnd FILL
XFILL_1__14770_ vdd gnd FILL
XFILL_1__11982_ vdd gnd FILL
X_14626_ _14626_/A _14626_/B _14626_/C _14626_/Y vdd gnd OAI21X1
XFILL_2__10203_ vdd gnd FILL
X_11838_ _11838_/A _11838_/B _11838_/C _11838_/Y vdd gnd OAI21X1
XFILL_1__10933_ vdd gnd FILL
XFILL_1__13721_ vdd gnd FILL
XFILL_0__12362_ vdd gnd FILL
X_14557_ _14557_/A _14557_/Y vdd gnd INVX1
XFILL_2__10134_ vdd gnd FILL
X_11769_ _11769_/A _11769_/B _11769_/Y vdd gnd NOR2X1
XFILL_0__14101_ vdd gnd FILL
XBUFX2_insert340 BUFX2_insert340/A BUFX2_insert340/Y vdd gnd BUFX2
XFILL_0__11313_ vdd gnd FILL
XFILL_1__13652_ vdd gnd FILL
XFILL_1__10864_ vdd gnd FILL
XBUFX2_insert351 BUFX2_insert351/A BUFX2_insert351/Y vdd gnd BUFX2
XBUFX2_insert362 BUFX2_insert362/A BUFX2_insert362/Y vdd gnd BUFX2
XFILL_0__7900_ vdd gnd FILL
XFILL_0__12293_ vdd gnd FILL
X_13508_ _13508_/A _13508_/B _13508_/Y vdd gnd AND2X2
XBUFX2_insert373 BUFX2_insert373/A BUFX2_insert373/Y vdd gnd BUFX2
X_14488_ _14488_/A _14488_/B _14488_/Y vdd gnd NAND2X1
XFILL_2__10065_ vdd gnd FILL
XFILL_0__14032_ vdd gnd FILL
XFILL_0__11244_ vdd gnd FILL
XFILL_1__13583_ vdd gnd FILL
XFILL_1__10795_ vdd gnd FILL
X_13439_ _13439_/D _13439_/CLK _13439_/Q vdd gnd DFFPOSX1
XFILL_0__7831_ vdd gnd FILL
XFILL_1__12534_ vdd gnd FILL
XFILL256350x216150 vdd gnd FILL
XFILL_0__11175_ vdd gnd FILL
XFILL_0__7762_ vdd gnd FILL
XFILL_0__10126_ vdd gnd FILL
XFILL_1__12465_ vdd gnd FILL
XFILL_0__9501_ vdd gnd FILL
X_8040_ _8040_/A _8040_/B _8040_/C _8040_/Y vdd gnd AOI21X1
XFILL_2__7629_ vdd gnd FILL
XFILL_0__7693_ vdd gnd FILL
XFILL_1__11416_ vdd gnd FILL
XFILL_2__10967_ vdd gnd FILL
XFILL_0__10057_ vdd gnd FILL
XFILL_1__12396_ vdd gnd FILL
XFILL_0__9432_ vdd gnd FILL
XFILL_1__11347_ vdd gnd FILL
XFILL_1__14135_ vdd gnd FILL
XFILL_0__14865_ vdd gnd FILL
XFILL_2__10898_ vdd gnd FILL
XFILL_0__9363_ vdd gnd FILL
X_9991_ _9991_/A _9991_/B _9991_/Y vdd gnd NAND2X1
XFILL_1__14066_ vdd gnd FILL
XFILL_1__11278_ vdd gnd FILL
XFILL_0__13816_ vdd gnd FILL
XFILL_0__14796_ vdd gnd FILL
XFILL_0__8314_ vdd gnd FILL
XFILL_0__9294_ vdd gnd FILL
X_8942_ _8942_/A _8942_/B _8942_/C _8942_/D _8942_/Y vdd gnd AOI22X1
XFILL_1__13017_ vdd gnd FILL
XFILL_1__10229_ vdd gnd FILL
XFILL_0__10959_ vdd gnd FILL
XFILL_0__13747_ vdd gnd FILL
XFILL_0__8245_ vdd gnd FILL
X_8873_ _8873_/D _8873_/CLK _8873_/Q vdd gnd DFFPOSX1
XFILL_2__12499_ vdd gnd FILL
XFILL_0__13678_ vdd gnd FILL
X_7824_ _7824_/A _7824_/B _7824_/Y vdd gnd NAND2X1
XFILL_0__8176_ vdd gnd FILL
XFILL_0__12629_ vdd gnd FILL
XFILL_0__7127_ vdd gnd FILL
X_7755_ _7755_/A _7755_/B _7755_/Y vdd gnd NAND2X1
XFILL_1__13919_ vdd gnd FILL
X_7686_ _7686_/A _7686_/B _7686_/C _7686_/Y vdd gnd OAI21X1
X_9425_ _9425_/A _9425_/B _9425_/C _9425_/Y vdd gnd NAND3X1
XFILL_1__7871_ vdd gnd FILL
XFILL_1__9610_ vdd gnd FILL
X_9356_ _9356_/A _9356_/B _9356_/C _9356_/Y vdd gnd OAI21X1
XFILL_1__9541_ vdd gnd FILL
X_8307_ _8307_/A _8307_/Y vdd gnd INVX1
X_9287_ _9287_/A _9287_/B _9287_/Y vdd gnd NOR2X1
X_8238_ _8238_/A _8238_/B _8238_/C _8238_/Y vdd gnd AOI21X1
XFILL_1__9472_ vdd gnd FILL
XFILL_1__8423_ vdd gnd FILL
X_8169_ _8169_/A _8169_/B _8169_/C _8169_/Y vdd gnd OAI21X1
XFILL_1__8354_ vdd gnd FILL
XFILL_1__7305_ vdd gnd FILL
XFILL_1__8285_ vdd gnd FILL
X_12810_ _12810_/A _12810_/B _12810_/Y vdd gnd AND2X2
XFILL_1__7236_ vdd gnd FILL
X_13790_ _13790_/A _13790_/Y vdd gnd INVX1
XFILL_1_BUFX2_insert304 vdd gnd FILL
XFILL_1_BUFX2_insert315 vdd gnd FILL
X_12741_ _12741_/A _12741_/Y vdd gnd INVX1
XFILL_1_BUFX2_insert326 vdd gnd FILL
XFILL_1__7167_ vdd gnd FILL
XFILL_1_BUFX2_insert337 vdd gnd FILL
XFILL_1_BUFX2_insert348 vdd gnd FILL
XFILL_1_BUFX2_insert359 vdd gnd FILL
X_12672_ _12672_/A _12672_/B _12672_/Y vdd gnd NAND2X1
XFILL_1__7098_ vdd gnd FILL
X_14411_ _14411_/A _14411_/B _14411_/Y vdd gnd AND2X2
X_11623_ _11623_/D _11623_/CLK _11623_/Q vdd gnd DFFPOSX1
X_14342_ _14342_/A _14342_/B _14342_/C _14342_/Y vdd gnd NAND3X1
X_11554_ _11554_/A _11554_/B _11554_/C _11554_/Y vdd gnd OAI21X1
X_10505_ _10505_/A _10505_/B _10505_/C _10505_/Y vdd gnd OAI21X1
XFILL_2__8601_ vdd gnd FILL
X_14273_ _14273_/A _14273_/B _14273_/Y vdd gnd OR2X2
X_11485_ _11485_/A _11485_/B _11485_/Y vdd gnd NAND2X1
XFILL_2__9581_ vdd gnd FILL
XFILL_1__10580_ vdd gnd FILL
X_13224_ _13224_/A _13224_/Y vdd gnd INVX1
X_10436_ _10436_/A _10436_/B _10436_/Y vdd gnd NAND2X1
XFILL_1__9739_ vdd gnd FILL
XFILL_2__8532_ vdd gnd FILL
X_13155_ _13155_/A _13155_/B _13155_/C _13155_/D _13155_/Y vdd gnd AOI22X1
X_10367_ _10367_/A _10367_/B _10367_/Y vdd gnd NOR2X1
XFILL_1__12250_ vdd gnd FILL
X_12106_ _12106_/A _12106_/B _12106_/C _12106_/Y vdd gnd AOI21X1
XFILL_0__12980_ vdd gnd FILL
X_13086_ _13086_/A _13086_/B _13086_/Y vdd gnd NAND2X1
X_10298_ _10298_/A _10298_/B _10298_/Y vdd gnd NAND2X1
XFILL_1__11201_ vdd gnd FILL
XFILL_0__11931_ vdd gnd FILL
XFILL_1__12181_ vdd gnd FILL
X_12037_ _12037_/A _12037_/B _12037_/C _12037_/D _12037_/Y vdd gnd AOI22X1
XFILL_1__11132_ vdd gnd FILL
XFILL_0__14650_ vdd gnd FILL
XFILL_0__11862_ vdd gnd FILL
XFILL_2__12422_ vdd gnd FILL
XFILL_0__13601_ vdd gnd FILL
XFILL256350x28950 vdd gnd FILL
XFILL_0__10813_ vdd gnd FILL
XFILL_1__11063_ vdd gnd FILL
XFILL_0__14581_ vdd gnd FILL
XFILL_0__11793_ vdd gnd FILL
XFILL_1__10014_ vdd gnd FILL
XFILL_2_BUFX2_insert160 vdd gnd FILL
X_13988_ _13988_/A _13988_/B _13988_/C _13988_/Y vdd gnd AOI21X1
XFILL_2__12353_ vdd gnd FILL
XFILL_0__13532_ vdd gnd FILL
XFILL_2_BUFX2_insert182 vdd gnd FILL
XFILL_0__8030_ vdd gnd FILL
X_12939_ _12939_/A _12939_/B _12939_/Y vdd gnd NAND2X1
XFILL_1__14822_ vdd gnd FILL
XFILL_2__12284_ vdd gnd FILL
XFILL_0__10675_ vdd gnd FILL
XFILL_2__14023_ vdd gnd FILL
XFILL_0__12414_ vdd gnd FILL
XFILL_1__14753_ vdd gnd FILL
XFILL256950x75750 vdd gnd FILL
X_14609_ _14609_/A _14609_/B _14609_/Y vdd gnd NOR2X1
XFILL_1__11965_ vdd gnd FILL
XFILL_0__13394_ vdd gnd FILL
X_7540_ _7540_/A _7540_/B _7540_/Y vdd gnd NOR2X1
XFILL_0__9981_ vdd gnd FILL
XFILL_1__13704_ vdd gnd FILL
XFILL_0__12345_ vdd gnd FILL
XFILL_1__10916_ vdd gnd FILL
XFILL_1__14684_ vdd gnd FILL
XFILL_0__8932_ vdd gnd FILL
XFILL_1__11896_ vdd gnd FILL
X_7471_ _7471_/A _7471_/B _7471_/C _7471_/Y vdd gnd OAI21X1
XFILL_2__10117_ vdd gnd FILL
XBUFX2_insert170 BUFX2_insert170/A BUFX2_insert170/Y vdd gnd BUFX2
XFILL_1__13635_ vdd gnd FILL
XBUFX2_insert181 BUFX2_insert181/A BUFX2_insert181/Y vdd gnd BUFX2
XFILL_0__12276_ vdd gnd FILL
XFILL_1__10847_ vdd gnd FILL
X_9210_ _9210_/A _9210_/B _9210_/C _9210_/Y vdd gnd NAND3X1
XBUFX2_insert192 BUFX2_insert192/A BUFX2_insert192/Y vdd gnd BUFX2
XFILL_2__10048_ vdd gnd FILL
XFILL_0__14015_ vdd gnd FILL
XFILL_0__11227_ vdd gnd FILL
XFILL_1__10778_ vdd gnd FILL
XFILL_1__13566_ vdd gnd FILL
X_9141_ _9141_/A _9141_/Y vdd gnd INVX1
XFILL_0__7814_ vdd gnd FILL
XFILL_0__8794_ vdd gnd FILL
XFILL_1__12517_ vdd gnd FILL
XFILL_0__11158_ vdd gnd FILL
X_9072_ _9072_/A _9072_/B _9072_/Y vdd gnd NOR2X1
XFILL_0__7745_ vdd gnd FILL
XFILL_0__10109_ vdd gnd FILL
XFILL_1__12448_ vdd gnd FILL
X_8023_ _8023_/A _8023_/Y vdd gnd INVX1
XFILL_0__11089_ vdd gnd FILL
XFILL_0__7676_ vdd gnd FILL
XFILL_0__14917_ vdd gnd FILL
XFILL_1__12379_ vdd gnd FILL
XFILL_0__9415_ vdd gnd FILL
XFILL_1__14118_ vdd gnd FILL
XFILL_0__14848_ vdd gnd FILL
XFILL_0__9346_ vdd gnd FILL
X_9974_ _9974_/A _9974_/B _9974_/C _9974_/Y vdd gnd AOI21X1
XFILL_1__14049_ vdd gnd FILL
XFILL_0__14779_ vdd gnd FILL
XFILL_0__9277_ vdd gnd FILL
X_8925_ _8925_/A _8925_/Y vdd gnd INVX4
XFILL_1__8070_ vdd gnd FILL
XFILL_0__8228_ vdd gnd FILL
X_8856_ _8856_/D _8856_/CLK _8856_/Q vdd gnd DFFPOSX1
X_7807_ _7807_/A _7807_/B _7807_/Y vdd gnd NAND2X1
XFILL_0__8159_ vdd gnd FILL
X_8787_ _8787_/A _8787_/B _8787_/C _8787_/Y vdd gnd OAI21X1
XFILL_1__8972_ vdd gnd FILL
X_7738_ _7738_/A _7738_/B _7738_/C _7738_/Y vdd gnd AOI21X1
X_7669_ _7669_/A _7669_/B _7669_/C _7669_/Y vdd gnd OAI21X1
X_9408_ _9408_/A _9408_/B _9408_/Y vdd gnd NOR2X1
XFILL_1__7854_ vdd gnd FILL
X_11270_ _11270_/A _11270_/B _11270_/C _11270_/Y vdd gnd AOI21X1
X_9339_ _9339_/A _9339_/B _9339_/C _9339_/Y vdd gnd OAI21X1
XFILL_1__7785_ vdd gnd FILL
X_10221_ _10221_/A _10221_/B _10221_/Y vdd gnd AND2X2
XFILL_1__9524_ vdd gnd FILL
X_10152_ _10152_/A _10152_/Y vdd gnd INVX1
XFILL_1__9455_ vdd gnd FILL
X_10083_ _10083_/A _10083_/B _10083_/Y vdd gnd NAND2X1
XFILL_1__8406_ vdd gnd FILL
XFILL_1__9386_ vdd gnd FILL
X_13911_ _13911_/A _13911_/B _13911_/C _13911_/Y vdd gnd NAND3X1
X_14891_ _14891_/D _14891_/CLK _14891_/Q vdd gnd DFFPOSX1
XFILL_1__8337_ vdd gnd FILL
X_13842_ _13842_/A _13842_/Y vdd gnd INVX1
XFILL_1__8268_ vdd gnd FILL
XFILL_1__7219_ vdd gnd FILL
X_13773_ _13773_/A _13773_/B _13773_/Y vdd gnd NOR2X1
X_10985_ _10985_/A _10985_/Y vdd gnd INVX1
XFILL_1_BUFX2_insert112 vdd gnd FILL
XFILL_1_BUFX2_insert123 vdd gnd FILL
XFILL_1__8199_ vdd gnd FILL
XFILL_1_BUFX2_insert134 vdd gnd FILL
XFILL_1_BUFX2_insert145 vdd gnd FILL
X_12724_ _12724_/A _12724_/B _12724_/C _12724_/Y vdd gnd NAND3X1
XFILL_1_BUFX2_insert156 vdd gnd FILL
XFILL_1_BUFX2_insert167 vdd gnd FILL
XFILL_1_BUFX2_insert178 vdd gnd FILL
XFILL_0__10460_ vdd gnd FILL
XFILL_1_BUFX2_insert189 vdd gnd FILL
X_12655_ _12655_/A _12655_/B _12655_/Y vdd gnd NAND2X1
XFILL_2__11020_ vdd gnd FILL
XFILL_1__11750_ vdd gnd FILL
XFILL_0__10391_ vdd gnd FILL
X_11606_ _11606_/A _11606_/B _11606_/C _11606_/Y vdd gnd OAI21X1
X_12586_ _12586_/D _12586_/CLK _12586_/Q vdd gnd DFFPOSX1
XFILL_0__12130_ vdd gnd FILL
XFILL_2__7894_ vdd gnd FILL
X_14325_ _14325_/A _14325_/B _14325_/Y vdd gnd AND2X2
X_11537_ _11537_/A _11537_/B _11537_/C _11537_/Y vdd gnd OAI21X1
XFILL_1__10632_ vdd gnd FILL
XFILL_1__13420_ vdd gnd FILL
XFILL_0__12061_ vdd gnd FILL
X_14256_ _14256_/A _14256_/B _14256_/C _14256_/Y vdd gnd NAND3X1
XFILL_2__14710_ vdd gnd FILL
X_11468_ _11468_/A _11468_/B _11468_/Y vdd gnd NAND2X1
XFILL_0__11012_ vdd gnd FILL
XFILL_2__11922_ vdd gnd FILL
XFILL_1__10563_ vdd gnd FILL
XFILL_1__13351_ vdd gnd FILL
X_13207_ _13207_/A _13207_/B _13207_/Y vdd gnd NAND2X1
X_10419_ _10419_/A _10419_/B _10419_/C _10419_/Y vdd gnd NAND3X1
XFILL_2__8515_ vdd gnd FILL
X_14187_ _14187_/D _14187_/CLK _14187_/Q vdd gnd DFFPOSX1
XFILL_2__14641_ vdd gnd FILL
XFILL_1__12302_ vdd gnd FILL
X_11399_ _11399_/A _11399_/B _11399_/Y vdd gnd NAND2X1
XFILL_2__11853_ vdd gnd FILL
XFILL_1__13282_ vdd gnd FILL
XFILL_1__10494_ vdd gnd FILL
X_13138_ _13138_/A _13138_/B _13138_/Y vdd gnd NAND2X1
XFILL_0__7530_ vdd gnd FILL
XFILL_2__8446_ vdd gnd FILL
XFILL_1__12233_ vdd gnd FILL
XFILL_2__14572_ vdd gnd FILL
XFILL_2__11784_ vdd gnd FILL
XFILL_0__12963_ vdd gnd FILL
XFILL_0__7461_ vdd gnd FILL
X_13069_ _13069_/A _13069_/B _13069_/Y vdd gnd NAND2X1
XFILL_0__14702_ vdd gnd FILL
XFILL_2__8377_ vdd gnd FILL
XFILL_1__12164_ vdd gnd FILL
XFILL_0__9200_ vdd gnd FILL
XFILL_0__11914_ vdd gnd FILL
XFILL_0__12894_ vdd gnd FILL
XFILL_0__7392_ vdd gnd FILL
XFILL_1__11115_ vdd gnd FILL
XFILL_0__14633_ vdd gnd FILL
XFILL_2__10666_ vdd gnd FILL
XFILL_0__11845_ vdd gnd FILL
XFILL_1__12095_ vdd gnd FILL
XFILL_0__9131_ vdd gnd FILL
XFILL_1__11046_ vdd gnd FILL
XFILL_0__14564_ vdd gnd FILL
XFILL_0__11776_ vdd gnd FILL
XFILL_0__9062_ vdd gnd FILL
X_8710_ _8710_/A _8710_/B _8710_/Y vdd gnd NAND2X1
X_9690_ _9690_/A _9690_/B _9690_/C _9690_/Y vdd gnd OAI21X1
XFILL_2__12336_ vdd gnd FILL
XFILL_0__13515_ vdd gnd FILL
XFILL_0__8013_ vdd gnd FILL
XFILL_0__14495_ vdd gnd FILL
X_8641_ _8641_/A _8641_/B _8641_/Y vdd gnd NOR2X1
XFILL_1__14805_ vdd gnd FILL
XFILL_2__12267_ vdd gnd FILL
XFILL_0__10658_ vdd gnd FILL
XFILL_1__12997_ vdd gnd FILL
XFILL_2__14006_ vdd gnd FILL
X_8572_ _8572_/A _8572_/B _8572_/Y vdd gnd NAND2X1
XFILL_1__14736_ vdd gnd FILL
XFILL_1__11948_ vdd gnd FILL
XFILL_2__12198_ vdd gnd FILL
XFILL_0__13377_ vdd gnd FILL
XFILL_0__10589_ vdd gnd FILL
X_7523_ _7523_/A _7523_/B _7523_/C _7523_/Y vdd gnd NAND3X1
XFILL_0__9964_ vdd gnd FILL
XFILL_0__12328_ vdd gnd FILL
XFILL_1__14667_ vdd gnd FILL
XFILL_1__11879_ vdd gnd FILL
X_7454_ _7454_/A _7454_/B _7454_/C _7454_/Y vdd gnd OAI21X1
XFILL_0__9895_ vdd gnd FILL
XFILL_1__13618_ vdd gnd FILL
XFILL_0__12259_ vdd gnd FILL
XFILL_1__14598_ vdd gnd FILL
X_7385_ _7385_/A _7385_/B _7385_/C _7385_/Y vdd gnd NAND3X1
XFILL_1__13549_ vdd gnd FILL
X_9124_ _9124_/A _9124_/B _9124_/C _9124_/Y vdd gnd AOI21X1
XFILL_1__7570_ vdd gnd FILL
XFILL_0__8777_ vdd gnd FILL
XFILL_2__14839_ vdd gnd FILL
X_9055_ _9055_/A _9055_/B _9055_/Y vdd gnd NAND2X1
XFILL_0__7728_ vdd gnd FILL
XFILL_1__9240_ vdd gnd FILL
X_8006_ _8006_/A _8006_/B _8006_/C _8006_/D _8006_/Y vdd gnd AOI22X1
XFILL_0__7659_ vdd gnd FILL
XFILL_1__9171_ vdd gnd FILL
XFILL_0__9329_ vdd gnd FILL
XFILL_1__8122_ vdd gnd FILL
X_9957_ _9957_/A _9957_/B _9957_/S _9957_/Y vdd gnd MUX2X1
XFILL_1__8053_ vdd gnd FILL
X_8908_ _8908_/D _8908_/CLK _8908_/Q vdd gnd DFFPOSX1
X_9888_ _9888_/A _9888_/B _9888_/C _9888_/Y vdd gnd AOI21X1
X_10770_ _10770_/A _10770_/B _10770_/Y vdd gnd NOR2X1
X_8839_ _8839_/A _8839_/B _8839_/C _8839_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert108 vdd gnd FILL
XFILL_0_BUFX2_insert119 vdd gnd FILL
X_12440_ _12440_/A _12440_/Y vdd gnd INVX1
XFILL_1__8955_ vdd gnd FILL
XFILL_1__7906_ vdd gnd FILL
X_12371_ _12371_/A _12371_/B _12371_/C _12371_/Y vdd gnd OAI21X1
X_14110_ _14110_/A _14110_/Y vdd gnd INVX1
X_11322_ _11322_/A _11322_/Y vdd gnd INVX1
XFILL_1__7837_ vdd gnd FILL
X_14041_ _14041_/A _14041_/B _14041_/C _14041_/Y vdd gnd NAND3X1
X_11253_ _11253_/A _11253_/B _11253_/C _11253_/Y vdd gnd OAI21X1
XFILL_1_CLKBUF1_insert388 vdd gnd FILL
XFILL_1__7768_ vdd gnd FILL
X_10204_ _10204_/A _10204_/B _10204_/C _10204_/Y vdd gnd OAI21X1
XFILL_1__9507_ vdd gnd FILL
XFILL_2__8300_ vdd gnd FILL
X_11184_ _11184_/A _11184_/B _11184_/Y vdd gnd NAND2X1
XFILL_1__7699_ vdd gnd FILL
X_10135_ _10135_/A _10135_/B _10135_/C _10135_/Y vdd gnd NAND3X1
XFILL_1__9438_ vdd gnd FILL
XFILL_2__8231_ vdd gnd FILL
X_10066_ _10066_/A _10066_/B _10066_/Y vdd gnd NAND2X1
XFILL_1__9369_ vdd gnd FILL
XFILL_2__10520_ vdd gnd FILL
XFILL_2__8162_ vdd gnd FILL
X_14874_ _14874_/D _14874_/CLK _14874_/Q vdd gnd DFFPOSX1
XFILL_2__10451_ vdd gnd FILL
XFILL_2__8093_ vdd gnd FILL
X_13825_ _13825_/A _13825_/B _13825_/C _13825_/Y vdd gnd AOI21X1
XFILL_2__13170_ vdd gnd FILL
XFILL_2__10382_ vdd gnd FILL
XFILL_1__12920_ vdd gnd FILL
XFILL_0__11561_ vdd gnd FILL
X_13756_ _13756_/A _13756_/B _13756_/Y vdd gnd NAND2X1
X_10968_ _10968_/A _10968_/B _10968_/Y vdd gnd NOR2X1
XFILL_0__13300_ vdd gnd FILL
XFILL_0__10512_ vdd gnd FILL
XFILL_0__14280_ vdd gnd FILL
XFILL_1__12851_ vdd gnd FILL
XFILL_0__11492_ vdd gnd FILL
X_12707_ _12707_/A _12707_/Y vdd gnd INVX1
X_13687_ _13687_/A _13687_/B _13687_/Y vdd gnd AND2X2
XFILL_1__11802_ vdd gnd FILL
XFILL_0__13231_ vdd gnd FILL
X_10899_ _10899_/A _10899_/B _10899_/C _10899_/Y vdd gnd OAI21X1
XFILL_2__8995_ vdd gnd FILL
XFILL_0__10443_ vdd gnd FILL
XFILL_1__12782_ vdd gnd FILL
X_12638_ _12638_/A _12638_/B _12638_/C _12638_/Y vdd gnd OAI21X1
XFILL_2__11003_ vdd gnd FILL
XFILL_0__13162_ vdd gnd FILL
XFILL_1__11733_ vdd gnd FILL
XFILL_0__10374_ vdd gnd FILL
X_12569_ _12569_/D _12569_/CLK _12569_/Q vdd gnd DFFPOSX1
XFILL_0__12113_ vdd gnd FILL
XFILL_2__7877_ vdd gnd FILL
XFILL_1__14452_ vdd gnd FILL
X_14308_ _14308_/A _14308_/B _14308_/C _14308_/Y vdd gnd OAI21X1
XFILL_0__8700_ vdd gnd FILL
XFILL_0__13093_ vdd gnd FILL
XFILL_0__9680_ vdd gnd FILL
XFILL_1__13403_ vdd gnd FILL
XFILL_1__10615_ vdd gnd FILL
XFILL_0__12044_ vdd gnd FILL
XFILL_1__14383_ vdd gnd FILL
XFILL_1__11595_ vdd gnd FILL
X_14239_ _14239_/A _14239_/B _14239_/C _14239_/Y vdd gnd OAI21X1
XFILL_0__8631_ vdd gnd FILL
X_7170_ _7170_/A _7170_/Y vdd gnd INVX1
XFILL_2__11905_ vdd gnd FILL
XFILL_1__13334_ vdd gnd FILL
XFILL_1__10546_ vdd gnd FILL
XFILL_0__8562_ vdd gnd FILL
XFILL_2__14624_ vdd gnd FILL
XFILL_2__11836_ vdd gnd FILL
XFILL_1__10477_ vdd gnd FILL
XFILL_1__13265_ vdd gnd FILL
XFILL_0__7513_ vdd gnd FILL
XFILL_0__13995_ vdd gnd FILL
XFILL_2__8429_ vdd gnd FILL
XFILL_0__8493_ vdd gnd FILL
XFILL_1__12216_ vdd gnd FILL
XFILL_1__13196_ vdd gnd FILL
XCLKBUF1_insert387 CLKBUF1_insert387/A CLKBUF1_insert387/Y vdd gnd CLKBUF1
XFILL_2__11767_ vdd gnd FILL
XFILL_0__12946_ vdd gnd FILL
XFILL_0__7444_ vdd gnd FILL
XFILL_2__13506_ vdd gnd FILL
XFILL_1__12147_ vdd gnd FILL
XFILL_2__11698_ vdd gnd FILL
X_9811_ _9811_/D _9811_/CLK _9811_/Q vdd gnd DFFPOSX1
XFILL_0__12877_ vdd gnd FILL
XFILL_0__7375_ vdd gnd FILL
XFILL_0__14616_ vdd gnd FILL
XFILL_2__10649_ vdd gnd FILL
XFILL_1__12078_ vdd gnd FILL
XFILL_0__9114_ vdd gnd FILL
XFILL_0__11828_ vdd gnd FILL
X_9742_ _9742_/A _9742_/Y vdd gnd INVX1
XFILL_1__11029_ vdd gnd FILL
XFILL_0__9045_ vdd gnd FILL
XFILL_0__11759_ vdd gnd FILL
X_9673_ _9673_/A _9673_/B _9673_/Y vdd gnd NAND2X1
XFILL_0__14478_ vdd gnd FILL
X_8624_ _8624_/A _8624_/B _8624_/Y vdd gnd OR2X2
X_8555_ _8555_/A _8555_/B _8555_/C _8555_/Y vdd gnd NAND3X1
XFILL_1__14719_ vdd gnd FILL
XFILL_0__9947_ vdd gnd FILL
X_7506_ _7506_/A _7506_/B _7506_/C _7506_/Y vdd gnd OAI21X1
XFILL_1__8740_ vdd gnd FILL
X_8486_ _8486_/A _8486_/B _8486_/C _8486_/Y vdd gnd OAI21X1
X_7437_ _7437_/A _7437_/B _7437_/C _7437_/Y vdd gnd OAI21X1
XFILL_0__9878_ vdd gnd FILL
XFILL_1__8671_ vdd gnd FILL
XFILL_1__7622_ vdd gnd FILL
XFILL_0__8829_ vdd gnd FILL
X_7368_ _7368_/A _7368_/B _7368_/C _7368_/Y vdd gnd AOI21X1
X_9107_ _9107_/A _9107_/Y vdd gnd INVX1
XFILL_1__7553_ vdd gnd FILL
X_7299_ _7299_/A _7299_/Y vdd gnd INVX1
X_9038_ _9038_/A _9038_/B _9038_/S _9038_/Y vdd gnd MUX2X1
XFILL_1__7484_ vdd gnd FILL
XFILL_1__9223_ vdd gnd FILL
X_11940_ _11940_/A _11940_/B _11940_/C _11940_/D _11940_/Y vdd gnd AOI22X1
XFILL_1__9154_ vdd gnd FILL
XFILL_1__8105_ vdd gnd FILL
X_11871_ _11871_/A _11871_/B _11871_/C _11871_/Y vdd gnd AOI21X1
XFILL_1__9085_ vdd gnd FILL
X_13610_ _13610_/A _13610_/B _13610_/C _13610_/Y vdd gnd AOI21X1
X_10822_ _10822_/A _10822_/B _10822_/C _10822_/D _10822_/Y vdd gnd AOI22X1
X_14590_ _14590_/A _14590_/B _14590_/Y vdd gnd NAND2X1
XFILL_1__8036_ vdd gnd FILL
X_13541_ _13541_/A _13541_/B _13541_/C _13541_/Y vdd gnd OAI21X1
X_10753_ _10753_/D _10753_/CLK _10753_/Q vdd gnd DFFPOSX1
X_13472_ _13472_/D _13472_/CLK _13472_/Q vdd gnd DFFPOSX1
X_10684_ _10684_/A _10684_/B _10684_/Y vdd gnd NAND2X1
XFILL_1__9987_ vdd gnd FILL
X_12423_ _12423_/A _12423_/B _12423_/C _12423_/Y vdd gnd AOI21X1
XFILL_1__8938_ vdd gnd FILL
X_12354_ _12354_/A _12354_/B _12354_/C _12354_/Y vdd gnd AOI21X1
XFILL_0__10090_ vdd gnd FILL
X_11305_ _11305_/A _11305_/B _11305_/C _11305_/Y vdd gnd NAND3X1
X_12285_ _12285_/A _12285_/B _12285_/Y vdd gnd OR2X2
XFILL_1__10400_ vdd gnd FILL
XFILL_1__11380_ vdd gnd FILL
X_14024_ _14024_/A _14024_/B _14024_/C _14024_/Y vdd gnd NAND3X1
X_11236_ _11236_/A _11236_/B _11236_/Y vdd gnd NOR2X1
XFILL_1__10331_ vdd gnd FILL
X_11167_ _11167_/A _11167_/B _11167_/C _11167_/Y vdd gnd OAI21X1
XFILL_1__13050_ vdd gnd FILL
XFILL_1__10262_ vdd gnd FILL
XFILL_0__12800_ vdd gnd FILL
XFILL_0__10992_ vdd gnd FILL
X_10118_ _10118_/A _10118_/B _10118_/C _10118_/Y vdd gnd OAI21X1
XFILL_0__13780_ vdd gnd FILL
XFILL_1__12001_ vdd gnd FILL
XFILL_2__14340_ vdd gnd FILL
X_11098_ _11098_/A _11098_/B _11098_/Y vdd gnd NAND2X1
XFILL_1__10193_ vdd gnd FILL
XFILL_0__12731_ vdd gnd FILL
X_10049_ _10049_/A _10049_/B _10049_/C _10049_/Y vdd gnd OAI21X1
XFILL_2__8145_ vdd gnd FILL
XFILL_0__12662_ vdd gnd FILL
XFILL_0__7160_ vdd gnd FILL
X_14857_ _14857_/A _14857_/B _14857_/C _14857_/Y vdd gnd AOI21X1
XFILL_2__13222_ vdd gnd FILL
XFILL_2__10434_ vdd gnd FILL
XFILL_0__14401_ vdd gnd FILL
XFILL_2__8076_ vdd gnd FILL
XFILL_1__13952_ vdd gnd FILL
X_13808_ _13808_/A _13808_/Y vdd gnd INVX1
X_14788_ _14788_/A _14788_/B _14788_/C _14788_/Y vdd gnd NAND3X1
XFILL_0__7091_ vdd gnd FILL
XFILL_2__13153_ vdd gnd FILL
XFILL_1__12903_ vdd gnd FILL
XFILL_2__10365_ vdd gnd FILL
XFILL_0__14332_ vdd gnd FILL
XFILL_0__11544_ vdd gnd FILL
XFILL_1__13883_ vdd gnd FILL
X_13739_ _13739_/A _13739_/B _13739_/C _13739_/Y vdd gnd AOI21X1
XFILL_2__13084_ vdd gnd FILL
XFILL_1__12834_ vdd gnd FILL
XFILL_2__10296_ vdd gnd FILL
XFILL_0__14263_ vdd gnd FILL
XFILL_0__11475_ vdd gnd FILL
XFILL_0__13214_ vdd gnd FILL
XFILL_0__10426_ vdd gnd FILL
XFILL256650x72150 vdd gnd FILL
XFILL_1__12765_ vdd gnd FILL
X_8340_ _8340_/A _8340_/B _8340_/Y vdd gnd OR2X2
XFILL_0__13145_ vdd gnd FILL
XFILL_1__11716_ vdd gnd FILL
XFILL_0__10357_ vdd gnd FILL
XFILL_0__9732_ vdd gnd FILL
XFILL_1__12696_ vdd gnd FILL
X_8271_ _8271_/A _8271_/B _8271_/C _8271_/Y vdd gnd OAI21X1
XFILL_1__14435_ vdd gnd FILL
XFILL_0__13076_ vdd gnd FILL
XFILL_0__10288_ vdd gnd FILL
X_7222_ _7222_/A _7222_/Y vdd gnd INVX1
XFILL_0__9663_ vdd gnd FILL
XFILL_0__12027_ vdd gnd FILL
XFILL_1__14366_ vdd gnd FILL
XFILL_0__8614_ vdd gnd FILL
XFILL_1__11578_ vdd gnd FILL
X_7153_ _7153_/A _7153_/B _7153_/C _7153_/Y vdd gnd OAI21X1
XFILL_0__9594_ vdd gnd FILL
XFILL_1__13317_ vdd gnd FILL
XFILL_1__10529_ vdd gnd FILL
XFILL_1__14297_ vdd gnd FILL
XFILL_0__8545_ vdd gnd FILL
X_7084_ _7084_/A _7084_/B _7084_/Y vdd gnd NOR2X1
XFILL_2__11819_ vdd gnd FILL
XFILL_1__13248_ vdd gnd FILL
XFILL_0__13978_ vdd gnd FILL
XFILL_0__8476_ vdd gnd FILL
XFILL_0__12929_ vdd gnd FILL
XFILL_1__13179_ vdd gnd FILL
XFILL_0__7427_ vdd gnd FILL
XFILL_0__7358_ vdd gnd FILL
X_7986_ _7986_/D _7986_/CLK _7986_/Q vdd gnd DFFPOSX1
X_9725_ _9725_/A _9725_/B _9725_/C _9725_/Y vdd gnd OAI21X1
XFILL_0__7289_ vdd gnd FILL
XFILL_0__9028_ vdd gnd FILL
XFILL_1__9910_ vdd gnd FILL
X_9656_ _9656_/A _9656_/B _9656_/Y vdd gnd NAND2X1
X_8607_ _8607_/A _8607_/B _8607_/C _8607_/Y vdd gnd OAI21X1
X_9587_ _9587_/A _9587_/B _9587_/C _9587_/Y vdd gnd OAI21X1
X_8538_ _8538_/A _8538_/B _8538_/C _8538_/Y vdd gnd OAI21X1
XFILL_1__8723_ vdd gnd FILL
X_8469_ _8469_/A _8469_/B _8469_/C _8469_/Y vdd gnd NAND3X1
XFILL_1__8654_ vdd gnd FILL
XFILL_1__7605_ vdd gnd FILL
X_12070_ _12070_/A _12070_/B _12070_/Y vdd gnd NOR2X1
XFILL_1__8585_ vdd gnd FILL
X_11021_ _11021_/A _11021_/B _11021_/C _11021_/Y vdd gnd AOI21X1
XFILL_1__7536_ vdd gnd FILL
XFILL_1__7467_ vdd gnd FILL
XFILL_1__9206_ vdd gnd FILL
X_12972_ _12972_/A _12972_/Y vdd gnd INVX1
XFILL_1__7398_ vdd gnd FILL
X_14711_ _14711_/A _14711_/B _14711_/Y vdd gnd NOR2X1
XFILL257550x57750 vdd gnd FILL
X_11923_ _11923_/A _11923_/B _11923_/Y vdd gnd NAND2X1
XFILL_1__9137_ vdd gnd FILL
X_14642_ _14642_/A _14642_/B _14642_/Y vdd gnd NAND2X1
X_11854_ _11854_/A _11854_/Y vdd gnd INVX1
XFILL_1__9068_ vdd gnd FILL
XFILL_2__9950_ vdd gnd FILL
X_10805_ _10805_/A _10805_/B _10805_/Y vdd gnd NAND2X1
X_14573_ _14573_/A _14573_/Y vdd gnd INVX1
XFILL_1__8019_ vdd gnd FILL
X_11785_ _11785_/A _11785_/B _11785_/C _11785_/Y vdd gnd AOI21X1
XFILL_2__9881_ vdd gnd FILL
X_13524_ _13524_/A _13524_/B _13524_/C _13524_/Y vdd gnd OAI21X1
XFILL_1__10880_ vdd gnd FILL
X_10736_ _10736_/D _10736_/CLK _10736_/Q vdd gnd DFFPOSX1
XFILL_2__8832_ vdd gnd FILL
XFILL_0__11260_ vdd gnd FILL
X_13455_ _13455_/D _13455_/CLK _13455_/Q vdd gnd DFFPOSX1
X_10667_ _10667_/A _10667_/B _10667_/C _10667_/Y vdd gnd OAI21X1
XFILL_0__10211_ vdd gnd FILL
XFILL_2__8763_ vdd gnd FILL
X_12406_ _12406_/A _12406_/B _12406_/Y vdd gnd NAND2X1
XFILL_0__11191_ vdd gnd FILL
X_13386_ _13386_/A _13386_/B _13386_/Y vdd gnd NAND2X1
X_10598_ _10598_/A _10598_/B _10598_/Y vdd gnd AND2X2
XFILL_1__11501_ vdd gnd FILL
XFILL_0__10142_ vdd gnd FILL
XFILL_2__8694_ vdd gnd FILL
XFILL_1__12481_ vdd gnd FILL
X_12337_ _12337_/A _12337_/B _12337_/Y vdd gnd NOR2X1
XFILL_1__14220_ vdd gnd FILL
XFILL_1__11432_ vdd gnd FILL
XFILL_0__10073_ vdd gnd FILL
X_12268_ _12268_/A _12268_/B _12268_/Y vdd gnd NAND2X1
XFILL_2__12722_ vdd gnd FILL
XFILL_0__13901_ vdd gnd FILL
XFILL_1__14151_ vdd gnd FILL
X_14007_ _14007_/A _14007_/B _14007_/C _14007_/Y vdd gnd AOI21X1
XFILL_1__11363_ vdd gnd FILL
X_11219_ _11219_/A _11219_/B _11219_/C _11219_/Y vdd gnd NAND3X1
XFILL_2__9315_ vdd gnd FILL
XFILL_1__13102_ vdd gnd FILL
X_12199_ _12199_/A _12199_/Y vdd gnd INVX1
XFILL_1__10314_ vdd gnd FILL
XFILL_1__11294_ vdd gnd FILL
XFILL_0__13832_ vdd gnd FILL
XFILL_1__14082_ vdd gnd FILL
XFILL_0__8330_ vdd gnd FILL
XFILL_2__11604_ vdd gnd FILL
XFILL_1__10245_ vdd gnd FILL
XFILL_1__13033_ vdd gnd FILL
XFILL_0__13763_ vdd gnd FILL
XFILL_0__10975_ vdd gnd FILL
XFILL_0__8261_ vdd gnd FILL
XFILL_2__14323_ vdd gnd FILL
XFILL_1__10176_ vdd gnd FILL
XFILL_0__12714_ vdd gnd FILL
XFILL_0__7212_ vdd gnd FILL
X_14909_ _14909_/A _14909_/Y vdd gnd BUFX2
XFILL_0__13694_ vdd gnd FILL
X_7840_ _7840_/A _7840_/B _7840_/Y vdd gnd OR2X2
XFILL_0__8192_ vdd gnd FILL
XFILL_2__14254_ vdd gnd FILL
XFILL_0__12645_ vdd gnd FILL
XFILL_0__7143_ vdd gnd FILL
XFILL_2__13205_ vdd gnd FILL
X_7771_ _7771_/A _7771_/B _7771_/C _7771_/Y vdd gnd OAI21X1
XFILL_1__13935_ vdd gnd FILL
X_9510_ _9510_/A _9510_/B _9510_/Y vdd gnd OR2X2
XFILL_0__7074_ vdd gnd FILL
XFILL_2__13136_ vdd gnd FILL
XFILL_0__14315_ vdd gnd FILL
XFILL_1__13866_ vdd gnd FILL
XFILL_0__11527_ vdd gnd FILL
X_9441_ _9441_/A _9441_/B _9441_/C _9441_/Y vdd gnd AOI21X1
XFILL_1__12817_ vdd gnd FILL
XFILL_2__13067_ vdd gnd FILL
XFILL_0__14246_ vdd gnd FILL
XFILL_0__11458_ vdd gnd FILL
XFILL_1__13797_ vdd gnd FILL
X_9372_ _9372_/A _9372_/B _9372_/Y vdd gnd NAND2X1
XFILL_0__10409_ vdd gnd FILL
XFILL_1__12748_ vdd gnd FILL
XFILL_0_BUFX2_insert280 vdd gnd FILL
XFILL_0__11389_ vdd gnd FILL
XFILL_0_BUFX2_insert291 vdd gnd FILL
X_8323_ _8323_/A _8323_/B _8323_/Y vdd gnd NAND2X1
XFILL_0__13128_ vdd gnd FILL
XFILL_1__12679_ vdd gnd FILL
XFILL_0__9715_ vdd gnd FILL
X_8254_ _8254_/A _8254_/Y vdd gnd INVX1
XFILL_1__14418_ vdd gnd FILL
XFILL_0__13059_ vdd gnd FILL
X_7205_ _7205_/A _7205_/B _7205_/Y vdd gnd NAND2X1
XFILL_0__9646_ vdd gnd FILL
X_8185_ _8185_/A _8185_/B _8185_/C _8185_/Y vdd gnd OAI21X1
XFILL_1__14349_ vdd gnd FILL
X_7136_ _7136_/A _7136_/B _7136_/C _7136_/Y vdd gnd OAI21X1
XFILL_0__9577_ vdd gnd FILL
XFILL_1__8370_ vdd gnd FILL
XFILL_1__7321_ vdd gnd FILL
XFILL_0__8528_ vdd gnd FILL
XFILL_1__7252_ vdd gnd FILL
XFILL_0__8459_ vdd gnd FILL
XFILL_1__7183_ vdd gnd FILL
X_7969_ _7969_/D _7969_/CLK _7969_/Q vdd gnd DFFPOSX1
X_9708_ _9708_/A _9708_/B _9708_/Y vdd gnd NAND2X1
X_11570_ _11570_/A _11570_/B _11570_/Y vdd gnd NAND2X1
X_9639_ _9639_/A _9639_/B _9639_/Y vdd gnd OR2X2
X_10521_ _10521_/A _10521_/Y vdd gnd INVX1
X_13240_ _13240_/A _13240_/Y vdd gnd INVX1
X_10452_ _10452_/A _10452_/B _10452_/C _10452_/Y vdd gnd AOI21X1
XFILL_1__9755_ vdd gnd FILL
XFILL257550x32550 vdd gnd FILL
X_13171_ _13171_/A _13171_/B _13171_/C _13171_/Y vdd gnd OAI21X1
X_10383_ _10383_/A _10383_/B _10383_/Y vdd gnd NAND2X1
XFILL_1__8706_ vdd gnd FILL
XFILL_1__9686_ vdd gnd FILL
X_12122_ _12122_/A _12122_/B _12122_/C _12122_/Y vdd gnd AOI21X1
XFILL_1__8637_ vdd gnd FILL
X_12053_ _12053_/A _12053_/B _12053_/Y vdd gnd NAND2X1
XFILL_1__8568_ vdd gnd FILL
X_11004_ _11004_/A _11004_/B _11004_/Y vdd gnd NAND2X1
XFILL_2__9100_ vdd gnd FILL
XFILL_1__7519_ vdd gnd FILL
XFILL_0_CLKBUF1_insert35 vdd gnd FILL
XFILL_0_CLKBUF1_insert46 vdd gnd FILL
XFILL_1__8499_ vdd gnd FILL
XFILL_0_CLKBUF1_insert57 vdd gnd FILL
XFILL_2__9031_ vdd gnd FILL
XFILL_0_CLKBUF1_insert68 vdd gnd FILL
XFILL_2_BUFX2_insert320 vdd gnd FILL
XFILL_0_CLKBUF1_insert79 vdd gnd FILL
XFILL_1__10030_ vdd gnd FILL
XFILL_2_BUFX2_insert353 vdd gnd FILL
X_12955_ _12955_/A _12955_/B _12955_/Y vdd gnd NAND2X1
XFILL_2__11320_ vdd gnd FILL
XFILL_2_BUFX2_insert375 vdd gnd FILL
X_11906_ _11906_/A _11906_/B _11906_/C _11906_/Y vdd gnd OAI21X1
X_12886_ _12886_/A _12886_/B _12886_/C _12886_/Y vdd gnd OAI21X1
XFILL_2__11251_ vdd gnd FILL
XFILL_0__12430_ vdd gnd FILL
XFILL_1__11981_ vdd gnd FILL
X_14625_ _14625_/A _14625_/B _14625_/C _14625_/Y vdd gnd AOI21X1
X_11837_ _11837_/A _11837_/Y vdd gnd INVX1
XFILL_2__9933_ vdd gnd FILL
XFILL_1__13720_ vdd gnd FILL
XFILL_0__12361_ vdd gnd FILL
XFILL_1__10932_ vdd gnd FILL
XFILL_2__11182_ vdd gnd FILL
X_14556_ _14556_/A _14556_/Y vdd gnd INVX1
X_11768_ _11768_/A _11768_/B _11768_/S _11768_/Y vdd gnd MUX2X1
XFILL_0__14100_ vdd gnd FILL
XFILL_0__11312_ vdd gnd FILL
XBUFX2_insert330 BUFX2_insert330/A BUFX2_insert330/Y vdd gnd BUFX2
XFILL_2__9864_ vdd gnd FILL
XFILL_1__13651_ vdd gnd FILL
XBUFX2_insert341 BUFX2_insert341/A BUFX2_insert341/Y vdd gnd BUFX2
XFILL_0__12292_ vdd gnd FILL
XFILL_1__10863_ vdd gnd FILL
X_10719_ _10719_/D _10719_/CLK _10719_/Q vdd gnd DFFPOSX1
X_13507_ _13507_/A _13507_/Y vdd gnd INVX1
XBUFX2_insert352 BUFX2_insert352/A BUFX2_insert352/Y vdd gnd BUFX2
XBUFX2_insert363 BUFX2_insert363/A BUFX2_insert363/Y vdd gnd BUFX2
X_14487_ _14487_/A _14487_/B _14487_/C _14487_/Y vdd gnd OAI21X1
XFILL_2__8815_ vdd gnd FILL
XBUFX2_insert374 BUFX2_insert374/A BUFX2_insert374/Y vdd gnd BUFX2
X_11699_ _11699_/A _11699_/B _11699_/C _11699_/Y vdd gnd OAI21X1
XFILL_0__11243_ vdd gnd FILL
XFILL_0__14031_ vdd gnd FILL
XFILL_1__13582_ vdd gnd FILL
X_13438_ _13438_/D _13438_/CLK _13438_/Q vdd gnd DFFPOSX1
XFILL_0__7830_ vdd gnd FILL
XFILL_1__10794_ vdd gnd FILL
XFILL_2__8746_ vdd gnd FILL
XFILL_1__12533_ vdd gnd FILL
XFILL_0__11174_ vdd gnd FILL
XFILL_0__7761_ vdd gnd FILL
X_13369_ _13369_/A _13369_/B _13369_/C _13369_/Y vdd gnd OAI21X1
XFILL_2__13823_ vdd gnd FILL
XFILL_0__10125_ vdd gnd FILL
XFILL_2__8677_ vdd gnd FILL
XFILL_0__9500_ vdd gnd FILL
XFILL_1__12464_ vdd gnd FILL
XFILL_0__7692_ vdd gnd FILL
XFILL_1__11415_ vdd gnd FILL
XFILL_2__13754_ vdd gnd FILL
XFILL_0__10056_ vdd gnd FILL
XFILL_0__9431_ vdd gnd FILL
XFILL_1__12395_ vdd gnd FILL
XFILL_2__12705_ vdd gnd FILL
XFILL_1__14134_ vdd gnd FILL
XFILL_1__11346_ vdd gnd FILL
XFILL_0__14864_ vdd gnd FILL
XFILL_0__9362_ vdd gnd FILL
X_9990_ _9990_/A _9990_/B _9990_/C _9990_/Y vdd gnd OAI21X1
XFILL_2__12636_ vdd gnd FILL
XFILL_1__14065_ vdd gnd FILL
XFILL_0__13815_ vdd gnd FILL
XFILL_0__8313_ vdd gnd FILL
XFILL_1__11277_ vdd gnd FILL
XFILL_0__14795_ vdd gnd FILL
XFILL_0__9293_ vdd gnd FILL
XFILL_2__9229_ vdd gnd FILL
X_8941_ _8941_/A _8941_/B _8941_/C _8941_/Y vdd gnd OAI21X1
XFILL_1__13016_ vdd gnd FILL
XFILL_1__10228_ vdd gnd FILL
XFILL_0__13746_ vdd gnd FILL
XFILL_0__10958_ vdd gnd FILL
XFILL_0__8244_ vdd gnd FILL
XFILL_2__14306_ vdd gnd FILL
X_8872_ _8872_/D _8872_/CLK _8872_/Q vdd gnd DFFPOSX1
XFILL_2__11518_ vdd gnd FILL
XFILL_1__10159_ vdd gnd FILL
XFILL_0__13677_ vdd gnd FILL
X_7823_ _7823_/A _7823_/B _7823_/Y vdd gnd NAND2X1
XFILL_0__8175_ vdd gnd FILL
XFILL_0__10889_ vdd gnd FILL
XFILL_2__14237_ vdd gnd FILL
XFILL_2__11449_ vdd gnd FILL
XFILL_0__12628_ vdd gnd FILL
XFILL_0__7126_ vdd gnd FILL
X_7754_ _7754_/A _7754_/B _7754_/Y vdd gnd OR2X2
XFILL_1__13918_ vdd gnd FILL
XFILL_2__13119_ vdd gnd FILL
X_7685_ _7685_/A _7685_/B _7685_/C _7685_/Y vdd gnd OAI21X1
XFILL_1__13849_ vdd gnd FILL
XFILL_2__14099_ vdd gnd FILL
X_9424_ _9424_/A _9424_/B _9424_/C _9424_/Y vdd gnd OAI21X1
XFILL_1__7870_ vdd gnd FILL
XFILL_0__14229_ vdd gnd FILL
X_9355_ _9355_/A _9355_/B _9355_/C _9355_/Y vdd gnd OAI21X1
XFILL_1__9540_ vdd gnd FILL
X_8306_ _8306_/A _8306_/B _8306_/C _8306_/Y vdd gnd NAND3X1
X_9286_ _9286_/A _9286_/B _9286_/Y vdd gnd NAND2X1
XFILL_1__9471_ vdd gnd FILL
X_8237_ _8237_/A _8237_/B _8237_/Y vdd gnd NAND2X1
XFILL_1__8422_ vdd gnd FILL
XFILL_0__9629_ vdd gnd FILL
X_8168_ _8168_/A _8168_/B _8168_/C _8168_/D _8168_/Y vdd gnd AOI22X1
X_7119_ _7119_/A _7119_/B _7119_/C _7119_/Y vdd gnd OAI21X1
XFILL_1__8353_ vdd gnd FILL
X_8099_ _8099_/A _8099_/Y vdd gnd INVX1
XFILL_1__7304_ vdd gnd FILL
XFILL_1__8284_ vdd gnd FILL
XFILL_1__7235_ vdd gnd FILL
XFILL_1_BUFX2_insert305 vdd gnd FILL
X_12740_ _12740_/A _12740_/B _12740_/C _12740_/Y vdd gnd OAI21X1
XFILL_1_BUFX2_insert316 vdd gnd FILL
XFILL_1__7166_ vdd gnd FILL
XFILL_1_BUFX2_insert327 vdd gnd FILL
XFILL_1_BUFX2_insert338 vdd gnd FILL
XFILL_1_BUFX2_insert349 vdd gnd FILL
X_12671_ _12671_/A _12671_/Y vdd gnd INVX1
XFILL_1__7097_ vdd gnd FILL
X_14410_ _14410_/A _14410_/B _14410_/C _14410_/D _14410_/Y vdd gnd AOI22X1
X_11622_ _11622_/D _11622_/CLK _11622_/Q vdd gnd DFFPOSX1
X_14341_ _14341_/A _14341_/B _14341_/Y vdd gnd NAND2X1
X_11553_ _11553_/A _11553_/B _11553_/C _11553_/Y vdd gnd OAI21X1
X_10504_ _10504_/A _10504_/B _10504_/Y vdd gnd NOR2X1
X_14272_ _14272_/A _14272_/B _14272_/Y vdd gnd NAND2X1
X_11484_ _11484_/A _11484_/Y vdd gnd INVX1
XFILL_1__7999_ vdd gnd FILL
X_13223_ _13223_/A _13223_/B _13223_/C _13223_/Y vdd gnd OAI21X1
X_10435_ _10435_/A _10435_/B _10435_/C _10435_/Y vdd gnd OAI21X1
XFILL_1__9738_ vdd gnd FILL
X_13154_ _13154_/A _13154_/B _13154_/C _13154_/Y vdd gnd AOI21X1
X_10366_ _10366_/A _10366_/B _10366_/C _10366_/Y vdd gnd OAI21X1
XFILL257250x79350 vdd gnd FILL
XFILL_2__8462_ vdd gnd FILL
XFILL_1__9669_ vdd gnd FILL
X_12105_ _12105_/A _12105_/B _12105_/Y vdd gnd NAND2X1
X_13085_ _13085_/A _13085_/B _13085_/Y vdd gnd NAND2X1
X_10297_ _10297_/A _10297_/B _10297_/Y vdd gnd OR2X2
XFILL_1__11200_ vdd gnd FILL
XFILL_2__8393_ vdd gnd FILL
XFILL_0__11930_ vdd gnd FILL
XFILL_1__12180_ vdd gnd FILL
X_12036_ _12036_/A _12036_/B _12036_/Y vdd gnd OR2X2
XFILL_1__11131_ vdd gnd FILL
XFILL_2__10682_ vdd gnd FILL
XFILL_0__11861_ vdd gnd FILL
XFILL_1__11062_ vdd gnd FILL
XFILL_0__13600_ vdd gnd FILL
XFILL_0__10812_ vdd gnd FILL
XFILL_0__14580_ vdd gnd FILL
XFILL_2__9014_ vdd gnd FILL
XFILL_0__11792_ vdd gnd FILL
X_13987_ _13987_/A _13987_/B _13987_/C _13987_/Y vdd gnd NAND3X1
XFILL_1__10013_ vdd gnd FILL
XFILL_0__13531_ vdd gnd FILL
XFILL_2_BUFX2_insert172 vdd gnd FILL
X_12938_ _12938_/A _12938_/B _12938_/C _12938_/Y vdd gnd OAI21X1
XFILL_2__11303_ vdd gnd FILL
XFILL_2_BUFX2_insert194 vdd gnd FILL
XFILL_1__14821_ vdd gnd FILL
XFILL_0__10674_ vdd gnd FILL
X_12869_ _12869_/A _12869_/Y vdd gnd INVX1
XFILL_2__11234_ vdd gnd FILL
XFILL_1__14752_ vdd gnd FILL
XFILL_0__12413_ vdd gnd FILL
XFILL_1__11964_ vdd gnd FILL
X_14608_ _14608_/A _14608_/Y vdd gnd INVX1
XFILL_0__13393_ vdd gnd FILL
XFILL_2__9916_ vdd gnd FILL
XFILL_0__9980_ vdd gnd FILL
XFILL_1__13703_ vdd gnd FILL
XFILL_2__11165_ vdd gnd FILL
XFILL_1__10915_ vdd gnd FILL
XFILL_1__14683_ vdd gnd FILL
XFILL_0__12344_ vdd gnd FILL
XFILL_1__11895_ vdd gnd FILL
XFILL_0__8931_ vdd gnd FILL
X_14539_ _14539_/D _14539_/CLK _14539_/Q vdd gnd DFFPOSX1
X_7470_ _7470_/A _7470_/B _7470_/Y vdd gnd NAND2X1
XBUFX2_insert160 BUFX2_insert160/A BUFX2_insert160/Y vdd gnd BUFX2
XFILL_1__13634_ vdd gnd FILL
XFILL_2__9847_ vdd gnd FILL
XFILL_0__12275_ vdd gnd FILL
XBUFX2_insert171 BUFX2_insert171/A BUFX2_insert171/Y vdd gnd BUFX2
XFILL_1__10846_ vdd gnd FILL
XFILL_2__11096_ vdd gnd FILL
XBUFX2_insert182 BUFX2_insert182/A BUFX2_insert182/Y vdd gnd BUFX2
XBUFX2_insert193 BUFX2_insert193/A BUFX2_insert193/Y vdd gnd BUFX2
XFILL_0__14014_ vdd gnd FILL
XFILL_1__13565_ vdd gnd FILL
XFILL_0__11226_ vdd gnd FILL
XFILL_0__7813_ vdd gnd FILL
XFILL_1__10777_ vdd gnd FILL
X_9140_ _9140_/A _9140_/B _9140_/C _9140_/Y vdd gnd AOI21X1
XFILL_0__8793_ vdd gnd FILL
XFILL_2__8729_ vdd gnd FILL
XFILL_1__12516_ vdd gnd FILL
XFILL_2__14855_ vdd gnd FILL
XFILL_0__11157_ vdd gnd FILL
XFILL_0__7744_ vdd gnd FILL
X_9071_ _9071_/A _9071_/B _9071_/Y vdd gnd OR2X2
XFILL_0__10108_ vdd gnd FILL
XFILL_2__13806_ vdd gnd FILL
XFILL_1__12447_ vdd gnd FILL
XFILL_0__11088_ vdd gnd FILL
XFILL_2__14786_ vdd gnd FILL
XFILL_2__11998_ vdd gnd FILL
X_8022_ _8022_/A _8022_/B _8022_/C _8022_/Y vdd gnd AOI21X1
XFILL_0__7675_ vdd gnd FILL
XFILL_0__10039_ vdd gnd FILL
XFILL_0__14916_ vdd gnd FILL
XFILL_2__13737_ vdd gnd FILL
XFILL_0__9414_ vdd gnd FILL
XFILL_1__12378_ vdd gnd FILL
XFILL_1__14117_ vdd gnd FILL
XFILL_2__13668_ vdd gnd FILL
XFILL_1__11329_ vdd gnd FILL
XFILL_0__14847_ vdd gnd FILL
XFILL_0__9345_ vdd gnd FILL
XFILL_2__12619_ vdd gnd FILL
X_9973_ _9973_/A _9973_/B _9973_/Y vdd gnd OR2X2
XFILL_1__14048_ vdd gnd FILL
XFILL_2__13599_ vdd gnd FILL
XFILL_0__14778_ vdd gnd FILL
XFILL_0__9276_ vdd gnd FILL
X_8924_ _8924_/A _8924_/B _8924_/Y vdd gnd NOR2X1
XFILL_0__13729_ vdd gnd FILL
XFILL_0__8227_ vdd gnd FILL
X_8855_ _8855_/D _8855_/CLK _8855_/Q vdd gnd DFFPOSX1
X_7806_ _7806_/A _7806_/B _7806_/Y vdd gnd NOR2X1
XFILL_0__8158_ vdd gnd FILL
X_8786_ _8786_/A _8786_/B _8786_/Y vdd gnd NAND2X1
XFILL_0__7109_ vdd gnd FILL
X_7737_ _7737_/A _7737_/Y vdd gnd INVX1
XFILL_0__8089_ vdd gnd FILL
XFILL_1__8971_ vdd gnd FILL
X_7668_ _7668_/A _7668_/B _7668_/Y vdd gnd NOR2X1
X_9407_ _9407_/A _9407_/B _9407_/C _9407_/Y vdd gnd NAND3X1
XFILL_1__7853_ vdd gnd FILL
X_7599_ _7599_/A _7599_/Y vdd gnd INVX1
X_9338_ _9338_/A _9338_/B _9338_/Y vdd gnd NAND2X1
XFILL_1__7784_ vdd gnd FILL
X_10220_ _10220_/A _10220_/B _10220_/Y vdd gnd NAND2X1
XFILL_1__9523_ vdd gnd FILL
X_9269_ _9269_/A _9269_/Y vdd gnd INVX1
X_10151_ _10151_/A _10151_/B _10151_/C _10151_/Y vdd gnd NOR3X1
XFILL_1__9454_ vdd gnd FILL
X_10082_ _10082_/A _10082_/B _10082_/C _10082_/Y vdd gnd NAND3X1
XFILL_1__8405_ vdd gnd FILL
XFILL_1__9385_ vdd gnd FILL
X_13910_ _13910_/A _13910_/Y vdd gnd INVX1
XFILL_1__8336_ vdd gnd FILL
X_14890_ _14890_/D _14890_/CLK _14890_/Q vdd gnd DFFPOSX1
X_13841_ _13841_/A _13841_/B _13841_/Y vdd gnd NAND2X1
XFILL_1__8267_ vdd gnd FILL
XFILL257550x183750 vdd gnd FILL
XFILL_1__7218_ vdd gnd FILL
X_13772_ _13772_/A _13772_/B _13772_/C _13772_/Y vdd gnd NAND3X1
X_10984_ _10984_/A _10984_/B _10984_/C _10984_/Y vdd gnd NOR3X1
XFILL_1__8198_ vdd gnd FILL
XFILL_1_BUFX2_insert113 vdd gnd FILL
XFILL_1_BUFX2_insert124 vdd gnd FILL
XFILL_1_BUFX2_insert135 vdd gnd FILL
XFILL257250x54150 vdd gnd FILL
X_12723_ _12723_/A _12723_/B _12723_/S _12723_/Y vdd gnd MUX2X1
XFILL_1__7149_ vdd gnd FILL
XFILL_1_BUFX2_insert146 vdd gnd FILL
XFILL_1_BUFX2_insert157 vdd gnd FILL
XFILL_1_BUFX2_insert168 vdd gnd FILL
X_12654_ _12654_/A _12654_/Y vdd gnd INVX1
XFILL_1_BUFX2_insert179 vdd gnd FILL
XFILL_0__10390_ vdd gnd FILL
X_11605_ _11605_/A _11605_/B _11605_/C _11605_/Y vdd gnd OAI21X1
XFILL_2__9701_ vdd gnd FILL
X_12585_ _12585_/D _12585_/CLK _12585_/Q vdd gnd DFFPOSX1
X_14324_ _14324_/A _14324_/Y vdd gnd INVX1
X_11536_ _11536_/A _11536_/B _11536_/Y vdd gnd OR2X2
XFILL_1__10631_ vdd gnd FILL
XFILL_0__12060_ vdd gnd FILL
X_14255_ _14255_/A _14255_/B _14255_/C _14255_/Y vdd gnd OAI21X1
X_11467_ _11467_/A _11467_/B _11467_/C _11467_/Y vdd gnd OAI21X1
XFILL_0__11011_ vdd gnd FILL
XFILL_1__13350_ vdd gnd FILL
X_13206_ _13206_/A _13206_/B _13206_/C _13206_/Y vdd gnd OAI21X1
XFILL_1__10562_ vdd gnd FILL
X_10418_ _10418_/A _10418_/B _10418_/Y vdd gnd OR2X2
X_14186_ _14186_/D _14186_/CLK _14186_/Q vdd gnd DFFPOSX1
XFILL_1__12301_ vdd gnd FILL
X_11398_ _11398_/A _11398_/B _11398_/C _11398_/Y vdd gnd OAI21X1
XFILL_1__13281_ vdd gnd FILL
X_13137_ _13137_/A _13137_/Y vdd gnd INVX1
XFILL_1__10493_ vdd gnd FILL
X_10349_ _10349_/A _10349_/B _10349_/C _10349_/Y vdd gnd NAND3X1
XFILL_2__10803_ vdd gnd FILL
XFILL_1__12232_ vdd gnd FILL
XFILL_0__12962_ vdd gnd FILL
XFILL_0__7460_ vdd gnd FILL
X_13068_ _13068_/A _13068_/B _13068_/C _13068_/Y vdd gnd OAI21X1
XFILL_2__13522_ vdd gnd FILL
XFILL_0__14701_ vdd gnd FILL
XFILL_0__11913_ vdd gnd FILL
XFILL_1__12163_ vdd gnd FILL
X_12019_ _12019_/A _12019_/B _12019_/Y vdd gnd NAND2X1
XFILL_0__12893_ vdd gnd FILL
XFILL_0__7391_ vdd gnd FILL
XFILL_2__7327_ vdd gnd FILL
XFILL_1__11114_ vdd gnd FILL
XFILL_0__14632_ vdd gnd FILL
XFILL_0__9130_ vdd gnd FILL
XFILL_0__11844_ vdd gnd FILL
XFILL_1__12094_ vdd gnd FILL
XFILL_2__7258_ vdd gnd FILL
XFILL_1__11045_ vdd gnd FILL
XFILL_2__13384_ vdd gnd FILL
XFILL_0__14563_ vdd gnd FILL
XFILL_2__10596_ vdd gnd FILL
XFILL_0__9061_ vdd gnd FILL
XFILL_0__11775_ vdd gnd FILL
XFILL_0__13514_ vdd gnd FILL
XFILL_0__8012_ vdd gnd FILL
XFILL_0__14494_ vdd gnd FILL
X_8640_ _8640_/A _8640_/Y vdd gnd INVX1
XFILL_1__14804_ vdd gnd FILL
XFILL_0__10657_ vdd gnd FILL
XFILL_1__12996_ vdd gnd FILL
X_8571_ _8571_/A _8571_/B _8571_/C _8571_/Y vdd gnd NAND3X1
XFILL_2__11217_ vdd gnd FILL
XFILL_1__14735_ vdd gnd FILL
XFILL_1__11947_ vdd gnd FILL
XFILL_0__13376_ vdd gnd FILL
X_7522_ _7522_/A _7522_/Y vdd gnd INVX1
XFILL_0__10588_ vdd gnd FILL
XFILL_0__9963_ vdd gnd FILL
XFILL_2__11148_ vdd gnd FILL
XFILL_1__14666_ vdd gnd FILL
XFILL_0__12327_ vdd gnd FILL
XFILL_1__11878_ vdd gnd FILL
X_7453_ _7453_/A _7453_/B _7453_/Y vdd gnd NAND2X1
XFILL_0__9894_ vdd gnd FILL
XFILL_1__13617_ vdd gnd FILL
XFILL_1__10829_ vdd gnd FILL
XFILL_2__11079_ vdd gnd FILL
XFILL_1__14597_ vdd gnd FILL
XFILL_0__12258_ vdd gnd FILL
X_7384_ _7384_/A _7384_/B _7384_/C _7384_/Y vdd gnd OAI21X1
XFILL_0__11209_ vdd gnd FILL
XFILL_1__13548_ vdd gnd FILL
X_9123_ _9123_/A _9123_/B _9123_/Y vdd gnd NAND2X1
XFILL_0__12189_ vdd gnd FILL
XFILL_0__8776_ vdd gnd FILL
XFILL_0__7727_ vdd gnd FILL
X_9054_ _9054_/A _9054_/B _9054_/C _9054_/Y vdd gnd OAI21X1
X_8005_ _8005_/A _8005_/B _8005_/Y vdd gnd AND2X2
XFILL_0__7658_ vdd gnd FILL
XFILL_1__9170_ vdd gnd FILL
XFILL_0__7589_ vdd gnd FILL
XFILL_1__8121_ vdd gnd FILL
XFILL_0__9328_ vdd gnd FILL
X_9956_ _9956_/A _9956_/B _9956_/C _9956_/Y vdd gnd OAI21X1
XFILL_0__9259_ vdd gnd FILL
XFILL_1__8052_ vdd gnd FILL
X_8907_ _8907_/D _8907_/CLK _8907_/Q vdd gnd DFFPOSX1
X_9887_ _9887_/A _9887_/B _9887_/C _9887_/Y vdd gnd OAI21X1
X_8838_ _8838_/A _8838_/B _8838_/Y vdd gnd NAND2X1
XFILL257550x115350 vdd gnd FILL
XFILL_0_BUFX2_insert109 vdd gnd FILL
X_8769_ _8769_/A _8769_/B _8769_/C _8769_/Y vdd gnd OAI21X1
XFILL_1__8954_ vdd gnd FILL
X_12370_ _12370_/A _12370_/B _12370_/C _12370_/Y vdd gnd OAI21X1
XFILL_1__7905_ vdd gnd FILL
X_11321_ _11321_/A _11321_/B _11321_/C _11321_/Y vdd gnd OAI21X1
XFILL_1__7836_ vdd gnd FILL
X_14040_ _14040_/A _14040_/Y vdd gnd INVX1
X_11252_ _11252_/A _11252_/B _11252_/Y vdd gnd NAND2X1
XFILL_1_CLKBUF1_insert389 vdd gnd FILL
XFILL_1__7767_ vdd gnd FILL
X_10203_ _10203_/A _10203_/B _10203_/C _10203_/Y vdd gnd OAI21X1
XFILL_1__9506_ vdd gnd FILL
X_11183_ _11183_/A _11183_/B _11183_/Y vdd gnd NAND2X1
XFILL_1__7698_ vdd gnd FILL
X_10134_ _10134_/A _10134_/B _10134_/C _10134_/Y vdd gnd NAND3X1
XFILL_1__9437_ vdd gnd FILL
X_10065_ _10065_/A _10065_/Y vdd gnd INVX1
XFILL_1__9368_ vdd gnd FILL
XFILL_2__7112_ vdd gnd FILL
X_14873_ _14873_/D _14873_/CLK _14873_/Q vdd gnd DFFPOSX1
XFILL_1__8319_ vdd gnd FILL
XFILL_1__9299_ vdd gnd FILL
X_13824_ _13824_/A _13824_/B _13824_/C _13824_/Y vdd gnd NAND3X1
XFILL_0__11560_ vdd gnd FILL
X_10967_ _10967_/A _10967_/B _10967_/C _10967_/Y vdd gnd NAND3X1
XFILL_2__12120_ vdd gnd FILL
X_13755_ _13755_/A _13755_/B _13755_/C _13755_/Y vdd gnd NAND3X1
XFILL_0__10511_ vdd gnd FILL
XFILL_1__12850_ vdd gnd FILL
XFILL_0__11491_ vdd gnd FILL
X_12706_ _12706_/A _12706_/B _12706_/C _12706_/D _12706_/Y vdd gnd OAI22X1
XFILL_2__12051_ vdd gnd FILL
XFILL_1__11801_ vdd gnd FILL
X_10898_ _10898_/A _10898_/B _10898_/C _10898_/Y vdd gnd AOI21X1
X_13686_ _13686_/A _13686_/B _13686_/Y vdd gnd NOR2X1
XFILL_0__13230_ vdd gnd FILL
XFILL_0__10442_ vdd gnd FILL
XFILL_1__12781_ vdd gnd FILL
X_12637_ _12637_/A _12637_/B _12637_/Y vdd gnd NAND2X1
XFILL_1__11732_ vdd gnd FILL
XFILL_0__13161_ vdd gnd FILL
XFILL_0__10373_ vdd gnd FILL
X_12568_ _12568_/D _12568_/CLK _12568_/Q vdd gnd DFFPOSX1
XFILL_0__12112_ vdd gnd FILL
XFILL_1__14451_ vdd gnd FILL
X_14307_ _14307_/A _14307_/B _14307_/C _14307_/Y vdd gnd NAND3X1
X_11519_ _11519_/A _11519_/B _11519_/Y vdd gnd NAND2X1
XFILL_0__13092_ vdd gnd FILL
XFILL_2__9615_ vdd gnd FILL
X_12499_ _12499_/A _12499_/B _12499_/C _12499_/Y vdd gnd OAI21X1
XFILL_1__13402_ vdd gnd FILL
XFILL_1__10614_ vdd gnd FILL
XFILL_2__12953_ vdd gnd FILL
XFILL_1__14382_ vdd gnd FILL
XFILL_0__12043_ vdd gnd FILL
XFILL_0__8630_ vdd gnd FILL
XFILL_1__11594_ vdd gnd FILL
X_14238_ _14238_/A _14238_/B _14238_/Y vdd gnd NAND2X1
XFILL_2__9546_ vdd gnd FILL
XFILL_1__13333_ vdd gnd FILL
XFILL_2__12884_ vdd gnd FILL
XFILL_1__10545_ vdd gnd FILL
XFILL_0__8561_ vdd gnd FILL
X_14169_ _14169_/D _14169_/CLK _14169_/Q vdd gnd DFFPOSX1
XFILL_2__9477_ vdd gnd FILL
XFILL_1__13264_ vdd gnd FILL
XFILL_0__7512_ vdd gnd FILL
XFILL_1__10476_ vdd gnd FILL
XFILL_0__13994_ vdd gnd FILL
XFILL_0__8492_ vdd gnd FILL
XFILL_1__12215_ vdd gnd FILL
XFILL_1__13195_ vdd gnd FILL
XFILL_0__12945_ vdd gnd FILL
XCLKBUF1_insert388 CLKBUF1_insert388/A CLKBUF1_insert388/Y vdd gnd CLKBUF1
XFILL_0__7443_ vdd gnd FILL
XFILL_2__14485_ vdd gnd FILL
XFILL_1__12146_ vdd gnd FILL
X_9810_ _9810_/D _9810_/CLK _9810_/Q vdd gnd DFFPOSX1
XFILL_0__12876_ vdd gnd FILL
XFILL_0__7374_ vdd gnd FILL
XFILL_0__14615_ vdd gnd FILL
XFILL_0__9113_ vdd gnd FILL
XFILL_0__11827_ vdd gnd FILL
XFILL_1__12077_ vdd gnd FILL
X_9741_ _9741_/A _9741_/B _9741_/C _9741_/Y vdd gnd OAI21X1
XFILL_1__11028_ vdd gnd FILL
XFILL_2__13367_ vdd gnd FILL
XFILL_0__9044_ vdd gnd FILL
XFILL_0__11758_ vdd gnd FILL
X_9672_ _9672_/A _9672_/B _9672_/Y vdd gnd NAND2X1
XFILL_2__13298_ vdd gnd FILL
XFILL_0__14477_ vdd gnd FILL
X_8623_ _8623_/A _8623_/B _8623_/Y vdd gnd AND2X2
XFILL_1__12979_ vdd gnd FILL
X_8554_ _8554_/A _8554_/B _8554_/C _8554_/Y vdd gnd AOI21X1
XFILL_1__14718_ vdd gnd FILL
XFILL_0__13359_ vdd gnd FILL
X_7505_ _7505_/A _7505_/B _7505_/Y vdd gnd NOR2X1
XFILL_0__9946_ vdd gnd FILL
X_8485_ _8485_/A _8485_/B _8485_/C _8485_/Y vdd gnd NAND3X1
XFILL_1__14649_ vdd gnd FILL
X_7436_ _7436_/A _7436_/B _7436_/Y vdd gnd NAND2X1
XFILL_1__8670_ vdd gnd FILL
XFILL_0__9877_ vdd gnd FILL
XFILL_1__7621_ vdd gnd FILL
XFILL_0__8828_ vdd gnd FILL
X_7367_ _7367_/A _7367_/Y vdd gnd INVX1
X_9106_ _9106_/A _9106_/Y vdd gnd INVX1
XFILL_1__7552_ vdd gnd FILL
XFILL_0__8759_ vdd gnd FILL
X_7298_ _7298_/A _7298_/B _7298_/C _7298_/Y vdd gnd OAI21X1
X_9037_ _9037_/A _9037_/B _9037_/S _9037_/Y vdd gnd MUX2X1
XFILL_1__7483_ vdd gnd FILL
XFILL_1__9222_ vdd gnd FILL
XFILL_1__9153_ vdd gnd FILL
XFILL_1__8104_ vdd gnd FILL
X_11870_ _11870_/A _11870_/B _11870_/C _11870_/Y vdd gnd NAND3X1
XFILL_1__9084_ vdd gnd FILL
X_9939_ _9939_/A _9939_/B _9939_/C _9939_/Y vdd gnd NAND3X1
X_10821_ _10821_/A _10821_/B _10821_/C _10821_/Y vdd gnd OAI21X1
XFILL_1__8035_ vdd gnd FILL
X_10752_ _10752_/D _10752_/CLK _10752_/Q vdd gnd DFFPOSX1
X_13540_ _13540_/A _13540_/B _13540_/C _13540_/D _13540_/Y vdd gnd AOI22X1
X_13471_ _13471_/D _13471_/CLK _13471_/Q vdd gnd DFFPOSX1
X_10683_ _10683_/A _10683_/B _10683_/C _10683_/Y vdd gnd OAI21X1
XFILL_1__9986_ vdd gnd FILL
X_12422_ _12422_/A _12422_/B _12422_/Y vdd gnd NOR2X1
XFILL_1__8937_ vdd gnd FILL
X_12353_ _12353_/A _12353_/B _12353_/C _12353_/Y vdd gnd OAI21X1
X_11304_ _11304_/A _11304_/B _11304_/Y vdd gnd NAND2X1
XFILL_2__9400_ vdd gnd FILL
X_12284_ _12284_/A _12284_/B _12284_/Y vdd gnd NAND2X1
XFILL_1__7819_ vdd gnd FILL
XFILL_1__8799_ vdd gnd FILL
X_14023_ _14023_/A _14023_/B _14023_/C _14023_/Y vdd gnd NAND3X1
X_11235_ _11235_/A _11235_/B _11235_/Y vdd gnd OR2X2
XFILL_2__9331_ vdd gnd FILL
XFILL_1__10330_ vdd gnd FILL
X_11166_ _11166_/A _11166_/B _11166_/Y vdd gnd NAND2X1
XFILL_2__9262_ vdd gnd FILL
XFILL_1__10261_ vdd gnd FILL
X_10117_ _10117_/A _10117_/B _10117_/C _10117_/Y vdd gnd OAI21X1
XFILL_0__10991_ vdd gnd FILL
XFILL_1__12000_ vdd gnd FILL
X_11097_ _11097_/A _11097_/B _11097_/C _11097_/Y vdd gnd OAI21X1
XFILL_2__9193_ vdd gnd FILL
XFILL_2__11551_ vdd gnd FILL
XFILL_0__12730_ vdd gnd FILL
XFILL_1__10192_ vdd gnd FILL
X_10048_ _10048_/A _10048_/B _10048_/C _10048_/Y vdd gnd AOI21X1
XFILL_2__14270_ vdd gnd FILL
XFILL_2__11482_ vdd gnd FILL
XFILL_0__12661_ vdd gnd FILL
X_14856_ _14856_/A _14856_/B _14856_/C _14856_/Y vdd gnd OAI21X1
XFILL_0__14400_ vdd gnd FILL
XFILL_1__13951_ vdd gnd FILL
X_13807_ _13807_/A _13807_/B _13807_/C _13807_/Y vdd gnd OAI21X1
XFILL_0__7090_ vdd gnd FILL
XFILL_1__12902_ vdd gnd FILL
X_14787_ _14787_/A _14787_/B _14787_/Y vdd gnd AND2X2
X_11999_ _11999_/A _11999_/B _11999_/C _11999_/Y vdd gnd NOR3X1
XFILL_0__14331_ vdd gnd FILL
XFILL_0__11543_ vdd gnd FILL
XFILL_1__13882_ vdd gnd FILL
XFILL_2__12103_ vdd gnd FILL
X_13738_ _13738_/A _13738_/B _13738_/C _13738_/Y vdd gnd NAND3X1
XFILL_1__12833_ vdd gnd FILL
XFILL_0__14262_ vdd gnd FILL
XFILL_0__11474_ vdd gnd FILL
X_13669_ _13669_/A _13669_/B _13669_/C _13669_/Y vdd gnd OAI21X1
XFILL_2__12034_ vdd gnd FILL
XFILL_0__13213_ vdd gnd FILL
XFILL_0__10425_ vdd gnd FILL
XFILL_1__12764_ vdd gnd FILL
XFILL_1__11715_ vdd gnd FILL
XFILL_0__13144_ vdd gnd FILL
XFILL_0__10356_ vdd gnd FILL
XFILL_1__12695_ vdd gnd FILL
XFILL_0__9731_ vdd gnd FILL
X_8270_ _8270_/A _8270_/B _8270_/C _8270_/Y vdd gnd OAI21X1
XFILL_1__14434_ vdd gnd FILL
XFILL_0__13075_ vdd gnd FILL
XFILL_0__10287_ vdd gnd FILL
XFILL_2__13985_ vdd gnd FILL
X_7221_ _7221_/A _7221_/B _7221_/C _7221_/Y vdd gnd NAND3X1
XFILL_0__9662_ vdd gnd FILL
XFILL_2__12936_ vdd gnd FILL
XFILL_0__12026_ vdd gnd FILL
XFILL_1__14365_ vdd gnd FILL
XFILL_1__11577_ vdd gnd FILL
XFILL_0__8613_ vdd gnd FILL
X_7152_ _7152_/A _7152_/B _7152_/Y vdd gnd NAND2X1
XFILL_2__9529_ vdd gnd FILL
XFILL_0__9593_ vdd gnd FILL
XFILL_1__13316_ vdd gnd FILL
XFILL_1__10528_ vdd gnd FILL
XFILL_1__14296_ vdd gnd FILL
XFILL_2__12867_ vdd gnd FILL
XFILL_0__8544_ vdd gnd FILL
X_7083_ _7083_/A _7083_/B _7083_/C _7083_/Y vdd gnd OAI21X1
XFILL_1__13247_ vdd gnd FILL
XFILL_1__10459_ vdd gnd FILL
XFILL_2__12798_ vdd gnd FILL
XFILL_0__13977_ vdd gnd FILL
XFILL_0__8475_ vdd gnd FILL
XFILL_1__13178_ vdd gnd FILL
XFILL_0__12928_ vdd gnd FILL
XFILL_0__7426_ vdd gnd FILL
XFILL_1__12129_ vdd gnd FILL
XFILL_2__14468_ vdd gnd FILL
XFILL_0__12859_ vdd gnd FILL
XFILL_0__7357_ vdd gnd FILL
X_7985_ _7985_/D _7985_/CLK _7985_/Q vdd gnd DFFPOSX1
XFILL_2__14399_ vdd gnd FILL
X_9724_ _9724_/A _9724_/B _9724_/Y vdd gnd NAND2X1
XFILL_0__7288_ vdd gnd FILL
XFILL_0__9027_ vdd gnd FILL
X_9655_ _9655_/A _9655_/B _9655_/Y vdd gnd NAND2X1
X_8606_ _8606_/A _8606_/B _8606_/Y vdd gnd AND2X2
X_9586_ _9586_/A _9586_/B _9586_/C _9586_/Y vdd gnd AOI21X1
X_8537_ _8537_/A _8537_/B _8537_/Y vdd gnd NAND2X1
XFILL_0__9929_ vdd gnd FILL
XFILL_1__8722_ vdd gnd FILL
X_8468_ _8468_/A _8468_/B _8468_/C _8468_/Y vdd gnd OAI21X1
X_7419_ _7419_/A _7419_/Y vdd gnd INVX1
XFILL_1__8653_ vdd gnd FILL
X_8399_ _8399_/A _8399_/B _8399_/S _8399_/Y vdd gnd MUX2X1
XFILL_1__7604_ vdd gnd FILL
XFILL_1__8584_ vdd gnd FILL
X_11020_ _11020_/A _11020_/B _11020_/C _11020_/Y vdd gnd NAND3X1
XFILL_1__7535_ vdd gnd FILL
XFILL_1__7466_ vdd gnd FILL
XFILL_1__9205_ vdd gnd FILL
X_12971_ _12971_/A _12971_/B _12971_/Y vdd gnd NAND2X1
XFILL_1__7397_ vdd gnd FILL
X_14710_ _14710_/A _14710_/B _14710_/C _14710_/Y vdd gnd AOI21X1
X_11922_ _11922_/A _11922_/B _11922_/C _11922_/Y vdd gnd AOI21X1
XFILL_1__9136_ vdd gnd FILL
X_14641_ _14641_/A _14641_/B _14641_/C _14641_/Y vdd gnd OAI21X1
XFILL_1__9067_ vdd gnd FILL
X_11853_ _11853_/A _11853_/B _11853_/C _11853_/Y vdd gnd OAI21X1
X_10804_ _10804_/A _10804_/Y vdd gnd INVX1
X_14572_ _14572_/A _14572_/B _14572_/C _14572_/Y vdd gnd OAI21X1
XFILL_1__8018_ vdd gnd FILL
X_11784_ _11784_/A _11784_/B _11784_/Y vdd gnd NAND2X1
X_13523_ _13523_/A _13523_/B _13523_/Y vdd gnd NAND2X1
X_10735_ _10735_/D _10735_/CLK _10735_/Q vdd gnd DFFPOSX1
X_10666_ _10666_/A _10666_/Y vdd gnd INVX1
X_13454_ _13454_/D _13454_/CLK _13454_/Q vdd gnd DFFPOSX1
XFILL_0__10210_ vdd gnd FILL
XFILL_1__9969_ vdd gnd FILL
XFILL_0__11190_ vdd gnd FILL
X_12405_ _12405_/A _12405_/B _12405_/Y vdd gnd OR2X2
X_13385_ _13385_/A _13385_/B _13385_/C _13385_/Y vdd gnd OAI21X1
XFILL_2__7713_ vdd gnd FILL
X_10597_ _10597_/A _10597_/B _10597_/Y vdd gnd NAND2X1
XFILL_1__11500_ vdd gnd FILL
XFILL_0__10141_ vdd gnd FILL
XFILL_1__12480_ vdd gnd FILL
X_12336_ _12336_/A _12336_/Y vdd gnd INVX1
XFILL_2__7644_ vdd gnd FILL
XFILL_1__11431_ vdd gnd FILL
XFILL_2__10982_ vdd gnd FILL
XFILL_0__10072_ vdd gnd FILL
XFILL_2__13770_ vdd gnd FILL
X_12267_ _12267_/A _12267_/B _12267_/C _12267_/Y vdd gnd NAND3X1
XFILL_0__13900_ vdd gnd FILL
XFILL_1__14150_ vdd gnd FILL
XFILL_2__7575_ vdd gnd FILL
XFILL_1__11362_ vdd gnd FILL
X_14006_ _14006_/A _14006_/B _14006_/C _14006_/Y vdd gnd NAND3X1
X_11218_ _11218_/A _11218_/Y vdd gnd INVX1
XFILL_1__13101_ vdd gnd FILL
X_12198_ _12198_/A _12198_/B _12198_/C _12198_/Y vdd gnd NOR3X1
XFILL_2__12652_ vdd gnd FILL
XFILL_1__10313_ vdd gnd FILL
XFILL_0__13831_ vdd gnd FILL
XFILL_1__14081_ vdd gnd FILL
XFILL_1__11293_ vdd gnd FILL
X_11149_ _11149_/A _11149_/B _11149_/Y vdd gnd NAND2X1
XFILL_2__9245_ vdd gnd FILL
XFILL_1__13032_ vdd gnd FILL
XFILL_1__10244_ vdd gnd FILL
XFILL_0__13762_ vdd gnd FILL
XFILL_0__8260_ vdd gnd FILL
XFILL_0__10974_ vdd gnd FILL
XFILL_2__11534_ vdd gnd FILL
XFILL_2__9176_ vdd gnd FILL
XFILL_0__12713_ vdd gnd FILL
XFILL_1__10175_ vdd gnd FILL
XFILL_0__7211_ vdd gnd FILL
X_14908_ _14908_/A _14908_/Y vdd gnd BUFX2
XFILL_0__13693_ vdd gnd FILL
XFILL_0__8191_ vdd gnd FILL
XFILL_2__11465_ vdd gnd FILL
XFILL_0__12644_ vdd gnd FILL
XFILL_0__7142_ vdd gnd FILL
X_14839_ _14839_/A _14839_/B _14839_/Y vdd gnd NAND2X1
X_7770_ _7770_/A _7770_/B _7770_/Y vdd gnd NAND2X1
XFILL_1__13934_ vdd gnd FILL
XFILL_2__11396_ vdd gnd FILL
XFILL_0__7073_ vdd gnd FILL
XFILL_0__14314_ vdd gnd FILL
XFILL_0__11526_ vdd gnd FILL
XFILL_1__13865_ vdd gnd FILL
X_9440_ _9440_/A _9440_/B _9440_/C _9440_/Y vdd gnd NAND3X1
XFILL_0__14245_ vdd gnd FILL
XFILL_1__12816_ vdd gnd FILL
XFILL_0__11457_ vdd gnd FILL
XFILL_1__13796_ vdd gnd FILL
X_9371_ _9371_/A _9371_/B _9371_/C _9371_/Y vdd gnd NAND3X1
XFILL_2__12017_ vdd gnd FILL
XFILL_0__10408_ vdd gnd FILL
XFILL_1__12747_ vdd gnd FILL
XFILL_0_BUFX2_insert270 vdd gnd FILL
X_8322_ _8322_/A _8322_/B _8322_/C _8322_/Y vdd gnd NAND3X1
XFILL_0__11388_ vdd gnd FILL
XFILL_0_BUFX2_insert281 vdd gnd FILL
XFILL_0_BUFX2_insert292 vdd gnd FILL
XFILL_0__13127_ vdd gnd FILL
XFILL_0__10339_ vdd gnd FILL
XFILL_1__12678_ vdd gnd FILL
XFILL_0__9714_ vdd gnd FILL
X_8253_ _8253_/A _8253_/B _8253_/C _8253_/Y vdd gnd NAND3X1
XFILL_1__14417_ vdd gnd FILL
XFILL_2__13968_ vdd gnd FILL
XFILL_0__13058_ vdd gnd FILL
X_7204_ _7204_/A _7204_/Y vdd gnd INVX1
XFILL_0__9645_ vdd gnd FILL
X_8184_ _8184_/A _8184_/B _8184_/Y vdd gnd NAND2X1
XFILL_1__14348_ vdd gnd FILL
XFILL_0__12009_ vdd gnd FILL
XFILL_2__12919_ vdd gnd FILL
XFILL_2__13899_ vdd gnd FILL
X_7135_ _7135_/A _7135_/B _7135_/Y vdd gnd NAND2X1
XFILL_0__9576_ vdd gnd FILL
XFILL_1__14279_ vdd gnd FILL
XFILL_1__7320_ vdd gnd FILL
XFILL_0__8527_ vdd gnd FILL
XFILL_1__7251_ vdd gnd FILL
XFILL_0__8458_ vdd gnd FILL
XFILL_0__7409_ vdd gnd FILL
XFILL_1__7182_ vdd gnd FILL
XFILL_0__8389_ vdd gnd FILL
X_7968_ _7968_/D _7968_/CLK _7968_/Q vdd gnd DFFPOSX1
X_9707_ _9707_/A _9707_/B _9707_/C _9707_/Y vdd gnd OAI21X1
X_7899_ _7899_/A _7899_/B _7899_/C _7899_/Y vdd gnd OAI21X1
X_9638_ _9638_/A _9638_/B _9638_/Y vdd gnd NAND2X1
X_10520_ _10520_/A _10520_/B _10520_/C _10520_/Y vdd gnd OAI21X1
X_9569_ _9569_/A _9569_/B _9569_/Y vdd gnd NOR2X1
X_10451_ _10451_/A _10451_/B _10451_/Y vdd gnd NOR2X1
XFILL_1__9754_ vdd gnd FILL
X_13170_ _13170_/A _13170_/B _13170_/C _13170_/Y vdd gnd AOI21X1
X_10382_ _10382_/A _10382_/B _10382_/C _10382_/Y vdd gnd NAND3X1
XFILL_1__8705_ vdd gnd FILL
XFILL_1__9685_ vdd gnd FILL
X_12121_ _12121_/A _12121_/Y vdd gnd INVX1
XFILL_1__8636_ vdd gnd FILL
X_12052_ _12052_/A _12052_/B _12052_/C _12052_/Y vdd gnd OAI21X1
XFILL_2__7360_ vdd gnd FILL
XFILL_1__8567_ vdd gnd FILL
X_11003_ _11003_/A _11003_/B _11003_/C _11003_/Y vdd gnd OAI21X1
XFILL_1__7518_ vdd gnd FILL
XFILL_2__7291_ vdd gnd FILL
XFILL_0_CLKBUF1_insert36 vdd gnd FILL
XFILL_1__8498_ vdd gnd FILL
XFILL_0_CLKBUF1_insert47 vdd gnd FILL
XFILL_0_CLKBUF1_insert58 vdd gnd FILL
XFILL_2_BUFX2_insert310 vdd gnd FILL
XFILL_0_CLKBUF1_insert69 vdd gnd FILL
XFILL_1__7449_ vdd gnd FILL
XFILL_2_BUFX2_insert332 vdd gnd FILL
X_12954_ _12954_/A _12954_/B _12954_/C _12954_/D _12954_/Y vdd gnd AOI22X1
XFILL_2_BUFX2_insert365 vdd gnd FILL
X_11905_ _11905_/A _11905_/B _11905_/Y vdd gnd NAND2X1
XFILL_1__9119_ vdd gnd FILL
X_12885_ _12885_/A _12885_/Y vdd gnd INVX1
XFILL_1__11980_ vdd gnd FILL
X_14624_ _14624_/A _14624_/B _14624_/Y vdd gnd NAND2X1
XFILL_2__10201_ vdd gnd FILL
X_11836_ _11836_/A _11836_/B _11836_/Y vdd gnd NAND2X1
XFILL_1__10931_ vdd gnd FILL
XFILL_0__12360_ vdd gnd FILL
X_14555_ _14555_/D _14555_/CLK _14555_/Q vdd gnd DFFPOSX1
XFILL_2__10132_ vdd gnd FILL
X_11767_ _11767_/A _11767_/B _11767_/S _11767_/Y vdd gnd MUX2X1
XBUFX2_insert320 BUFX2_insert320/A BUFX2_insert320/Y vdd gnd BUFX2
XFILL_0__11311_ vdd gnd FILL
XFILL_1__13650_ vdd gnd FILL
XFILL_1__10862_ vdd gnd FILL
XBUFX2_insert331 BUFX2_insert331/A BUFX2_insert331/Y vdd gnd BUFX2
XBUFX2_insert342 BUFX2_insert342/A BUFX2_insert342/Y vdd gnd BUFX2
XFILL_0__12291_ vdd gnd FILL
X_13506_ _13506_/A _13506_/B _13506_/Y vdd gnd NOR2X1
X_10718_ _10718_/D _10718_/CLK _10718_/Q vdd gnd DFFPOSX1
XBUFX2_insert353 BUFX2_insert353/A BUFX2_insert353/Y vdd gnd BUFX2
X_14486_ _14486_/A _14486_/B _14486_/Y vdd gnd NAND2X1
XFILL_2__10063_ vdd gnd FILL
X_11698_ _11698_/A _11698_/B _11698_/Y vdd gnd NOR2X1
XBUFX2_insert364 BUFX2_insert364/A BUFX2_insert364/Y vdd gnd BUFX2
XFILL_0__14030_ vdd gnd FILL
XBUFX2_insert375 BUFX2_insert375/A BUFX2_insert375/Y vdd gnd BUFX2
XFILL_0__11242_ vdd gnd FILL
XFILL_1__13581_ vdd gnd FILL
XFILL_1__10793_ vdd gnd FILL
X_13437_ _13437_/D _13437_/CLK _13437_/Q vdd gnd DFFPOSX1
X_10649_ _10649_/A _10649_/B _10649_/C _10649_/Y vdd gnd OAI21X1
XFILL_1__12532_ vdd gnd FILL
XFILL_0__11173_ vdd gnd FILL
XFILL_0__7760_ vdd gnd FILL
X_13368_ _13368_/A _13368_/B _13368_/C _13368_/Y vdd gnd OAI21X1
XFILL_0__10124_ vdd gnd FILL
XFILL_1__12463_ vdd gnd FILL
X_12319_ _12319_/A _12319_/B _12319_/Y vdd gnd AND2X2
XFILL_0__7691_ vdd gnd FILL
XFILL_2__7627_ vdd gnd FILL
XFILL_1__11414_ vdd gnd FILL
X_13299_ _13299_/A _13299_/B _13299_/Y vdd gnd NAND2X1
XFILL_2__10965_ vdd gnd FILL
XFILL_0__10055_ vdd gnd FILL
XFILL_1__12394_ vdd gnd FILL
XFILL_0__9430_ vdd gnd FILL
XFILL_1__14133_ vdd gnd FILL
XFILL_2__7558_ vdd gnd FILL
XFILL_1__11345_ vdd gnd FILL
XFILL_0__14863_ vdd gnd FILL
XFILL_2__10896_ vdd gnd FILL
XFILL_2__13684_ vdd gnd FILL
XFILL_0__9361_ vdd gnd FILL
XFILL_1__14064_ vdd gnd FILL
XFILL_0__13814_ vdd gnd FILL
XFILL_2__7489_ vdd gnd FILL
XFILL_1__11276_ vdd gnd FILL
XFILL_0__14794_ vdd gnd FILL
XFILL_0__8312_ vdd gnd FILL
XFILL_0__9292_ vdd gnd FILL
X_8940_ _8940_/A _8940_/B _8940_/C _8940_/Y vdd gnd OAI21X1
XFILL_1__13015_ vdd gnd FILL
XFILL_1__10227_ vdd gnd FILL
XFILL_0__13745_ vdd gnd FILL
XFILL_0__10957_ vdd gnd FILL
XFILL_0__8243_ vdd gnd FILL
XFILL257250x216150 vdd gnd FILL
X_8871_ _8871_/D _8871_/CLK _8871_/Q vdd gnd DFFPOSX1
XFILL_1__10158_ vdd gnd FILL
XFILL_0__13676_ vdd gnd FILL
X_7822_ _7822_/A _7822_/Y vdd gnd INVX1
XFILL_0__8174_ vdd gnd FILL
XFILL_0__10888_ vdd gnd FILL
XFILL_0__12627_ vdd gnd FILL
XFILL_0__7125_ vdd gnd FILL
XFILL_1__10089_ vdd gnd FILL
X_7753_ _7753_/A _7753_/B _7753_/Y vdd gnd NAND2X1
XFILL_1__13917_ vdd gnd FILL
XFILL_2__11379_ vdd gnd FILL
X_7684_ _7684_/A _7684_/B _7684_/C _7684_/Y vdd gnd OAI21X1
XFILL_0__11509_ vdd gnd FILL
XFILL_1__13848_ vdd gnd FILL
X_9423_ _9423_/A _9423_/B _9423_/Y vdd gnd NAND2X1
XFILL_0__12489_ vdd gnd FILL
XFILL_0__14228_ vdd gnd FILL
XFILL_1__13779_ vdd gnd FILL
X_9354_ _9354_/A _9354_/B _9354_/C _9354_/Y vdd gnd OAI21X1
X_8305_ _8305_/A _8305_/B _8305_/C _8305_/Y vdd gnd OAI21X1
X_9285_ _9285_/A _9285_/B _9285_/C _9285_/Y vdd gnd OAI21X1
X_8236_ _8236_/A _8236_/B _8236_/C _8236_/Y vdd gnd NAND3X1
XFILL_1__9470_ vdd gnd FILL
XFILL_0__7889_ vdd gnd FILL
XFILL_0__9628_ vdd gnd FILL
XFILL_1__8421_ vdd gnd FILL
X_8167_ _8167_/A _8167_/B _8167_/Y vdd gnd NOR2X1
X_7118_ _7118_/A _7118_/B _7118_/Y vdd gnd NAND2X1
XFILL_0__9559_ vdd gnd FILL
XFILL_1__8352_ vdd gnd FILL
X_8098_ _8098_/A _8098_/B _8098_/C _8098_/Y vdd gnd OAI21X1
XFILL_1__7303_ vdd gnd FILL
XFILL_1__8283_ vdd gnd FILL
XFILL257250x126150 vdd gnd FILL
XFILL_1__7234_ vdd gnd FILL
XFILL_1__7165_ vdd gnd FILL
XFILL_1_BUFX2_insert306 vdd gnd FILL
XFILL_1_BUFX2_insert317 vdd gnd FILL
XFILL_1_BUFX2_insert328 vdd gnd FILL
XFILL_1_BUFX2_insert339 vdd gnd FILL
X_12670_ _12670_/A _12670_/Y vdd gnd INVX8
XFILL_1__7096_ vdd gnd FILL
X_11621_ _11621_/D _11621_/CLK _11621_/Q vdd gnd DFFPOSX1
X_14340_ _14340_/A _14340_/Y vdd gnd INVX1
X_11552_ _11552_/A _11552_/B _11552_/C _11552_/Y vdd gnd OAI21X1
X_10503_ _10503_/A _10503_/Y vdd gnd INVX1
X_14271_ _14271_/A _14271_/B _14271_/C _14271_/Y vdd gnd OAI21X1
X_11483_ _11483_/A _11483_/B _11483_/Y vdd gnd NOR2X1
XFILL_1__7998_ vdd gnd FILL
X_10434_ _10434_/A _10434_/B _10434_/Y vdd gnd OR2X2
X_13222_ _13222_/A _13222_/B _13222_/C _13222_/Y vdd gnd OAI21X1
XFILL_1__9737_ vdd gnd FILL
X_13153_ _13153_/A _13153_/Y vdd gnd INVX1
X_10365_ _10365_/A _10365_/B _10365_/C _10365_/Y vdd gnd AOI21X1
XFILL_1__9668_ vdd gnd FILL
X_12104_ _12104_/A _12104_/B _12104_/C _12104_/Y vdd gnd OAI21X1
X_13084_ _13084_/A _13084_/B _13084_/Y vdd gnd OR2X2
X_10296_ _10296_/A _10296_/B _10296_/Y vdd gnd NAND2X1
XFILL_2__7412_ vdd gnd FILL
XFILL_1__8619_ vdd gnd FILL
XFILL_1__9599_ vdd gnd FILL
X_12035_ _12035_/A _12035_/B _12035_/C _12035_/Y vdd gnd OAI21X1
XFILL_2__7343_ vdd gnd FILL
XFILL_1__11130_ vdd gnd FILL
XFILL_0__11860_ vdd gnd FILL
XFILL_2__12420_ vdd gnd FILL
XFILL_1__11061_ vdd gnd FILL
XFILL_2__7274_ vdd gnd FILL
XFILL_0__10811_ vdd gnd FILL
XFILL256950x10950 vdd gnd FILL
XFILL_0__11791_ vdd gnd FILL
XFILL_1__10012_ vdd gnd FILL
XFILL_2__12351_ vdd gnd FILL
X_13986_ _13986_/A _13986_/Y vdd gnd INVX1
XFILL_0__13530_ vdd gnd FILL
XFILL_2_BUFX2_insert151 vdd gnd FILL
X_12937_ _12937_/A _12937_/B _12937_/Y vdd gnd NAND2X1
XFILL_2_BUFX2_insert184 vdd gnd FILL
XFILL_1__14820_ vdd gnd FILL
XFILL_2__12282_ vdd gnd FILL
XFILL_0__10673_ vdd gnd FILL
X_12868_ _12868_/A _12868_/B _12868_/Y vdd gnd NOR2X1
XFILL_0__12412_ vdd gnd FILL
XFILL_1__14751_ vdd gnd FILL
XFILL_1__11963_ vdd gnd FILL
X_14607_ _14607_/A _14607_/B _14607_/Y vdd gnd NAND2X1
XFILL_0__13392_ vdd gnd FILL
X_11819_ _11819_/A _11819_/B _11819_/Y vdd gnd AND2X2
X_12799_ _12799_/A _12799_/B _12799_/Y vdd gnd NAND2X1
XFILL_1__10914_ vdd gnd FILL
XFILL_1__13702_ vdd gnd FILL
XFILL_0__12343_ vdd gnd FILL
XFILL_1__14682_ vdd gnd FILL
XFILL_1__11894_ vdd gnd FILL
XFILL_0__8930_ vdd gnd FILL
X_14538_ _14538_/D _14538_/CLK _14538_/Q vdd gnd DFFPOSX1
XFILL_2__10115_ vdd gnd FILL
XBUFX2_insert150 BUFX2_insert150/A BUFX2_insert150/Y vdd gnd BUFX2
XFILL_1__13633_ vdd gnd FILL
XBUFX2_insert161 BUFX2_insert161/A BUFX2_insert161/Y vdd gnd BUFX2
XFILL_1__10845_ vdd gnd FILL
XFILL_0__12274_ vdd gnd FILL
XBUFX2_insert172 BUFX2_insert172/A BUFX2_insert172/Y vdd gnd BUFX2
XBUFX2_insert183 BUFX2_insert183/A BUFX2_insert183/Y vdd gnd BUFX2
X_14469_ _14469_/A _14469_/B _14469_/C _14469_/Y vdd gnd OAI21X1
XFILL_2__10046_ vdd gnd FILL
XFILL_0__14013_ vdd gnd FILL
XBUFX2_insert194 BUFX2_insert194/A BUFX2_insert194/Y vdd gnd BUFX2
XFILL_1__13564_ vdd gnd FILL
XFILL_0__11225_ vdd gnd FILL
XFILL_1__10776_ vdd gnd FILL
XFILL_0__7812_ vdd gnd FILL
XFILL_1__12515_ vdd gnd FILL
XFILL_0__8792_ vdd gnd FILL
XFILL_0__11156_ vdd gnd FILL
X_9070_ _9070_/A _9070_/Y vdd gnd INVX1
XFILL_0__7743_ vdd gnd FILL
XFILL_0__10107_ vdd gnd FILL
XFILL_1__12446_ vdd gnd FILL
XFILL_0__11087_ vdd gnd FILL
X_8021_ _8021_/A _8021_/B _8021_/C _8021_/Y vdd gnd OAI21X1
XFILL_0__7674_ vdd gnd FILL
XFILL_0__14915_ vdd gnd FILL
XFILL_0__10038_ vdd gnd FILL
XFILL_1__12377_ vdd gnd FILL
XFILL_2__10948_ vdd gnd FILL
XFILL_0__9413_ vdd gnd FILL
XFILL_1__14116_ vdd gnd FILL
XFILL_1__11328_ vdd gnd FILL
XFILL_0__14846_ vdd gnd FILL
XFILL_2__10879_ vdd gnd FILL
XFILL_0__9344_ vdd gnd FILL
X_9972_ _9972_/A _9972_/B _9972_/C _9972_/Y vdd gnd OAI21X1
XFILL_1__14047_ vdd gnd FILL
XFILL_1__11259_ vdd gnd FILL
XFILL_0__14777_ vdd gnd FILL
XFILL_0__11989_ vdd gnd FILL
XFILL_0__9275_ vdd gnd FILL
X_8923_ _8923_/A _8923_/Y vdd gnd INVX2
XFILL_0__13728_ vdd gnd FILL
XFILL_0__8226_ vdd gnd FILL
X_8854_ _8854_/D _8854_/CLK _8854_/Q vdd gnd DFFPOSX1
XFILL_0__13659_ vdd gnd FILL
X_7805_ _7805_/A _7805_/B _7805_/C _7805_/Y vdd gnd OAI21X1
XFILL_0__8157_ vdd gnd FILL
X_8785_ _8785_/A _8785_/B _8785_/C _8785_/Y vdd gnd OAI21X1
XFILL_0__7108_ vdd gnd FILL
X_7736_ _7736_/A _7736_/B _7736_/Y vdd gnd NAND2X1
XFILL_0__8088_ vdd gnd FILL
XFILL_1__8970_ vdd gnd FILL
X_7667_ _7667_/A _7667_/B _7667_/Y vdd gnd AND2X2
X_9406_ _9406_/A _9406_/Y vdd gnd INVX1
XFILL_1__7852_ vdd gnd FILL
X_7598_ _7598_/A _7598_/B _7598_/C _7598_/Y vdd gnd OAI21X1
X_9337_ _9337_/A _9337_/B _9337_/C _9337_/Y vdd gnd OAI21X1
XFILL_1__7783_ vdd gnd FILL
XFILL_1__9522_ vdd gnd FILL
X_9268_ _9268_/A _9268_/B _9268_/Y vdd gnd NAND2X1
X_10150_ _10150_/A _10150_/Y vdd gnd INVX1
X_8219_ _8219_/A _8219_/B _8219_/Y vdd gnd AND2X2
XFILL_1__9453_ vdd gnd FILL
X_9199_ _9199_/A _9199_/Y vdd gnd INVX1
X_10081_ _10081_/A _10081_/B _10081_/C _10081_/Y vdd gnd NAND3X1
XFILL_1__8404_ vdd gnd FILL
XFILL_1__9384_ vdd gnd FILL
XFILL_1__8335_ vdd gnd FILL
X_13840_ _13840_/A _13840_/B _13840_/Y vdd gnd NAND2X1
XFILL_1__8266_ vdd gnd FILL
XFILL_1__7217_ vdd gnd FILL
X_13771_ _13771_/A _13771_/B _13771_/C _13771_/Y vdd gnd OAI21X1
X_10983_ _10983_/A _10983_/B _10983_/C _10983_/Y vdd gnd NAND3X1
XFILL_1__8197_ vdd gnd FILL
XFILL_1_BUFX2_insert114 vdd gnd FILL
XFILL_1_BUFX2_insert125 vdd gnd FILL
X_12722_ _12722_/A _12722_/B _12722_/S _12722_/Y vdd gnd MUX2X1
XFILL_1_BUFX2_insert136 vdd gnd FILL
XFILL_1_BUFX2_insert147 vdd gnd FILL
XFILL_1__7148_ vdd gnd FILL
XFILL_1_BUFX2_insert158 vdd gnd FILL
XFILL_1_BUFX2_insert169 vdd gnd FILL
X_12653_ _12653_/A _12653_/B _12653_/C _12653_/Y vdd gnd AOI21X1
XFILL_1__7079_ vdd gnd FILL
X_11604_ _11604_/A _11604_/B _11604_/C _11604_/Y vdd gnd OAI21X1
X_12584_ _12584_/D _12584_/CLK _12584_/Q vdd gnd DFFPOSX1
X_14323_ _14323_/A _14323_/B _14323_/C _14323_/D _14323_/Y vdd gnd AOI22X1
X_11535_ _11535_/A _11535_/Y vdd gnd INVX1
XFILL_2__9631_ vdd gnd FILL
XFILL_1__10630_ vdd gnd FILL
X_14254_ _14254_/A _14254_/B _14254_/Y vdd gnd NAND2X1
X_11466_ _11466_/A _11466_/B _11466_/Y vdd gnd NAND2X1
XFILL_0__11010_ vdd gnd FILL
XFILL_2__9562_ vdd gnd FILL
XFILL_1__10561_ vdd gnd FILL
X_13205_ _13205_/A _13205_/B _13205_/Y vdd gnd NOR2X1
X_10417_ _10417_/A _10417_/B _10417_/Y vdd gnd NAND2X1
XFILL_1__12300_ vdd gnd FILL
X_11397_ _11397_/A _11397_/B _11397_/Y vdd gnd OR2X2
X_14185_ _14185_/D _14185_/CLK _14185_/Q vdd gnd DFFPOSX1
XFILL_2__9493_ vdd gnd FILL
XFILL_1__13280_ vdd gnd FILL
XFILL_1__10492_ vdd gnd FILL
X_13136_ _13136_/A _13136_/Y vdd gnd INVX1
X_10348_ _10348_/A _10348_/B _10348_/C _10348_/Y vdd gnd OAI21X1
XFILL_1__12231_ vdd gnd FILL
XFILL_2__14570_ vdd gnd FILL
XFILL_0__12961_ vdd gnd FILL
X_10279_ _10279_/A _10279_/B _10279_/C _10279_/Y vdd gnd OAI21X1
X_13067_ _13067_/A _13067_/B _13067_/Y vdd gnd NAND2X1
XFILL_0__14700_ vdd gnd FILL
XFILL_0__11912_ vdd gnd FILL
XFILL_1__12162_ vdd gnd FILL
X_12018_ _12018_/A _12018_/B _12018_/C _12018_/Y vdd gnd NAND3X1
XFILL_0__12892_ vdd gnd FILL
XFILL_0__7390_ vdd gnd FILL
XFILL_1__11113_ vdd gnd FILL
XFILL_0__14631_ vdd gnd FILL
XFILL_0__11843_ vdd gnd FILL
XFILL_1__12093_ vdd gnd FILL
XFILL_2__12403_ vdd gnd FILL
XFILL_1__11044_ vdd gnd FILL
XFILL_0__14562_ vdd gnd FILL
XFILL_0__11774_ vdd gnd FILL
XFILL_0__9060_ vdd gnd FILL
XFILL256650x57750 vdd gnd FILL
X_13969_ _13969_/A _13969_/B _13969_/C _13969_/Y vdd gnd AOI21X1
XFILL_2__12334_ vdd gnd FILL
XFILL_0__13513_ vdd gnd FILL
XFILL_2__7188_ vdd gnd FILL
XFILL_0__8011_ vdd gnd FILL
XFILL_0__14493_ vdd gnd FILL
XFILL_1__14803_ vdd gnd FILL
XFILL_2__12265_ vdd gnd FILL
XFILL_0__10656_ vdd gnd FILL
XFILL_1__12995_ vdd gnd FILL
X_8570_ _8570_/A _8570_/B _8570_/Y vdd gnd OR2X2
XFILL_2__14004_ vdd gnd FILL
XFILL_1__14734_ vdd gnd FILL
XFILL_2__12196_ vdd gnd FILL
XFILL_1__11946_ vdd gnd FILL
XFILL_0__13375_ vdd gnd FILL
X_7521_ _7521_/A _7521_/B _7521_/C _7521_/Y vdd gnd AOI21X1
XFILL_0__10587_ vdd gnd FILL
XFILL_0__9962_ vdd gnd FILL
XFILL_0__12326_ vdd gnd FILL
XFILL_1__14665_ vdd gnd FILL
XFILL_1__11877_ vdd gnd FILL
X_7452_ _7452_/A _7452_/B _7452_/Y vdd gnd NAND2X1
XFILL_0__9893_ vdd gnd FILL
XFILL_1__13616_ vdd gnd FILL
XFILL_0__12257_ vdd gnd FILL
XFILL_1__10828_ vdd gnd FILL
XFILL_1__14596_ vdd gnd FILL
X_7383_ _7383_/A _7383_/Y vdd gnd INVX1
XFILL_2__10029_ vdd gnd FILL
XFILL_0__11208_ vdd gnd FILL
XFILL_1__13547_ vdd gnd FILL
X_9122_ _9122_/A _9122_/B _9122_/C _9122_/Y vdd gnd OAI21X1
XFILL_0__12188_ vdd gnd FILL
XFILL_0__8775_ vdd gnd FILL
XFILL_0__11139_ vdd gnd FILL
XFILL_0__7726_ vdd gnd FILL
X_9053_ _9053_/A _9053_/B _9053_/Y vdd gnd NAND2X1
XFILL_1__12429_ vdd gnd FILL
X_8004_ _8004_/A _8004_/Y vdd gnd INVX2
XFILL_0__7657_ vdd gnd FILL
XFILL_0__7588_ vdd gnd FILL
XFILL_0__14829_ vdd gnd FILL
XFILL_0__9327_ vdd gnd FILL
XFILL_1__8120_ vdd gnd FILL
X_9955_ _9955_/A _9955_/B _9955_/Y vdd gnd NAND2X1
XFILL_0__9258_ vdd gnd FILL
XFILL_1__8051_ vdd gnd FILL
X_8906_ _8906_/D _8906_/CLK _8906_/Q vdd gnd DFFPOSX1
X_9886_ _9886_/A _9886_/Y vdd gnd INVX1
XFILL_0__8209_ vdd gnd FILL
XFILL_0__9189_ vdd gnd FILL
X_8837_ _8837_/A _8837_/B _8837_/C _8837_/Y vdd gnd OAI21X1
X_8768_ _8768_/A _8768_/B _8768_/C _8768_/Y vdd gnd OAI21X1
XFILL_1__8953_ vdd gnd FILL
X_7719_ _7719_/A _7719_/B _7719_/Y vdd gnd NAND2X1
X_8699_ _8699_/A _8699_/B _8699_/Y vdd gnd NAND2X1
XFILL_1__7904_ vdd gnd FILL
X_11320_ _11320_/A _11320_/Y vdd gnd INVX1
XFILL_1__7835_ vdd gnd FILL
X_11251_ _11251_/A _11251_/B _11251_/C _11251_/Y vdd gnd AOI21X1
XFILL_1__7766_ vdd gnd FILL
X_10202_ _10202_/A _10202_/B _10202_/C _10202_/Y vdd gnd AOI21X1
XFILL_1__9505_ vdd gnd FILL
X_11182_ _11182_/A _11182_/B _11182_/C _11182_/Y vdd gnd AOI21X1
XFILL_1__7697_ vdd gnd FILL
X_10133_ _10133_/A _10133_/B _10133_/C _10133_/Y vdd gnd OAI21X1
XFILL_1__9436_ vdd gnd FILL
X_10064_ _10064_/A _10064_/B _10064_/C _10064_/Y vdd gnd AOI21X1
XFILL_1__9367_ vdd gnd FILL
XFILL_2__8160_ vdd gnd FILL
X_14872_ _14872_/D _14872_/CLK _14872_/Q vdd gnd DFFPOSX1
XFILL_1__8318_ vdd gnd FILL
XFILL_1__9298_ vdd gnd FILL
XFILL_2__8091_ vdd gnd FILL
X_13823_ _13823_/A _13823_/B _13823_/C _13823_/Y vdd gnd AOI21X1
XFILL_1__8249_ vdd gnd FILL
XFILL_2__10380_ vdd gnd FILL
X_13754_ _13754_/A _13754_/B _13754_/Y vdd gnd NAND2X1
X_10966_ _10966_/A _10966_/B _10966_/C _10966_/Y vdd gnd OAI21X1
XFILL_0__10510_ vdd gnd FILL
XFILL_0__11490_ vdd gnd FILL
X_12705_ _12705_/A _12705_/B _12705_/C _12705_/Y vdd gnd NAND3X1
X_13685_ _13685_/A _13685_/B _13685_/C _13685_/Y vdd gnd NAND3X1
XFILL_1__11800_ vdd gnd FILL
X_10897_ _10897_/A _10897_/B _10897_/Y vdd gnd OR2X2
XFILL_2__8993_ vdd gnd FILL
XFILL_0__10441_ vdd gnd FILL
XFILL_1__12780_ vdd gnd FILL
XFILL_2__11001_ vdd gnd FILL
X_12636_ _12636_/A _12636_/Y vdd gnd INVX1
XFILL_0__13160_ vdd gnd FILL
XFILL_1__11731_ vdd gnd FILL
XFILL_0__10372_ vdd gnd FILL
X_12567_ _12567_/D _12567_/CLK _12567_/Q vdd gnd DFFPOSX1
XFILL_0__12111_ vdd gnd FILL
XFILL_2__7875_ vdd gnd FILL
XFILL_1__14450_ vdd gnd FILL
X_14306_ _14306_/A _14306_/B _14306_/C _14306_/Y vdd gnd NAND3X1
XFILL_0__13091_ vdd gnd FILL
X_11518_ _11518_/A _11518_/Y vdd gnd INVX1
XFILL_1__10613_ vdd gnd FILL
X_12498_ _12498_/A _12498_/B _12498_/Y vdd gnd NAND2X1
XFILL_1__13401_ vdd gnd FILL
XFILL_1__14381_ vdd gnd FILL
XFILL_0__12042_ vdd gnd FILL
XFILL_1__11593_ vdd gnd FILL
X_14237_ _14237_/A _14237_/Y vdd gnd INVX1
X_11449_ _11449_/A _11449_/B _11449_/Y vdd gnd NAND2X1
XFILL_2__11903_ vdd gnd FILL
XFILL_1__10544_ vdd gnd FILL
XFILL_1__13332_ vdd gnd FILL
XFILL_0__8560_ vdd gnd FILL
X_14168_ _14168_/D _14168_/CLK _14168_/Q vdd gnd DFFPOSX1
XFILL_2__14622_ vdd gnd FILL
XFILL_2__11834_ vdd gnd FILL
XFILL_1__13263_ vdd gnd FILL
XFILL_1__10475_ vdd gnd FILL
X_13119_ _13119_/A _13119_/B _13119_/Y vdd gnd NAND2X1
XFILL_0__7511_ vdd gnd FILL
XFILL_0__13993_ vdd gnd FILL
XFILL_2__8427_ vdd gnd FILL
XFILL_0__8491_ vdd gnd FILL
X_14099_ _14099_/A _14099_/B _14099_/Y vdd gnd NAND2X1
XFILL_1__12214_ vdd gnd FILL
XFILL_1__13194_ vdd gnd FILL
XFILL_2__11765_ vdd gnd FILL
XFILL_0__12944_ vdd gnd FILL
XFILL_0__7442_ vdd gnd FILL
XCLKBUF1_insert389 CLKBUF1_insert389/A CLKBUF1_insert389/Y vdd gnd CLKBUF1
XFILL_2__8358_ vdd gnd FILL
XFILL_1__12145_ vdd gnd FILL
XFILL_0__12875_ vdd gnd FILL
XFILL_0__7373_ vdd gnd FILL
XFILL_0__14614_ vdd gnd FILL
XFILL_2__10647_ vdd gnd FILL
XFILL_1__12076_ vdd gnd FILL
XFILL_0__11826_ vdd gnd FILL
XFILL_0__9112_ vdd gnd FILL
X_9740_ _9740_/A _9740_/B _9740_/Y vdd gnd NAND2X1
XFILL_1__11027_ vdd gnd FILL
XFILL_0__11757_ vdd gnd FILL
XFILL_0__9043_ vdd gnd FILL
X_9671_ _9671_/A _9671_/B _9671_/Y vdd gnd NAND2X1
XFILL_2__12317_ vdd gnd FILL
XFILL_0__14476_ vdd gnd FILL
X_8622_ _8622_/A _8622_/B _8622_/C _8622_/Y vdd gnd OAI21X1
XFILL_2__12248_ vdd gnd FILL
XFILL_0__13427_ vdd gnd FILL
XFILL_0__10639_ vdd gnd FILL
XFILL_1__12978_ vdd gnd FILL
X_8553_ _8553_/A _8553_/B _8553_/Y vdd gnd NAND2X1
XFILL_1__14717_ vdd gnd FILL
XFILL_1__11929_ vdd gnd FILL
XFILL_2__12179_ vdd gnd FILL
XFILL_0__13358_ vdd gnd FILL
XFILL_0__9945_ vdd gnd FILL
X_7504_ _7504_/A _7504_/B _7504_/Y vdd gnd AND2X2
X_8484_ _8484_/A _8484_/B _8484_/Y vdd gnd NOR2X1
XFILL_0__12309_ vdd gnd FILL
XFILL_1__14648_ vdd gnd FILL
XFILL_0__13289_ vdd gnd FILL
X_7435_ _7435_/A _7435_/Y vdd gnd INVX1
XFILL_0__9876_ vdd gnd FILL
XFILL_1__14579_ vdd gnd FILL
XFILL_1__7620_ vdd gnd FILL
XFILL_0__8827_ vdd gnd FILL
X_7366_ _7366_/A _7366_/B _7366_/Y vdd gnd AND2X2
X_9105_ _9105_/A _9105_/B _9105_/C _9105_/Y vdd gnd AOI21X1
XFILL_1__7551_ vdd gnd FILL
XFILL_0__8758_ vdd gnd FILL
X_7297_ _7297_/A _7297_/B _7297_/C _7297_/Y vdd gnd OAI21X1
X_9036_ _9036_/A _9036_/B _9036_/S _9036_/Y vdd gnd MUX2X1
XFILL_0__7709_ vdd gnd FILL
XFILL_1__7482_ vdd gnd FILL
XFILL_0__8689_ vdd gnd FILL
XFILL_1__9221_ vdd gnd FILL
XFILL_1__9152_ vdd gnd FILL
XFILL_1__8103_ vdd gnd FILL
XFILL_1__9083_ vdd gnd FILL
X_9938_ _9938_/A _9938_/B _9938_/C _9938_/Y vdd gnd NAND3X1
X_10820_ _10820_/A _10820_/B _10820_/Y vdd gnd NOR2X1
XFILL_1__8034_ vdd gnd FILL
X_9869_ _9869_/A _9869_/B _9869_/C _9869_/Y vdd gnd OAI21X1
X_10751_ _10751_/D _10751_/CLK _10751_/Q vdd gnd DFFPOSX1
X_13470_ _13470_/D _13470_/CLK _13470_/Q vdd gnd DFFPOSX1
X_10682_ _10682_/A _10682_/B _10682_/C _10682_/Y vdd gnd OAI21X1
XFILL_1__9985_ vdd gnd FILL
X_12421_ _12421_/A _12421_/B _12421_/C _12421_/Y vdd gnd OAI21X1
XFILL_1__8936_ vdd gnd FILL
X_12352_ _12352_/A _12352_/B _12352_/Y vdd gnd NOR2X1
XFILL_2__7660_ vdd gnd FILL
X_11303_ _11303_/A _11303_/B _11303_/C _11303_/Y vdd gnd OAI21X1
XFILL_1__7818_ vdd gnd FILL
X_12283_ _12283_/A _12283_/B _12283_/C _12283_/Y vdd gnd OAI21X1
XFILL_2__7591_ vdd gnd FILL
XFILL_1__8798_ vdd gnd FILL
X_14022_ _14022_/A _14022_/B _14022_/Y vdd gnd NAND2X1
X_11234_ _11234_/A _11234_/B _11234_/C _11234_/Y vdd gnd OAI21X1
XFILL_1__7749_ vdd gnd FILL
XFILL_2_BUFX2_insert8 vdd gnd FILL
X_11165_ _11165_/A _11165_/B _11165_/C _11165_/Y vdd gnd OAI21X1
XFILL_1__10260_ vdd gnd FILL
XFILL_0__10990_ vdd gnd FILL
X_10116_ _10116_/A _10116_/B _10116_/Y vdd gnd NOR2X1
XFILL_1__9419_ vdd gnd FILL
XFILL_2__8212_ vdd gnd FILL
X_11096_ _11096_/A _11096_/B _11096_/Y vdd gnd NAND2X1
XFILL_1__10191_ vdd gnd FILL
X_10047_ _10047_/A _10047_/B _10047_/Y vdd gnd NAND2X1
XFILL_2__10501_ vdd gnd FILL
XFILL_2__8143_ vdd gnd FILL
XFILL_0__12660_ vdd gnd FILL
X_14855_ _14855_/A _14855_/B _14855_/C _14855_/Y vdd gnd AOI21X1
XFILL_2__13220_ vdd gnd FILL
XFILL_2__10432_ vdd gnd FILL
XFILL_2__8074_ vdd gnd FILL
XFILL_0__11611_ vdd gnd FILL
XFILL_1__13950_ vdd gnd FILL
X_13806_ _13806_/A _13806_/B _13806_/C _13806_/Y vdd gnd OAI21X1
X_14786_ _14786_/A _14786_/B _14786_/Y vdd gnd NOR2X1
XFILL_2__10363_ vdd gnd FILL
X_11998_ _11998_/A _11998_/Y vdd gnd INVX1
XFILL_0__14330_ vdd gnd FILL
XFILL_1__12901_ vdd gnd FILL
XFILL_0__11542_ vdd gnd FILL
XFILL_1__13881_ vdd gnd FILL
X_13737_ _13737_/A _13737_/B _13737_/Y vdd gnd AND2X2
X_10949_ _10949_/A _10949_/B _10949_/Y vdd gnd NAND2X1
XFILL_2__10294_ vdd gnd FILL
XFILL_0__14261_ vdd gnd FILL
XFILL_1__12832_ vdd gnd FILL
XFILL_0__11473_ vdd gnd FILL
X_13668_ _13668_/A _13668_/B _13668_/C _13668_/Y vdd gnd AOI21X1
XFILL_0__13212_ vdd gnd FILL
XFILL_2__8976_ vdd gnd FILL
XFILL_0__10424_ vdd gnd FILL
XFILL_1__12763_ vdd gnd FILL
X_12619_ _12619_/A _12619_/Y vdd gnd INVX4
X_13599_ _13599_/A _13599_/B _13599_/S _13599_/Y vdd gnd MUX2X1
XFILL_0__13143_ vdd gnd FILL
XFILL_1__11714_ vdd gnd FILL
XFILL_0__10355_ vdd gnd FILL
XFILL_0__9730_ vdd gnd FILL
XFILL_1__12694_ vdd gnd FILL
XFILL_2__7858_ vdd gnd FILL
XFILL_1__14433_ vdd gnd FILL
XFILL_0__13074_ vdd gnd FILL
X_7220_ _7220_/A _7220_/B _7220_/C _7220_/Y vdd gnd AOI21X1
XFILL_0__10286_ vdd gnd FILL
XFILL_0__9661_ vdd gnd FILL
XFILL_0__12025_ vdd gnd FILL
XFILL_2__7789_ vdd gnd FILL
XFILL_1__14364_ vdd gnd FILL
XFILL_1__11576_ vdd gnd FILL
XFILL_0__8612_ vdd gnd FILL
X_7151_ _7151_/A _7151_/Y vdd gnd INVX1
XFILL_0__9592_ vdd gnd FILL
XFILL_1__10527_ vdd gnd FILL
XFILL_1__13315_ vdd gnd FILL
XFILL_1__14295_ vdd gnd FILL
XFILL_0__8543_ vdd gnd FILL
XFILL_2__14605_ vdd gnd FILL
X_7082_ _7082_/A _7082_/B _7082_/C _7082_/D _7082_/Y vdd gnd AOI22X1
XFILL_2__11817_ vdd gnd FILL
XFILL_1__10458_ vdd gnd FILL
XFILL_1__13246_ vdd gnd FILL
XFILL_0__13976_ vdd gnd FILL
XFILL_0__8474_ vdd gnd FILL
XFILL_1__13177_ vdd gnd FILL
XFILL_2__11748_ vdd gnd FILL
XFILL_0__12927_ vdd gnd FILL
XFILL_1__10389_ vdd gnd FILL
XFILL_0__7425_ vdd gnd FILL
XFILL_1__12128_ vdd gnd FILL
XFILL_0__12858_ vdd gnd FILL
XFILL_0__7356_ vdd gnd FILL
X_7984_ _7984_/D _7984_/CLK _7984_/Q vdd gnd DFFPOSX1
XFILL_1__12059_ vdd gnd FILL
XFILL_0__11809_ vdd gnd FILL
XFILL_0__12789_ vdd gnd FILL
X_9723_ _9723_/A _9723_/B _9723_/C _9723_/Y vdd gnd OAI21X1
XFILL_0__7287_ vdd gnd FILL
XFILL_0__9026_ vdd gnd FILL
X_9654_ _9654_/A _9654_/B _9654_/Y vdd gnd NOR2X1
XFILL_0__14459_ vdd gnd FILL
X_8605_ _8605_/A _8605_/B _8605_/Y vdd gnd NOR2X1
X_9585_ _9585_/A _9585_/Y vdd gnd INVX1
X_8536_ _8536_/A _8536_/B _8536_/C _8536_/Y vdd gnd NAND3X1
XCLKBUF1_insert90 CLKBUF1_insert90/A CLKBUF1_insert90/Y vdd gnd CLKBUF1
XFILL_0__9928_ vdd gnd FILL
XFILL_1__8721_ vdd gnd FILL
X_8467_ _8467_/A _8467_/B _8467_/Y vdd gnd OR2X2
X_7418_ _7418_/A _7418_/B _7418_/Y vdd gnd NAND2X1
XFILL_0__9859_ vdd gnd FILL
XFILL_1__8652_ vdd gnd FILL
X_8398_ _8398_/A _8398_/B _8398_/S _8398_/Y vdd gnd MUX2X1
XFILL_1__7603_ vdd gnd FILL
X_7349_ _7349_/A _7349_/B _7349_/C _7349_/Y vdd gnd OAI21X1
XFILL_1__8583_ vdd gnd FILL
XFILL_1__7534_ vdd gnd FILL
X_9019_ _9019_/A _9019_/Y vdd gnd INVX8
XFILL_1__7465_ vdd gnd FILL
XFILL_1__9204_ vdd gnd FILL
X_12970_ _12970_/A _12970_/B _12970_/Y vdd gnd NAND2X1
XFILL_1__7396_ vdd gnd FILL
X_11921_ _11921_/A _11921_/B _11921_/C _11921_/Y vdd gnd NAND3X1
XFILL_1__9135_ vdd gnd FILL
X_14640_ _14640_/A _14640_/B _14640_/Y vdd gnd NOR2X1
X_11852_ _11852_/A _11852_/Y vdd gnd INVX2
XFILL_1__9066_ vdd gnd FILL
X_10803_ _10803_/A _10803_/B _10803_/C _10803_/Y vdd gnd AOI21X1
X_14571_ _14571_/A _14571_/B _14571_/Y vdd gnd NAND2X1
XFILL_1__8017_ vdd gnd FILL
X_11783_ _11783_/A _11783_/Y vdd gnd INVX2
X_13522_ _13522_/A _13522_/Y vdd gnd INVX1
X_10734_ _10734_/D _10734_/CLK _10734_/Q vdd gnd DFFPOSX1
X_13453_ _13453_/D _13453_/CLK _13453_/Q vdd gnd DFFPOSX1
X_10665_ _10665_/A _10665_/B _10665_/C _10665_/Y vdd gnd OAI21X1
XFILL_1__9968_ vdd gnd FILL
X_12404_ _12404_/A _12404_/B _12404_/Y vdd gnd NAND2X1
X_13384_ _13384_/A _13384_/B _13384_/C _13384_/Y vdd gnd OAI21X1
X_10596_ _10596_/A _10596_/B _10596_/Y vdd gnd NAND2X1
XFILL_1__9899_ vdd gnd FILL
XFILL_0__10140_ vdd gnd FILL
X_12335_ _12335_/A _12335_/B _12335_/Y vdd gnd NAND2X1
XFILL_1__11430_ vdd gnd FILL
XFILL_0__10071_ vdd gnd FILL
X_12266_ _12266_/A _12266_/B _12266_/Y vdd gnd OR2X2
XFILL_1__11361_ vdd gnd FILL
X_14005_ _14005_/A _14005_/B _14005_/Y vdd gnd AND2X2
X_11217_ _11217_/A _11217_/B _11217_/C _11217_/Y vdd gnd AOI21X1
XFILL_1__13100_ vdd gnd FILL
XFILL_1__10312_ vdd gnd FILL
X_12197_ _12197_/A _12197_/B _12197_/C _12197_/Y vdd gnd NAND3X1
XFILL_1__14080_ vdd gnd FILL
XFILL_1__11292_ vdd gnd FILL
XFILL_0__13830_ vdd gnd FILL
X_11148_ _11148_/A _11148_/B _11148_/Y vdd gnd NAND2X1
XFILL_1__13031_ vdd gnd FILL
XFILL_1__10243_ vdd gnd FILL
XFILL_0__10973_ vdd gnd FILL
XFILL_0__13761_ vdd gnd FILL
X_11079_ _11079_/A _11079_/Y vdd gnd INVX1
XFILL_1__10174_ vdd gnd FILL
XFILL_0__12712_ vdd gnd FILL
XFILL_0__7210_ vdd gnd FILL
XFILL_0__13692_ vdd gnd FILL
X_14907_ _14907_/D _14907_/CLK _14907_/Q vdd gnd DFFPOSX1
XFILL_2__8126_ vdd gnd FILL
XFILL_0__8190_ vdd gnd FILL
XFILL_0__12643_ vdd gnd FILL
XFILL_0__7141_ vdd gnd FILL
XFILL_2__13203_ vdd gnd FILL
X_14838_ _14838_/A _14838_/B _14838_/Y vdd gnd NAND2X1
XFILL_2__10415_ vdd gnd FILL
XFILL_2__8057_ vdd gnd FILL
XFILL_1__13933_ vdd gnd FILL
X_14769_ _14769_/A _14769_/B _14769_/C _14769_/Y vdd gnd AOI21X1
XFILL_0__7072_ vdd gnd FILL
XFILL_2__13134_ vdd gnd FILL
XFILL_2__10346_ vdd gnd FILL
XFILL_0__14313_ vdd gnd FILL
XFILL_0__11525_ vdd gnd FILL
XFILL_1__13864_ vdd gnd FILL
XFILL_2__10277_ vdd gnd FILL
XFILL_0__14244_ vdd gnd FILL
XFILL_2__13065_ vdd gnd FILL
XFILL_1__12815_ vdd gnd FILL
XFILL_0__11456_ vdd gnd FILL
XFILL_1__13795_ vdd gnd FILL
X_9370_ _9370_/A _9370_/Y vdd gnd INVX1
XFILL_2__8959_ vdd gnd FILL
XFILL_0__10407_ vdd gnd FILL
XFILL_0_BUFX2_insert260 vdd gnd FILL
XFILL_1__12746_ vdd gnd FILL
XFILL_0_BUFX2_insert271 vdd gnd FILL
XFILL_0__11387_ vdd gnd FILL
X_8321_ _8321_/A _8321_/B _8321_/C _8321_/Y vdd gnd AOI21X1
XFILL_0_BUFX2_insert282 vdd gnd FILL
XFILL_0__13126_ vdd gnd FILL
XFILL_0_BUFX2_insert293 vdd gnd FILL
XFILL_0__10338_ vdd gnd FILL
XFILL_0__9713_ vdd gnd FILL
XFILL_1__12677_ vdd gnd FILL
X_8252_ _8252_/A _8252_/Y vdd gnd INVX1
XFILL_1__14416_ vdd gnd FILL
XFILL_0__13057_ vdd gnd FILL
X_7203_ _7203_/A _7203_/B _7203_/C _7203_/Y vdd gnd OAI21X1
XFILL_0__10269_ vdd gnd FILL
XFILL_0__9644_ vdd gnd FILL
X_8183_ _8183_/A _8183_/Y vdd gnd INVX1
XFILL_0__12008_ vdd gnd FILL
XFILL_2_BUFX2_insert20 vdd gnd FILL
XFILL_1__14347_ vdd gnd FILL
XFILL_1__11559_ vdd gnd FILL
X_7134_ _7134_/A _7134_/Y vdd gnd INVX1
XFILL_0__9575_ vdd gnd FILL
XFILL_1__14278_ vdd gnd FILL
XFILL_0__8526_ vdd gnd FILL
XFILL_1__13229_ vdd gnd FILL
XFILL_0__13959_ vdd gnd FILL
XFILL_1__7250_ vdd gnd FILL
XFILL_0__8457_ vdd gnd FILL
XFILL_0__7408_ vdd gnd FILL
XFILL_1__7181_ vdd gnd FILL
XFILL_0__8388_ vdd gnd FILL
XFILL_0__7339_ vdd gnd FILL
X_7967_ _7967_/D _7967_/CLK _7967_/Q vdd gnd DFFPOSX1
X_9706_ _9706_/A _9706_/B _9706_/C _9706_/Y vdd gnd OAI21X1
X_7898_ _7898_/A _7898_/B _7898_/C _7898_/Y vdd gnd OAI21X1
XFILL_0__9009_ vdd gnd FILL
X_9637_ _9637_/A _9637_/B _9637_/Y vdd gnd NAND2X1
X_9568_ _9568_/A _9568_/B _9568_/C _9568_/D _9568_/Y vdd gnd OAI22X1
X_10450_ _10450_/A _10450_/B _10450_/Y vdd gnd NAND2X1
XFILL_1__9753_ vdd gnd FILL
X_8519_ _8519_/A _8519_/B _8519_/Y vdd gnd NOR2X1
X_9499_ _9499_/A _9499_/B _9499_/Y vdd gnd AND2X2
XFILL_1__8704_ vdd gnd FILL
X_10381_ _10381_/A _10381_/B _10381_/C _10381_/Y vdd gnd NAND3X1
XFILL_1__9684_ vdd gnd FILL
X_12120_ _12120_/A _12120_/B _12120_/C _12120_/Y vdd gnd NAND3X1
XFILL_1__8635_ vdd gnd FILL
XFILL256950x183750 vdd gnd FILL
X_12051_ _12051_/A _12051_/B _12051_/C _12051_/Y vdd gnd OAI21X1
XFILL_1__8566_ vdd gnd FILL
X_11002_ _11002_/A _11002_/Y vdd gnd INVX1
XFILL_1__7517_ vdd gnd FILL
XFILL_1__8497_ vdd gnd FILL
XFILL_0_CLKBUF1_insert37 vdd gnd FILL
XFILL_0_CLKBUF1_insert48 vdd gnd FILL
XFILL_1__7448_ vdd gnd FILL
XFILL_0_CLKBUF1_insert59 vdd gnd FILL
XFILL_2_BUFX2_insert322 vdd gnd FILL
X_12953_ _12953_/A _12953_/B _12953_/Y vdd gnd OR2X2
XFILL_2_BUFX2_insert344 vdd gnd FILL
XFILL_1__7379_ vdd gnd FILL
X_11904_ _11904_/A _11904_/B _11904_/C _11904_/Y vdd gnd AOI21X1
XFILL_2_BUFX2_insert377 vdd gnd FILL
XFILL_1__9118_ vdd gnd FILL
X_12884_ _12884_/A _12884_/B _12884_/C _12884_/Y vdd gnd OAI21X1
X_14623_ _14623_/A _14623_/B _14623_/C _14623_/Y vdd gnd OAI21X1
X_11835_ _11835_/A _11835_/B _11835_/C _11835_/Y vdd gnd AOI21X1
XFILL_1__9049_ vdd gnd FILL
XFILL_2__9931_ vdd gnd FILL
XFILL_1__10930_ vdd gnd FILL
X_14554_ _14554_/D _14554_/CLK _14554_/Q vdd gnd DFFPOSX1
X_11766_ _11766_/A _11766_/B _11766_/C _11766_/Y vdd gnd OAI21X1
XBUFX2_insert310 BUFX2_insert310/A BUFX2_insert310/Y vdd gnd BUFX2
XFILL_2__9862_ vdd gnd FILL
XFILL_0__11310_ vdd gnd FILL
XBUFX2_insert321 BUFX2_insert321/A BUFX2_insert321/Y vdd gnd BUFX2
XFILL_0__12290_ vdd gnd FILL
X_13505_ _13505_/A _13505_/Y vdd gnd INVX2
XFILL_1__10861_ vdd gnd FILL
X_10717_ _10717_/D _10717_/CLK _10717_/Q vdd gnd DFFPOSX1
XBUFX2_insert332 BUFX2_insert332/A BUFX2_insert332/Y vdd gnd BUFX2
XBUFX2_insert343 BUFX2_insert343/A BUFX2_insert343/Y vdd gnd BUFX2
X_14485_ _14485_/A _14485_/B _14485_/C _14485_/Y vdd gnd OAI21X1
XFILL_2__8813_ vdd gnd FILL
XBUFX2_insert354 BUFX2_insert354/A BUFX2_insert354/Y vdd gnd BUFX2
X_11697_ _11697_/A _11697_/Y vdd gnd INVX4
XBUFX2_insert365 BUFX2_insert365/A BUFX2_insert365/Y vdd gnd BUFX2
XFILL_0__11241_ vdd gnd FILL
XBUFX2_insert376 BUFX2_insert376/A BUFX2_insert376/Y vdd gnd BUFX2
XFILL_1__10792_ vdd gnd FILL
XFILL_1__13580_ vdd gnd FILL
X_13436_ _13436_/D _13436_/CLK _13436_/Q vdd gnd DFFPOSX1
X_10648_ _10648_/A _10648_/B _10648_/Y vdd gnd NAND2X1
XFILL_2__8744_ vdd gnd FILL
XFILL_1__12531_ vdd gnd FILL
XFILL_0__11172_ vdd gnd FILL
X_13367_ _13367_/A _13367_/B _13367_/C _13367_/Y vdd gnd OAI21X1
X_10579_ _10579_/A _10579_/B _10579_/Y vdd gnd NAND2X1
XFILL_0__10123_ vdd gnd FILL
XFILL_2__8675_ vdd gnd FILL
XFILL_1__12462_ vdd gnd FILL
X_12318_ _12318_/A _12318_/B _12318_/C _12318_/Y vdd gnd OAI21X1
XFILL_0__7690_ vdd gnd FILL
X_13298_ _13298_/A _13298_/B _13298_/Y vdd gnd OR2X2
XFILL_1__11413_ vdd gnd FILL
XFILL_0__10054_ vdd gnd FILL
XFILL_1__12393_ vdd gnd FILL
X_12249_ _12249_/A _12249_/B _12249_/Y vdd gnd NAND2X1
XFILL_1__14132_ vdd gnd FILL
XFILL_1__11344_ vdd gnd FILL
XFILL_0__14862_ vdd gnd FILL
XFILL_0__9360_ vdd gnd FILL
XFILL_1__14063_ vdd gnd FILL
XFILL_0__13813_ vdd gnd FILL
XFILL_1__11275_ vdd gnd FILL
XFILL_0__8311_ vdd gnd FILL
XFILL_0__14793_ vdd gnd FILL
XFILL_0__9291_ vdd gnd FILL
XFILL_1__10226_ vdd gnd FILL
XFILL_1__13014_ vdd gnd FILL
XFILL_0__13744_ vdd gnd FILL
XFILL_0__10956_ vdd gnd FILL
XFILL_0__8242_ vdd gnd FILL
XFILL_2__14304_ vdd gnd FILL
X_8870_ _8870_/D _8870_/CLK _8870_/Q vdd gnd DFFPOSX1
XFILL_1__10157_ vdd gnd FILL
XFILL_2__12496_ vdd gnd FILL
XFILL_0__10887_ vdd gnd FILL
XFILL_0__13675_ vdd gnd FILL
X_7821_ _7821_/A _7821_/B _7821_/C _7821_/Y vdd gnd AOI21X1
XFILL_0__8173_ vdd gnd FILL
XFILL_2__14235_ vdd gnd FILL
XFILL_1__10088_ vdd gnd FILL
XFILL_0__12626_ vdd gnd FILL
XFILL_0__7124_ vdd gnd FILL
X_7752_ _7752_/A _7752_/B _7752_/Y vdd gnd OR2X2
XFILL_1__13916_ vdd gnd FILL
XFILL_2__13117_ vdd gnd FILL
X_7683_ _7683_/A _7683_/B _7683_/C _7683_/Y vdd gnd OAI21X1
XFILL_2__14097_ vdd gnd FILL
XFILL_1__13847_ vdd gnd FILL
XFILL_0__11508_ vdd gnd FILL
XFILL_0__12488_ vdd gnd FILL
X_9422_ _9422_/A _9422_/B _9422_/C _9422_/Y vdd gnd AOI21X1
XFILL_2__13048_ vdd gnd FILL
XFILL_0__14227_ vdd gnd FILL
XFILL_0__11439_ vdd gnd FILL
XFILL_1__13778_ vdd gnd FILL
X_9353_ _9353_/A _9353_/B _9353_/Y vdd gnd NOR2X1
XFILL_1__12729_ vdd gnd FILL
XFILL_0__14158_ vdd gnd FILL
X_8304_ _8304_/A _8304_/Y vdd gnd INVX1
X_9284_ _9284_/A _9284_/B _9284_/Y vdd gnd NAND2X1
XFILL_0__13109_ vdd gnd FILL
XFILL_0__14089_ vdd gnd FILL
X_8235_ _8235_/A _8235_/B _8235_/Y vdd gnd NAND2X1
XFILL_0__7888_ vdd gnd FILL
XFILL_0__9627_ vdd gnd FILL
XFILL_1__8420_ vdd gnd FILL
X_8166_ _8166_/A _8166_/B _8166_/Y vdd gnd NOR2X1
X_7117_ _7117_/A _7117_/Y vdd gnd INVX1
XFILL_0__9558_ vdd gnd FILL
XFILL_1__8351_ vdd gnd FILL
X_8097_ _8097_/A _8097_/B _8097_/Y vdd gnd NAND2X1
XFILL256950x115350 vdd gnd FILL
XFILL_1__7302_ vdd gnd FILL
XFILL_0__8509_ vdd gnd FILL
XFILL_0__9489_ vdd gnd FILL
XFILL_1__8282_ vdd gnd FILL
XFILL_1__7233_ vdd gnd FILL
XFILL_1__7164_ vdd gnd FILL
XFILL_1_BUFX2_insert307 vdd gnd FILL
X_8999_ _8999_/A _8999_/Y vdd gnd INVX1
XFILL_1_BUFX2_insert318 vdd gnd FILL
XFILL_1_BUFX2_insert329 vdd gnd FILL
XFILL_1__7095_ vdd gnd FILL
X_11620_ _11620_/D _11620_/CLK _11620_/Q vdd gnd DFFPOSX1
X_11551_ _11551_/A _11551_/B _11551_/C _11551_/Y vdd gnd OAI21X1
X_10502_ _10502_/A _10502_/B _10502_/Y vdd gnd NAND2X1
X_14270_ _14270_/A _14270_/B _14270_/C _14270_/Y vdd gnd OAI21X1
X_11482_ _11482_/A _11482_/B _11482_/Y vdd gnd NAND2X1
XFILL_1__7997_ vdd gnd FILL
X_13221_ _13221_/A _13221_/B _13221_/C _13221_/Y vdd gnd OAI21X1
X_10433_ _10433_/A _10433_/Y vdd gnd INVX1
XFILL_1__9736_ vdd gnd FILL
X_13152_ _13152_/A _13152_/B _13152_/Y vdd gnd NOR2X1
X_10364_ _10364_/A _10364_/B _10364_/C _10364_/Y vdd gnd NAND3X1
XFILL_1__9667_ vdd gnd FILL
XFILL_2__8460_ vdd gnd FILL
X_12103_ _12103_/A _12103_/B _12103_/C _12103_/Y vdd gnd AOI21X1
X_13083_ _13083_/A _13083_/B _13083_/Y vdd gnd NAND2X1
XFILL_1__8618_ vdd gnd FILL
X_10295_ _10295_/A _10295_/B _10295_/C _10295_/Y vdd gnd NAND3X1
XFILL_1__9598_ vdd gnd FILL
XFILL_2__8391_ vdd gnd FILL
X_12034_ _12034_/A _12034_/B _12034_/C _12034_/Y vdd gnd OAI21X1
XFILL_1__8549_ vdd gnd FILL
XFILL_2__10680_ vdd gnd FILL
XFILL_1__11060_ vdd gnd FILL
XFILL_0__10810_ vdd gnd FILL
XFILL_0__11790_ vdd gnd FILL
XFILL_2__9012_ vdd gnd FILL
XFILL_1__10011_ vdd gnd FILL
X_13985_ _13985_/A _13985_/B _13985_/C _13985_/Y vdd gnd OAI21X1
XFILL_2_BUFX2_insert141 vdd gnd FILL
XFILL_2_BUFX2_insert163 vdd gnd FILL
X_12936_ _12936_/A _12936_/B _12936_/Y vdd gnd NAND2X1
XFILL_2__11301_ vdd gnd FILL
XFILL_2_BUFX2_insert196 vdd gnd FILL
XFILL_0__10672_ vdd gnd FILL
X_12867_ _12867_/A _12867_/Y vdd gnd INVX1
XFILL_2__14020_ vdd gnd FILL
XFILL_2__11232_ vdd gnd FILL
XFILL_1__14750_ vdd gnd FILL
XFILL_0__12411_ vdd gnd FILL
XFILL_1__11962_ vdd gnd FILL
XFILL_0__13391_ vdd gnd FILL
X_14606_ _14606_/A _14606_/B _14606_/Y vdd gnd NAND2X1
X_11818_ _11818_/A _11818_/B _11818_/C _11818_/Y vdd gnd NAND3X1
XFILL_2__9914_ vdd gnd FILL
X_12798_ _12798_/A _12798_/B _12798_/C _12798_/Y vdd gnd OAI21X1
XFILL_1__13701_ vdd gnd FILL
XFILL_2__11163_ vdd gnd FILL
XFILL_0__12342_ vdd gnd FILL
XFILL_1__10913_ vdd gnd FILL
XFILL_1__14681_ vdd gnd FILL
XFILL_1__11893_ vdd gnd FILL
X_14537_ _14537_/D _14537_/CLK _14537_/Q vdd gnd DFFPOSX1
X_11749_ _11749_/A _11749_/B _11749_/C _11749_/Y vdd gnd OAI21X1
XBUFX2_insert140 BUFX2_insert140/A BUFX2_insert140/Y vdd gnd BUFX2
XFILL_1__13632_ vdd gnd FILL
XFILL_2__9845_ vdd gnd FILL
XBUFX2_insert151 BUFX2_insert151/A BUFX2_insert151/Y vdd gnd BUFX2
XFILL_2__11094_ vdd gnd FILL
XFILL_0__12273_ vdd gnd FILL
XFILL_1__10844_ vdd gnd FILL
XBUFX2_insert162 BUFX2_insert162/A BUFX2_insert162/Y vdd gnd BUFX2
X_14468_ _14468_/A _14468_/B _14468_/Y vdd gnd NAND2X1
XBUFX2_insert173 BUFX2_insert173/A BUFX2_insert173/Y vdd gnd BUFX2
XBUFX2_insert184 BUFX2_insert184/A BUFX2_insert184/Y vdd gnd BUFX2
XFILL_0__11224_ vdd gnd FILL
XFILL_0__14012_ vdd gnd FILL
XBUFX2_insert195 BUFX2_insert195/A BUFX2_insert195/Y vdd gnd BUFX2
XFILL_1__13563_ vdd gnd FILL
XFILL_0__7811_ vdd gnd FILL
X_13419_ _13419_/A _13419_/B _13419_/C _13419_/Y vdd gnd OAI21X1
XFILL_1__10775_ vdd gnd FILL
XFILL_0__8791_ vdd gnd FILL
X_14399_ _14399_/A _14399_/B _14399_/Y vdd gnd NAND2X1
XFILL_2__14853_ vdd gnd FILL
XFILL_2__8727_ vdd gnd FILL
XFILL_1__12514_ vdd gnd FILL
XFILL_0__11155_ vdd gnd FILL
XFILL_0__7742_ vdd gnd FILL
XFILL_2__13804_ vdd gnd FILL
XFILL_0__10106_ vdd gnd FILL
XFILL_2__8658_ vdd gnd FILL
XFILL_2__14784_ vdd gnd FILL
XFILL_1__12445_ vdd gnd FILL
XFILL_0__11086_ vdd gnd FILL
XFILL_2__11996_ vdd gnd FILL
X_8020_ _8020_/A _8020_/Y vdd gnd INVX1
XFILL_0__7673_ vdd gnd FILL
XFILL_0__10037_ vdd gnd FILL
XFILL_0__14914_ vdd gnd FILL
XFILL_2__8589_ vdd gnd FILL
XFILL_0__9412_ vdd gnd FILL
XFILL_1__12376_ vdd gnd FILL
XFILL_1__14115_ vdd gnd FILL
XFILL_1__11327_ vdd gnd FILL
XFILL_0__14845_ vdd gnd FILL
XFILL_0__9343_ vdd gnd FILL
X_9971_ _9971_/A _9971_/B _9971_/Y vdd gnd AND2X2
XFILL_2__12617_ vdd gnd FILL
XFILL_1__14046_ vdd gnd FILL
XFILL_1__11258_ vdd gnd FILL
XFILL_0__14776_ vdd gnd FILL
XFILL_0__9274_ vdd gnd FILL
X_8922_ _8922_/A _8922_/B _8922_/Y vdd gnd NOR2X1
XFILL_0__11988_ vdd gnd FILL
XFILL_1__10209_ vdd gnd FILL
XFILL_0__13727_ vdd gnd FILL
XFILL_1__11189_ vdd gnd FILL
XFILL_0__8225_ vdd gnd FILL
XFILL_0__10939_ vdd gnd FILL
X_8853_ _8853_/D _8853_/CLK _8853_/Q vdd gnd DFFPOSX1
XFILL_2__12479_ vdd gnd FILL
XFILL_0__13658_ vdd gnd FILL
X_7804_ _7804_/A _7804_/B _7804_/C _7804_/Y vdd gnd NAND3X1
XFILL_0__8156_ vdd gnd FILL
XFILL_2__14218_ vdd gnd FILL
X_8784_ _8784_/A _8784_/B _8784_/Y vdd gnd NAND2X1
XFILL_0__7107_ vdd gnd FILL
XFILL_0__13589_ vdd gnd FILL
X_7735_ _7735_/A _7735_/B _7735_/Y vdd gnd NOR2X1
XFILL_0__8087_ vdd gnd FILL
XFILL_2__14149_ vdd gnd FILL
X_7666_ _7666_/A _7666_/B _7666_/C _7666_/Y vdd gnd NAND3X1
X_9405_ _9405_/A _9405_/B _9405_/C _9405_/Y vdd gnd OAI21X1
XFILL_1__7851_ vdd gnd FILL
X_7597_ _7597_/A _7597_/B _7597_/Y vdd gnd NAND2X1
X_9336_ _9336_/A _9336_/B _9336_/Y vdd gnd NAND2X1
XFILL_0__8989_ vdd gnd FILL
XFILL_1__7782_ vdd gnd FILL
XFILL_1__9521_ vdd gnd FILL
X_9267_ _9267_/A _9267_/Y vdd gnd INVX1
XFILL_1__9452_ vdd gnd FILL
X_8218_ _8218_/A _8218_/B _8218_/Y vdd gnd NAND2X1
X_9198_ _9198_/A _9198_/B _9198_/C _9198_/Y vdd gnd OAI21X1
XFILL_1__8403_ vdd gnd FILL
X_10080_ _10080_/A _10080_/B _10080_/Y vdd gnd NAND2X1
XFILL_1__9383_ vdd gnd FILL
X_8149_ _8149_/A _8149_/Y vdd gnd INVX1
XFILL_1__8334_ vdd gnd FILL
XFILL_1__8265_ vdd gnd FILL
XFILL_1__7216_ vdd gnd FILL
X_13770_ _13770_/A _13770_/B _13770_/Y vdd gnd OR2X2
X_10982_ _10982_/A _10982_/B _10982_/C _10982_/Y vdd gnd OAI21X1
XFILL_1__8196_ vdd gnd FILL
X_12721_ _12721_/A _12721_/B _12721_/C _12721_/Y vdd gnd OAI21X1
XFILL_1_BUFX2_insert115 vdd gnd FILL
XFILL_1__7147_ vdd gnd FILL
XFILL_1_BUFX2_insert126 vdd gnd FILL
XFILL_1_BUFX2_insert137 vdd gnd FILL
XFILL_1_BUFX2_insert148 vdd gnd FILL
XFILL_1_BUFX2_insert159 vdd gnd FILL
X_12652_ _12652_/A _12652_/B _12652_/C _12652_/Y vdd gnd OAI21X1
XFILL_1__7078_ vdd gnd FILL
X_11603_ _11603_/A _11603_/B _11603_/C _11603_/Y vdd gnd OAI21X1
X_12583_ _12583_/D _12583_/CLK _12583_/Q vdd gnd DFFPOSX1
XFILL_2__7891_ vdd gnd FILL
X_14322_ _14322_/A _14322_/B _14322_/C _14322_/Y vdd gnd AOI21X1
X_11534_ _11534_/A _11534_/B _11534_/C _11534_/Y vdd gnd OAI21X1
X_14253_ _14253_/A _14253_/Y vdd gnd INVX8
X_11465_ _11465_/A _11465_/B _11465_/Y vdd gnd NOR2X1
X_13204_ _13204_/A _13204_/B _13204_/Y vdd gnd AND2X2
XFILL_1__10560_ vdd gnd FILL
X_10416_ _10416_/A _10416_/B _10416_/C _10416_/Y vdd gnd OAI21X1
XFILL_2__8512_ vdd gnd FILL
X_14184_ _14184_/D _14184_/CLK _14184_/Q vdd gnd DFFPOSX1
XFILL_1__9719_ vdd gnd FILL
X_11396_ _11396_/A _11396_/B _11396_/Y vdd gnd OR2X2
XFILL_2__11850_ vdd gnd FILL
XFILL_1__10491_ vdd gnd FILL
X_13135_ _13135_/A _13135_/B _13135_/C _13135_/Y vdd gnd OAI21X1
X_10347_ _10347_/A _10347_/B _10347_/Y vdd gnd NAND2X1
XFILL_2__8443_ vdd gnd FILL
XFILL_1__12230_ vdd gnd FILL
XFILL_2__11781_ vdd gnd FILL
XFILL_0__12960_ vdd gnd FILL
X_13066_ _13066_/A _13066_/B _13066_/C _13066_/Y vdd gnd AOI21X1
X_10278_ _10278_/A _10278_/B _10278_/C _10278_/Y vdd gnd OAI21X1
XFILL_2__13520_ vdd gnd FILL
XFILL_2__8374_ vdd gnd FILL
XFILL_0__11911_ vdd gnd FILL
XFILL_1__12161_ vdd gnd FILL
X_12017_ _12017_/A _12017_/B _12017_/C _12017_/Y vdd gnd AOI21X1
XFILL_0__12891_ vdd gnd FILL
XFILL_1__11112_ vdd gnd FILL
XFILL_0__14630_ vdd gnd FILL
XFILL_2__10663_ vdd gnd FILL
XFILL_1__12092_ vdd gnd FILL
XFILL_0__11842_ vdd gnd FILL
XFILL_1__11043_ vdd gnd FILL
XFILL_2__13382_ vdd gnd FILL
XFILL_0__14561_ vdd gnd FILL
XFILL_2__10594_ vdd gnd FILL
XFILL_0__11773_ vdd gnd FILL
X_13968_ _13968_/A _13968_/B _13968_/Y vdd gnd NOR2X1
XFILL_0__13512_ vdd gnd FILL
XFILL_0__8010_ vdd gnd FILL
XFILL_0__14492_ vdd gnd FILL
X_12919_ _12919_/A _12919_/B _12919_/C _12919_/Y vdd gnd NAND3X1
XFILL_1__14802_ vdd gnd FILL
X_13899_ _13899_/A _13899_/B _13899_/Y vdd gnd NAND2X1
XFILL_0__10655_ vdd gnd FILL
XFILL_1__12994_ vdd gnd FILL
XFILL_2__11215_ vdd gnd FILL
XFILL_1__14733_ vdd gnd FILL
XFILL_1__11945_ vdd gnd FILL
XFILL_0__10586_ vdd gnd FILL
XFILL_0__13374_ vdd gnd FILL
X_7520_ _7520_/A _7520_/B _7520_/C _7520_/Y vdd gnd OAI21X1
XFILL_0__9961_ vdd gnd FILL
XFILL_2__11146_ vdd gnd FILL
XFILL_1__14664_ vdd gnd FILL
XFILL_0__12325_ vdd gnd FILL
XFILL_1__11876_ vdd gnd FILL
X_7451_ _7451_/A _7451_/B _7451_/Y vdd gnd NAND2X1
XFILL_0__9892_ vdd gnd FILL
XFILL_1__13615_ vdd gnd FILL
XFILL_2__11077_ vdd gnd FILL
XFILL_0__12256_ vdd gnd FILL
XFILL_1__10827_ vdd gnd FILL
XFILL_1__14595_ vdd gnd FILL
X_7382_ _7382_/A _7382_/B _7382_/C _7382_/Y vdd gnd NAND3X1
XFILL_0__11207_ vdd gnd FILL
XFILL_1__13546_ vdd gnd FILL
XFILL_0__12187_ vdd gnd FILL
X_9121_ _9121_/A _9121_/B _9121_/Y vdd gnd AND2X2
XFILL_0__8774_ vdd gnd FILL
XFILL_2__14836_ vdd gnd FILL
XFILL_0__11138_ vdd gnd FILL
XFILL_0__7725_ vdd gnd FILL
X_9052_ _9052_/A _9052_/Y vdd gnd INVX1
XFILL_2__14767_ vdd gnd FILL
XFILL_1__12428_ vdd gnd FILL
XFILL_0__11069_ vdd gnd FILL
XFILL_2__11979_ vdd gnd FILL
X_8003_ _8003_/A _8003_/B _8003_/C _8003_/Y vdd gnd OAI21X1
XFILL_0__7656_ vdd gnd FILL
XFILL_2__13718_ vdd gnd FILL
XFILL_2__14698_ vdd gnd FILL
XFILL_1__12359_ vdd gnd FILL
XFILL_0__7587_ vdd gnd FILL
XFILL_2__13649_ vdd gnd FILL
XFILL_0__14828_ vdd gnd FILL
XFILL_0__9326_ vdd gnd FILL
X_9954_ _9954_/A _9954_/Y vdd gnd INVX1
XFILL_1__14029_ vdd gnd FILL
XFILL_0__14759_ vdd gnd FILL
XFILL_0__9257_ vdd gnd FILL
XFILL_1__8050_ vdd gnd FILL
X_8905_ _8905_/D _8905_/CLK _8905_/Q vdd gnd DFFPOSX1
X_9885_ _9885_/A _9885_/B _9885_/Y vdd gnd NAND2X1
XFILL_0__8208_ vdd gnd FILL
XFILL_0__9188_ vdd gnd FILL
X_8836_ _8836_/A _8836_/B _8836_/Y vdd gnd NAND2X1
XFILL_0__8139_ vdd gnd FILL
X_8767_ _8767_/A _8767_/Y vdd gnd INVX1
X_7718_ _7718_/A _7718_/B _7718_/Y vdd gnd NAND2X1
XFILL_1__8952_ vdd gnd FILL
X_8698_ _8698_/A _8698_/B _8698_/Y vdd gnd OR2X2
XFILL_1__7903_ vdd gnd FILL
X_7649_ _7649_/A _7649_/B _7649_/Y vdd gnd NAND2X1
XFILL_1__7834_ vdd gnd FILL
X_11250_ _11250_/A _11250_/B _11250_/Y vdd gnd NOR2X1
X_9319_ _9319_/A _9319_/B _9319_/C _9319_/Y vdd gnd OAI21X1
XFILL_1__7765_ vdd gnd FILL
X_10201_ _10201_/A _10201_/B _10201_/C _10201_/Y vdd gnd NOR3X1
XFILL_1__9504_ vdd gnd FILL
X_11181_ _11181_/A _11181_/B _11181_/Y vdd gnd NAND2X1
XFILL_1__7696_ vdd gnd FILL
X_10132_ _10132_/A _10132_/Y vdd gnd INVX1
XFILL_1__9435_ vdd gnd FILL
X_10063_ _10063_/A _10063_/B _10063_/C _10063_/Y vdd gnd NAND3X1
XFILL_1__9366_ vdd gnd FILL
XFILL_2__7110_ vdd gnd FILL
XFILL_1__8317_ vdd gnd FILL
X_14871_ _14871_/D _14871_/CLK _14871_/Q vdd gnd DFFPOSX1
XFILL_1__9297_ vdd gnd FILL
X_13822_ _13822_/A _13822_/B _13822_/C _13822_/Y vdd gnd AOI21X1
XFILL_1__8248_ vdd gnd FILL
X_13753_ _13753_/A _13753_/B _13753_/C _13753_/Y vdd gnd NAND3X1
X_10965_ _10965_/A _10965_/B _10965_/Y vdd gnd NOR2X1
XFILL_1__8179_ vdd gnd FILL
X_12704_ _12704_/A _12704_/B _12704_/C _12704_/Y vdd gnd NAND3X1
X_13684_ _13684_/A _13684_/B _13684_/C _13684_/Y vdd gnd OAI21X1
X_10896_ _10896_/A _10896_/B _10896_/C _10896_/Y vdd gnd OAI21X1
XFILL_0__10440_ vdd gnd FILL
X_12635_ _12635_/A _12635_/B _12635_/C _12635_/Y vdd gnd AOI21X1
XFILL_1__11730_ vdd gnd FILL
XFILL_0__10371_ vdd gnd FILL
X_12566_ _12566_/D _12566_/CLK _12566_/Q vdd gnd DFFPOSX1
XFILL_0__12110_ vdd gnd FILL
XFILL_0__13090_ vdd gnd FILL
X_14305_ _14305_/A _14305_/B _14305_/Y vdd gnd NAND2X1
X_11517_ _11517_/A _11517_/B _11517_/C _11517_/Y vdd gnd AOI21X1
X_12497_ _12497_/A _12497_/B _12497_/C _12497_/Y vdd gnd OAI21X1
XFILL_1__13400_ vdd gnd FILL
XFILL_1__10612_ vdd gnd FILL
XFILL_0__12041_ vdd gnd FILL
XFILL_1__14380_ vdd gnd FILL
X_14236_ _14236_/A _14236_/B _14236_/C _14236_/Y vdd gnd OAI21X1
XFILL_1__11592_ vdd gnd FILL
X_11448_ _11448_/A _11448_/B _11448_/Y vdd gnd OR2X2
XFILL_1__13331_ vdd gnd FILL
XFILL_1__10543_ vdd gnd FILL
X_14167_ _14167_/D _14167_/CLK _14167_/Q vdd gnd DFFPOSX1
X_11379_ _11379_/A _11379_/B _11379_/C _11379_/Y vdd gnd OAI21X1
XFILL_1__13262_ vdd gnd FILL
X_13118_ _13118_/A _13118_/B _13118_/Y vdd gnd NAND2X1
XFILL_0__7510_ vdd gnd FILL
XFILL_1__10474_ vdd gnd FILL
XFILL_0__13992_ vdd gnd FILL
XFILL_0__8490_ vdd gnd FILL
X_14098_ _14098_/A _14098_/B _14098_/C _14098_/Y vdd gnd OAI21X1
XFILL_1__12213_ vdd gnd FILL
XFILL_1__13193_ vdd gnd FILL
XFILL_0__12943_ vdd gnd FILL
XFILL_0__7441_ vdd gnd FILL
X_13049_ _13049_/A _13049_/B _13049_/S _13049_/Y vdd gnd MUX2X1
XFILL_2__13503_ vdd gnd FILL
XFILL_2__14483_ vdd gnd FILL
XFILL_1__12144_ vdd gnd FILL
XFILL_2__11695_ vdd gnd FILL
XFILL_0__12874_ vdd gnd FILL
XFILL_0__7372_ vdd gnd FILL
XFILL_2__7308_ vdd gnd FILL
XFILL_0__14613_ vdd gnd FILL
XFILL_2__8288_ vdd gnd FILL
XFILL_0__9111_ vdd gnd FILL
XFILL_1__12075_ vdd gnd FILL
XFILL_0__11825_ vdd gnd FILL
XFILL_2__7239_ vdd gnd FILL
XFILL_2__13365_ vdd gnd FILL
XFILL_1__11026_ vdd gnd FILL
XFILL_2__10577_ vdd gnd FILL
XFILL_0__9042_ vdd gnd FILL
XFILL_0__11756_ vdd gnd FILL
X_9670_ _9670_/A _9670_/Y vdd gnd INVX1
XFILL_2__13296_ vdd gnd FILL
XFILL_0__14475_ vdd gnd FILL
X_8621_ _8621_/A _8621_/B _8621_/Y vdd gnd NOR2X1
XFILL_0__13426_ vdd gnd FILL
XFILL_0__10638_ vdd gnd FILL
XFILL_1__12977_ vdd gnd FILL
X_8552_ _8552_/A _8552_/B _8552_/C _8552_/Y vdd gnd OAI21X1
XFILL_1__14716_ vdd gnd FILL
XFILL_1__11928_ vdd gnd FILL
XFILL_0__13357_ vdd gnd FILL
X_7503_ _7503_/A _7503_/B _7503_/Y vdd gnd NOR2X1
XFILL_0__10569_ vdd gnd FILL
XFILL_0__9944_ vdd gnd FILL
X_8483_ _8483_/A _8483_/B _8483_/C _8483_/Y vdd gnd NAND3X1
XFILL_2__11129_ vdd gnd FILL
XFILL_1__14647_ vdd gnd FILL
XFILL_0__12308_ vdd gnd FILL
XFILL_1__11859_ vdd gnd FILL
XFILL_0__13288_ vdd gnd FILL
X_7434_ _7434_/A _7434_/B _7434_/Y vdd gnd NAND2X1
XFILL_0__9875_ vdd gnd FILL
XFILL_1__14578_ vdd gnd FILL
XFILL_0__12239_ vdd gnd FILL
XFILL_0__8826_ vdd gnd FILL
X_7365_ _7365_/A _7365_/B _7365_/C _7365_/Y vdd gnd NAND3X1
XFILL_1__13529_ vdd gnd FILL
X_9104_ _9104_/A _9104_/B _9104_/C _9104_/D _9104_/Y vdd gnd AOI22X1
XFILL_1__7550_ vdd gnd FILL
XFILL_0__8757_ vdd gnd FILL
X_7296_ _7296_/A _7296_/B _7296_/C _7296_/Y vdd gnd OAI21X1
XFILL_0__7708_ vdd gnd FILL
X_9035_ _9035_/A _9035_/B _9035_/C _9035_/Y vdd gnd NAND3X1
XFILL_1__7481_ vdd gnd FILL
XFILL_0__8688_ vdd gnd FILL
XFILL_1__9220_ vdd gnd FILL
XFILL_0__7639_ vdd gnd FILL
XFILL_1__9151_ vdd gnd FILL
XFILL_1__8102_ vdd gnd FILL
XFILL_0__9309_ vdd gnd FILL
XFILL_1__9082_ vdd gnd FILL
X_9937_ _9937_/A _9937_/B _9937_/C _9937_/Y vdd gnd AOI21X1
XFILL_1__8033_ vdd gnd FILL
X_9868_ _9868_/A _9868_/Y vdd gnd INVX1
X_10750_ _10750_/D _10750_/CLK _10750_/Q vdd gnd DFFPOSX1
X_8819_ _8819_/A _8819_/B _8819_/C _8819_/Y vdd gnd OAI21X1
X_9799_ _9799_/D _9799_/CLK _9799_/Q vdd gnd DFFPOSX1
X_10681_ _10681_/A _10681_/B _10681_/C _10681_/Y vdd gnd OAI21X1
XFILL_1__9984_ vdd gnd FILL
X_12420_ _12420_/A _12420_/B _12420_/Y vdd gnd NOR2X1
XFILL_1__8935_ vdd gnd FILL
X_12351_ _12351_/A _12351_/Y vdd gnd INVX1
XFILL_1_CLKBUF1_insert100 vdd gnd FILL
X_11302_ _11302_/A _11302_/Y vdd gnd INVX1
X_12282_ _12282_/A _12282_/B _12282_/Y vdd gnd OR2X2
XFILL_1__7817_ vdd gnd FILL
XFILL_1__8797_ vdd gnd FILL
X_14021_ _14021_/A _14021_/B _14021_/C _14021_/Y vdd gnd OAI21X1
X_11233_ _11233_/A _11233_/B _11233_/C _11233_/Y vdd gnd NAND3X1
XFILL_1__7748_ vdd gnd FILL
X_11164_ _11164_/A _11164_/B _11164_/Y vdd gnd NAND2X1
XFILL_2__9260_ vdd gnd FILL
XFILL_1__7679_ vdd gnd FILL
X_10115_ _10115_/A _10115_/Y vdd gnd INVX1
XFILL_1__9418_ vdd gnd FILL
X_11095_ _11095_/A _11095_/B _11095_/Y vdd gnd NAND2X1
XFILL_2__9191_ vdd gnd FILL
XFILL_1__10190_ vdd gnd FILL
X_10046_ _10046_/A _10046_/B _10046_/C _10046_/Y vdd gnd OAI21X1
XFILL_1__9349_ vdd gnd FILL
XFILL_2__11480_ vdd gnd FILL
X_14854_ _14854_/A _14854_/B _14854_/C _14854_/Y vdd gnd OAI21X1
XFILL_0__11610_ vdd gnd FILL
X_13805_ _13805_/A _13805_/B _13805_/C _13805_/Y vdd gnd OAI21X1
XFILL_2__13150_ vdd gnd FILL
X_14785_ _14785_/A _14785_/B _14785_/Y vdd gnd NAND2X1
X_11997_ _11997_/A _11997_/B _11997_/C _11997_/Y vdd gnd AOI21X1
XFILL_1__12900_ vdd gnd FILL
XFILL_0__11541_ vdd gnd FILL
XFILL_1__13880_ vdd gnd FILL
XFILL_2__12101_ vdd gnd FILL
X_13736_ _13736_/A _13736_/B _13736_/C _13736_/Y vdd gnd AOI21X1
X_10948_ _10948_/A _10948_/Y vdd gnd INVX1
XFILL_2__13081_ vdd gnd FILL
XFILL_1__12831_ vdd gnd FILL
XFILL_0__14260_ vdd gnd FILL
XFILL_0__11472_ vdd gnd FILL
X_13667_ _13667_/A _13667_/B _13667_/Y vdd gnd NAND2X1
X_10879_ _10879_/A _10879_/B _10879_/Y vdd gnd NAND2X1
XFILL_0__13211_ vdd gnd FILL
XFILL_0__10423_ vdd gnd FILL
XFILL_1__12762_ vdd gnd FILL
X_12618_ _12618_/A _12618_/Y vdd gnd INVX2
X_13598_ _13598_/A _13598_/B _13598_/C _13598_/Y vdd gnd OAI21X1
XFILL_1__11713_ vdd gnd FILL
XFILL_0__13142_ vdd gnd FILL
XFILL_0__10354_ vdd gnd FILL
XFILL_1__12693_ vdd gnd FILL
X_12549_ _12549_/D _12549_/CLK _12549_/Q vdd gnd DFFPOSX1
XFILL_1__14432_ vdd gnd FILL
XFILL_0__13073_ vdd gnd FILL
XFILL_0__10285_ vdd gnd FILL
XFILL_0__9660_ vdd gnd FILL
XFILL_2__12934_ vdd gnd FILL
XFILL_0__12024_ vdd gnd FILL
XFILL_1__14363_ vdd gnd FILL
XFILL_0__8611_ vdd gnd FILL
XFILL_1__11575_ vdd gnd FILL
X_14219_ _14219_/A _14219_/Y vdd gnd INVX1
X_7150_ _7150_/A _7150_/B _7150_/Y vdd gnd NAND2X1
XFILL_0__9591_ vdd gnd FILL
XFILL256650x216150 vdd gnd FILL
XFILL_2__9527_ vdd gnd FILL
XFILL_1__13314_ vdd gnd FILL
XFILL_1__10526_ vdd gnd FILL
XFILL_1__14294_ vdd gnd FILL
XFILL_0__8542_ vdd gnd FILL
X_7081_ _7081_/A _7081_/B _7081_/Y vdd gnd AND2X2
XFILL_2__9458_ vdd gnd FILL
XFILL_1__13245_ vdd gnd FILL
XFILL_1__10457_ vdd gnd FILL
XFILL_0__13975_ vdd gnd FILL
XFILL_0__8473_ vdd gnd FILL
XFILL_1__13176_ vdd gnd FILL
XFILL_0__12926_ vdd gnd FILL
XFILL_1__10388_ vdd gnd FILL
XFILL_0__7424_ vdd gnd FILL
XFILL_2__14466_ vdd gnd FILL
XFILL_1__12127_ vdd gnd FILL
XFILL_0__12857_ vdd gnd FILL
XFILL_0__7355_ vdd gnd FILL
XFILL257250x244950 vdd gnd FILL
XFILL_2__13417_ vdd gnd FILL
X_7983_ _7983_/D _7983_/CLK _7983_/Q vdd gnd DFFPOSX1
XFILL_2__14397_ vdd gnd FILL
XFILL_1__12058_ vdd gnd FILL
XFILL_0__11808_ vdd gnd FILL
X_9722_ _9722_/A _9722_/B _9722_/Y vdd gnd NAND2X1
XFILL_0__12788_ vdd gnd FILL
XFILL_0__7286_ vdd gnd FILL
XFILL_1__11009_ vdd gnd FILL
XFILL_2__13348_ vdd gnd FILL
XFILL_0__9025_ vdd gnd FILL
XFILL_0__11739_ vdd gnd FILL
X_9653_ _9653_/A _9653_/B _9653_/C _9653_/Y vdd gnd OAI21X1
XFILL_2__13279_ vdd gnd FILL
XFILL_0__14458_ vdd gnd FILL
X_8604_ _8604_/A _8604_/B _8604_/C _8604_/Y vdd gnd AOI21X1
X_9584_ _9584_/A _9584_/B _9584_/Y vdd gnd NAND2X1
XFILL_0__13409_ vdd gnd FILL
XFILL_0__14389_ vdd gnd FILL
X_8535_ _8535_/A _8535_/B _8535_/Y vdd gnd NAND2X1
XCLKBUF1_insert80 CLKBUF1_insert80/A CLKBUF1_insert80/Y vdd gnd CLKBUF1
XCLKBUF1_insert91 CLKBUF1_insert91/A CLKBUF1_insert91/Y vdd gnd CLKBUF1
XFILL_0__9927_ vdd gnd FILL
XFILL_1__8720_ vdd gnd FILL
X_8466_ _8466_/A _8466_/B _8466_/C _8466_/Y vdd gnd NAND3X1
X_7417_ _7417_/A _7417_/B _7417_/C _7417_/D _7417_/Y vdd gnd AOI22X1
XFILL_1__8651_ vdd gnd FILL
XFILL_0__9858_ vdd gnd FILL
X_8397_ _8397_/A _8397_/B _8397_/C _8397_/Y vdd gnd NAND3X1
XFILL_1__7602_ vdd gnd FILL
XFILL_0__8809_ vdd gnd FILL
X_7348_ _7348_/A _7348_/Y vdd gnd INVX1
XFILL_1__8582_ vdd gnd FILL
XFILL256650x126150 vdd gnd FILL
XFILL_1__7533_ vdd gnd FILL
X_7279_ _7279_/A _7279_/B _7279_/C _7279_/Y vdd gnd OAI21X1
X_9018_ _9018_/A _9018_/Y vdd gnd INVX1
XFILL_1__7464_ vdd gnd FILL
XFILL_1__9203_ vdd gnd FILL
XFILL_1__7395_ vdd gnd FILL
XFILL_1__9134_ vdd gnd FILL
X_11920_ _11920_/A _11920_/Y vdd gnd INVX1
X_11851_ _11851_/A _11851_/Y vdd gnd INVX1
XFILL_1__9065_ vdd gnd FILL
X_10802_ _10802_/A _10802_/B _10802_/C _10802_/Y vdd gnd OAI21X1
X_14570_ _14570_/A _14570_/B _14570_/C _14570_/Y vdd gnd OAI21X1
XFILL_1__8016_ vdd gnd FILL
X_11782_ _11782_/A _11782_/B _11782_/S _11782_/Y vdd gnd MUX2X1
X_10733_ _10733_/D _10733_/CLK _10733_/Q vdd gnd DFFPOSX1
X_13521_ _13521_/A _13521_/B _13521_/C _13521_/Y vdd gnd AOI21X1
XFILL256650x3750 vdd gnd FILL
X_13452_ _13452_/D _13452_/CLK _13452_/Q vdd gnd DFFPOSX1
X_10664_ _10664_/A _10664_/B _10664_/Y vdd gnd NAND2X1
XFILL_1__9967_ vdd gnd FILL
XFILL_2__8760_ vdd gnd FILL
X_12403_ _12403_/A _12403_/Y vdd gnd INVX1
X_13383_ _13383_/A _13383_/Y vdd gnd INVX1
X_10595_ _10595_/A _10595_/B _10595_/Y vdd gnd NAND2X1
XFILL_2__8691_ vdd gnd FILL
XFILL_1__9898_ vdd gnd FILL
X_12334_ _12334_/A _12334_/B _12334_/Y vdd gnd OR2X2
XFILL_0__10070_ vdd gnd FILL
X_12265_ _12265_/A _12265_/B _12265_/Y vdd gnd NAND2X1
XFILL_1__11360_ vdd gnd FILL
X_14004_ _14004_/A _14004_/B _14004_/Y vdd gnd AND2X2
X_11216_ _11216_/A _11216_/B _11216_/C _11216_/Y vdd gnd OAI21X1
XFILL_2__9312_ vdd gnd FILL
X_12196_ _12196_/A _12196_/B _12196_/C _12196_/Y vdd gnd OAI21X1
XFILL_1__10311_ vdd gnd FILL
XFILL_2__12650_ vdd gnd FILL
XFILL_1__11291_ vdd gnd FILL
X_11147_ _11147_/A _11147_/B _11147_/Y vdd gnd NAND2X1
XFILL_2__11601_ vdd gnd FILL
XFILL_2__9243_ vdd gnd FILL
XFILL_1__13030_ vdd gnd FILL
XFILL_1__10242_ vdd gnd FILL
XFILL_0__13760_ vdd gnd FILL
XFILL_0__10972_ vdd gnd FILL
X_11078_ _11078_/A _11078_/B _11078_/C _11078_/Y vdd gnd NAND3X1
XFILL_2__14320_ vdd gnd FILL
XFILL_2__9174_ vdd gnd FILL
XFILL_2__11532_ vdd gnd FILL
XFILL_0__12711_ vdd gnd FILL
XFILL_1__10173_ vdd gnd FILL
X_14906_ _14906_/D _14906_/CLK _14906_/Q vdd gnd DFFPOSX1
X_10029_ _10029_/A _10029_/B _10029_/C _10029_/Y vdd gnd AOI21X1
XFILL_0__13691_ vdd gnd FILL
XFILL_2__14251_ vdd gnd FILL
XFILL_2__11463_ vdd gnd FILL
XFILL_0__12642_ vdd gnd FILL
XFILL_0__7140_ vdd gnd FILL
X_14837_ _14837_/A _14837_/B _14837_/Y vdd gnd OR2X2
XFILL_1__13932_ vdd gnd FILL
XFILL_2__11394_ vdd gnd FILL
X_14768_ _14768_/A _14768_/B _14768_/C _14768_/Y vdd gnd OAI21X1
XFILL_0__14312_ vdd gnd FILL
XFILL_1__13863_ vdd gnd FILL
XFILL_0__11524_ vdd gnd FILL
X_13719_ _13719_/A _13719_/B _13719_/C _13719_/Y vdd gnd NAND3X1
X_14699_ _14699_/A _14699_/B _14699_/C _14699_/Y vdd gnd AOI21X1
XFILL_1__12814_ vdd gnd FILL
XFILL_0__14243_ vdd gnd FILL
XFILL_0__11455_ vdd gnd FILL
XFILL_1__13794_ vdd gnd FILL
XFILL_2__12015_ vdd gnd FILL
XFILL_0_BUFX2_insert250 vdd gnd FILL
XFILL_0__10406_ vdd gnd FILL
XFILL_1__12745_ vdd gnd FILL
XFILL_0_BUFX2_insert261 vdd gnd FILL
X_8320_ _8320_/A _8320_/Y vdd gnd INVX1
XFILL_0__11386_ vdd gnd FILL
XFILL_0_BUFX2_insert272 vdd gnd FILL
XFILL_0_BUFX2_insert283 vdd gnd FILL
XFILL_0__13125_ vdd gnd FILL
XFILL_0_BUFX2_insert294 vdd gnd FILL
XFILL_0__10337_ vdd gnd FILL
XFILL_1__12676_ vdd gnd FILL
XFILL_0__9712_ vdd gnd FILL
X_8251_ _8251_/A _8251_/B _8251_/C _8251_/Y vdd gnd AOI21X1
XFILL_1__14415_ vdd gnd FILL
XFILL_0__13056_ vdd gnd FILL
XFILL_2__13966_ vdd gnd FILL
XFILL_0__10268_ vdd gnd FILL
X_7202_ _7202_/A _7202_/B _7202_/C _7202_/Y vdd gnd AOI21X1
XFILL_0__9643_ vdd gnd FILL
XFILL_2_BUFX2_insert10 vdd gnd FILL
X_8182_ _8182_/A _8182_/Y vdd gnd INVX1
XFILL_0__12007_ vdd gnd FILL
XFILL_1__14346_ vdd gnd FILL
XFILL_2__12917_ vdd gnd FILL
XFILL_1__11558_ vdd gnd FILL
XFILL_0__10199_ vdd gnd FILL
X_7133_ _7133_/A _7133_/Y vdd gnd INVX8
XFILL_0__9574_ vdd gnd FILL
XFILL_1__10509_ vdd gnd FILL
XFILL_1__14277_ vdd gnd FILL
XFILL_2__12848_ vdd gnd FILL
XFILL_1__11489_ vdd gnd FILL
XFILL_0__8525_ vdd gnd FILL
XFILL_1__13228_ vdd gnd FILL
XFILL_2__12779_ vdd gnd FILL
XFILL_0__13958_ vdd gnd FILL
XFILL_0__8456_ vdd gnd FILL
XFILL_1__13159_ vdd gnd FILL
XFILL_0__12909_ vdd gnd FILL
XFILL_0__7407_ vdd gnd FILL
XFILL_0__13889_ vdd gnd FILL
XFILL_1__7180_ vdd gnd FILL
XFILL_0__8387_ vdd gnd FILL
XFILL_2__14449_ vdd gnd FILL
XFILL_0__7338_ vdd gnd FILL
X_7966_ _7966_/D _7966_/CLK _7966_/Q vdd gnd DFFPOSX1
X_9705_ _9705_/A _9705_/B _9705_/C _9705_/Y vdd gnd OAI21X1
XFILL_0__7269_ vdd gnd FILL
X_7897_ _7897_/A _7897_/Y vdd gnd INVX1
XFILL_0__9008_ vdd gnd FILL
X_9636_ _9636_/A _9636_/Y vdd gnd INVX1
X_9567_ _9567_/A _9567_/B _9567_/Y vdd gnd NAND2X1
X_8518_ _8518_/A _8518_/B _8518_/C _8518_/Y vdd gnd OAI21X1
XFILL_1__9752_ vdd gnd FILL
X_9498_ _9498_/A _9498_/B _9498_/Y vdd gnd NAND2X1
X_10380_ _10380_/A _10380_/B _10380_/Y vdd gnd NAND2X1
XFILL_1__8703_ vdd gnd FILL
X_8449_ _8449_/A _8449_/B _8449_/Y vdd gnd OR2X2
XFILL_1__9683_ vdd gnd FILL
XFILL_1__8634_ vdd gnd FILL
X_12050_ _12050_/A _12050_/B _12050_/C _12050_/Y vdd gnd AOI21X1
XFILL_1__8565_ vdd gnd FILL
X_11001_ _11001_/A _11001_/B _11001_/C _11001_/Y vdd gnd NAND3X1
XFILL_1__7516_ vdd gnd FILL
XFILL_1__8496_ vdd gnd FILL
XFILL_0_CLKBUF1_insert38 vdd gnd FILL
XFILL_1__7447_ vdd gnd FILL
XFILL_0_CLKBUF1_insert49 vdd gnd FILL
XFILL_2_BUFX2_insert301 vdd gnd FILL
X_12952_ _12952_/A _12952_/B _12952_/C _12952_/Y vdd gnd OAI21X1
XFILL_2_BUFX2_insert334 vdd gnd FILL
XFILL_1__7378_ vdd gnd FILL
XFILL_2_BUFX2_insert356 vdd gnd FILL
X_11903_ _11903_/A _11903_/Y vdd gnd INVX1
XFILL_1__9117_ vdd gnd FILL
X_12883_ _12883_/A _12883_/B _12883_/C _12883_/Y vdd gnd OAI21X1
X_14622_ _14622_/A _14622_/B _14622_/Y vdd gnd NOR2X1
XFILL_1__9048_ vdd gnd FILL
X_11834_ _11834_/A _11834_/B _11834_/C _11834_/Y vdd gnd AOI21X1
X_11765_ _11765_/A _11765_/B _11765_/Y vdd gnd NAND2X1
X_14553_ _14553_/D _14553_/CLK _14553_/Q vdd gnd DFFPOSX1
XBUFX2_insert300 BUFX2_insert300/A BUFX2_insert300/Y vdd gnd BUFX2
XBUFX2_insert311 BUFX2_insert311/A BUFX2_insert311/Y vdd gnd BUFX2
XFILL_1__10860_ vdd gnd FILL
XBUFX2_insert322 BUFX2_insert322/A BUFX2_insert322/Y vdd gnd BUFX2
X_10716_ _10716_/D _10716_/CLK _10716_/Q vdd gnd DFFPOSX1
X_13504_ _13504_/A _13504_/Y vdd gnd INVX2
XBUFX2_insert333 BUFX2_insert333/A BUFX2_insert333/Y vdd gnd BUFX2
XBUFX2_insert344 BUFX2_insert344/A BUFX2_insert344/Y vdd gnd BUFX2
X_14484_ _14484_/A _14484_/B _14484_/Y vdd gnd NAND2X1
X_11696_ _11696_/A _11696_/B _11696_/Y vdd gnd NOR2X1
XBUFX2_insert355 BUFX2_insert355/A BUFX2_insert355/Y vdd gnd BUFX2
XFILL_0__11240_ vdd gnd FILL
XFILL_1__10791_ vdd gnd FILL
XBUFX2_insert366 BUFX2_insert366/A BUFX2_insert366/Y vdd gnd BUFX2
X_10647_ _10647_/A _10647_/B _10647_/C _10647_/Y vdd gnd OAI21X1
XBUFX2_insert377 BUFX2_insert377/A BUFX2_insert377/Y vdd gnd BUFX2
X_13435_ _13435_/D _13435_/CLK _13435_/Q vdd gnd DFFPOSX1
XFILL_1__12530_ vdd gnd FILL
XFILL_0__11171_ vdd gnd FILL
X_13366_ _13366_/A _13366_/B _13366_/Y vdd gnd NAND2X1
X_10578_ _10578_/A _10578_/B _10578_/Y vdd gnd NOR2X1
XFILL_0__10122_ vdd gnd FILL
XFILL_2__13820_ vdd gnd FILL
XFILL_1__12461_ vdd gnd FILL
X_12317_ _12317_/A _12317_/B _12317_/Y vdd gnd NOR2X1
X_13297_ _13297_/A _13297_/B _13297_/Y vdd gnd NAND2X1
XFILL_2__7625_ vdd gnd FILL
XFILL_1__11412_ vdd gnd FILL
XFILL_0__10053_ vdd gnd FILL
XFILL_2__13751_ vdd gnd FILL
XFILL_1__12392_ vdd gnd FILL
X_12248_ _12248_/A _12248_/B _12248_/C _12248_/Y vdd gnd OAI21X1
XFILL_2__12702_ vdd gnd FILL
XFILL_1__14131_ vdd gnd FILL
XFILL_1__11343_ vdd gnd FILL
XFILL_2__13682_ vdd gnd FILL
XFILL_0__14861_ vdd gnd FILL
X_12179_ _12179_/A _12179_/B _12179_/C _12179_/Y vdd gnd NAND3X1
XFILL_2__12633_ vdd gnd FILL
XFILL_1__14062_ vdd gnd FILL
XFILL_0__13812_ vdd gnd FILL
XFILL_0__8310_ vdd gnd FILL
XFILL_1__11274_ vdd gnd FILL
XFILL_0__14792_ vdd gnd FILL
XFILL_0__9290_ vdd gnd FILL
XFILL_2__9226_ vdd gnd FILL
XFILL_1__13013_ vdd gnd FILL
XFILL_1__10225_ vdd gnd FILL
XFILL_0__13743_ vdd gnd FILL
XFILL_0__8241_ vdd gnd FILL
XFILL_0__10955_ vdd gnd FILL
XFILL_2__11515_ vdd gnd FILL
XFILL_2__9157_ vdd gnd FILL
XFILL_1__10156_ vdd gnd FILL
XFILL_0__13674_ vdd gnd FILL
X_7820_ _7820_/A _7820_/Y vdd gnd INVX1
XFILL_0__8172_ vdd gnd FILL
XFILL_0__10886_ vdd gnd FILL
XFILL_2__9088_ vdd gnd FILL
XFILL_2__11446_ vdd gnd FILL
XFILL_0__12625_ vdd gnd FILL
XFILL_0__7123_ vdd gnd FILL
XFILL_1__10087_ vdd gnd FILL
X_7751_ _7751_/A _7751_/B _7751_/C _7751_/Y vdd gnd OAI21X1
XFILL_1__13915_ vdd gnd FILL
XFILL_2__11377_ vdd gnd FILL
X_7682_ _7682_/A _7682_/B _7682_/Y vdd gnd AND2X2
XFILL_0__11507_ vdd gnd FILL
XFILL_1__13846_ vdd gnd FILL
X_9421_ _9421_/A _9421_/B _9421_/C _9421_/Y vdd gnd NAND3X1
XFILL_0__12487_ vdd gnd FILL
XFILL_0__14226_ vdd gnd FILL
XFILL_0__11438_ vdd gnd FILL
XFILL_1__13777_ vdd gnd FILL
XFILL_1__10989_ vdd gnd FILL
X_9352_ _9352_/A _9352_/B _9352_/Y vdd gnd AND2X2
XFILL_1__12728_ vdd gnd FILL
XFILL_0__14157_ vdd gnd FILL
X_8303_ _8303_/A _8303_/B _8303_/C _8303_/Y vdd gnd NOR3X1
XFILL_0__11369_ vdd gnd FILL
X_9283_ _9283_/A _9283_/Y vdd gnd INVX1
XFILL_0__13108_ vdd gnd FILL
XFILL_1__12659_ vdd gnd FILL
XFILL_0__14088_ vdd gnd FILL
X_8234_ _8234_/A _8234_/B _8234_/C _8234_/Y vdd gnd NAND3X1
XFILL_0__7887_ vdd gnd FILL
XFILL_2__13949_ vdd gnd FILL
XFILL_0__13039_ vdd gnd FILL
XFILL_0__9626_ vdd gnd FILL
X_8165_ _8165_/A _8165_/B _8165_/C _8165_/Y vdd gnd OAI21X1
XFILL_1__14329_ vdd gnd FILL
X_7116_ _7116_/A _7116_/B _7116_/C _7116_/Y vdd gnd AOI21X1
XFILL_1__8350_ vdd gnd FILL
XFILL_0__9557_ vdd gnd FILL
X_8096_ _8096_/A _8096_/Y vdd gnd INVX1
XFILL_1__7301_ vdd gnd FILL
XFILL_0__8508_ vdd gnd FILL
XFILL_1__8281_ vdd gnd FILL
XFILL_0__9488_ vdd gnd FILL
XFILL_1__7232_ vdd gnd FILL
XFILL_0__8439_ vdd gnd FILL
XFILL_1__7163_ vdd gnd FILL
X_8998_ _8998_/A _8998_/B _8998_/Y vdd gnd NAND2X1
XFILL_1_BUFX2_insert308 vdd gnd FILL
XFILL_1_BUFX2_insert319 vdd gnd FILL
X_7949_ _7949_/D _7949_/CLK _7949_/Q vdd gnd DFFPOSX1
XFILL_1__7094_ vdd gnd FILL
X_11550_ _11550_/A _11550_/B _11550_/Y vdd gnd NAND2X1
X_9619_ _9619_/A _9619_/B _9619_/C _9619_/Y vdd gnd OAI21X1
X_10501_ _10501_/A _10501_/B _10501_/Y vdd gnd NOR2X1
X_11481_ _11481_/A _11481_/B _11481_/Y vdd gnd OR2X2
X_13220_ _13220_/A _13220_/B _13220_/C _13220_/Y vdd gnd OAI21X1
XFILL_1__7996_ vdd gnd FILL
X_10432_ _10432_/A _10432_/B _10432_/C _10432_/Y vdd gnd OAI21X1
XFILL_1__9735_ vdd gnd FILL
X_13151_ _13151_/A _13151_/B _13151_/C _13151_/Y vdd gnd OAI21X1
X_10363_ _10363_/A _10363_/B _10363_/Y vdd gnd AND2X2
XFILL_1__9666_ vdd gnd FILL
X_12102_ _12102_/A _12102_/B _12102_/Y vdd gnd OR2X2
X_13082_ _13082_/A _13082_/B _13082_/C _13082_/Y vdd gnd NAND3X1
X_10294_ _10294_/A _10294_/Y vdd gnd INVX1
XFILL_2__7410_ vdd gnd FILL
XFILL_1__8617_ vdd gnd FILL
XFILL_1__9597_ vdd gnd FILL
X_12033_ _12033_/A _12033_/B _12033_/C _12033_/Y vdd gnd NAND3X1
XFILL_2__7341_ vdd gnd FILL
XFILL_1__8548_ vdd gnd FILL
XFILL_2__7272_ vdd gnd FILL
XFILL_1__8479_ vdd gnd FILL
XFILL_2_BUFX2_insert120 vdd gnd FILL
X_13984_ _13984_/A _13984_/B _13984_/C _13984_/Y vdd gnd OAI21X1
XFILL_1__10010_ vdd gnd FILL
XFILL_2_BUFX2_insert153 vdd gnd FILL
X_12935_ _12935_/A _12935_/B _12935_/C _12935_/Y vdd gnd NAND3X1
XFILL_2_BUFX2_insert175 vdd gnd FILL
XFILL_0__10671_ vdd gnd FILL
X_12866_ _12866_/A _12866_/B _12866_/C _12866_/Y vdd gnd NAND3X1
XFILL_0__12410_ vdd gnd FILL
XFILL_1__11961_ vdd gnd FILL
X_14605_ _14605_/A _14605_/B _14605_/C _14605_/Y vdd gnd AOI21X1
XFILL_0__13390_ vdd gnd FILL
X_11817_ _11817_/A _11817_/Y vdd gnd INVX1
XFILL_1__13700_ vdd gnd FILL
X_12797_ _12797_/A _12797_/B _12797_/Y vdd gnd NAND2X1
XFILL_1__10912_ vdd gnd FILL
XFILL_1__14680_ vdd gnd FILL
XFILL_0__12341_ vdd gnd FILL
XFILL_1__11892_ vdd gnd FILL
X_14536_ _14536_/D _14536_/CLK _14536_/Q vdd gnd DFFPOSX1
XFILL_2__10113_ vdd gnd FILL
X_11748_ _11748_/A _11748_/B _11748_/C _11748_/D _11748_/Y vdd gnd AOI22X1
XFILL_1__13631_ vdd gnd FILL
XBUFX2_insert130 BUFX2_insert130/A BUFX2_insert130/Y vdd gnd BUFX2
XBUFX2_insert141 BUFX2_insert141/A BUFX2_insert141/Y vdd gnd BUFX2
XFILL_1__10843_ vdd gnd FILL
XFILL_0__12272_ vdd gnd FILL
XBUFX2_insert152 BUFX2_insert152/A BUFX2_insert152/Y vdd gnd BUFX2
XBUFX2_insert163 BUFX2_insert163/A BUFX2_insert163/Y vdd gnd BUFX2
X_14467_ _14467_/A _14467_/B _14467_/C _14467_/Y vdd gnd OAI21X1
XFILL_2__10044_ vdd gnd FILL
X_11679_ _11679_/D _11679_/CLK _11679_/Q vdd gnd DFFPOSX1
XFILL_0__14011_ vdd gnd FILL
XBUFX2_insert174 BUFX2_insert174/A BUFX2_insert174/Y vdd gnd BUFX2
XBUFX2_insert185 BUFX2_insert185/A BUFX2_insert185/Y vdd gnd BUFX2
XFILL_0__11223_ vdd gnd FILL
XFILL_1__13562_ vdd gnd FILL
XBUFX2_insert196 BUFX2_insert196/A BUFX2_insert196/Y vdd gnd BUFX2
XFILL_1__10774_ vdd gnd FILL
XFILL_0__7810_ vdd gnd FILL
X_13418_ _13418_/A _13418_/B _13418_/Y vdd gnd NAND2X1
XFILL_0__8790_ vdd gnd FILL
XFILL_1__12513_ vdd gnd FILL
X_14398_ _14398_/A _14398_/B _14398_/Y vdd gnd NOR2X1
XFILL_0__11154_ vdd gnd FILL
XFILL_0__7741_ vdd gnd FILL
X_13349_ _13349_/A _13349_/B _13349_/Y vdd gnd NAND2X1
XFILL_0__10105_ vdd gnd FILL
XFILL_1__12444_ vdd gnd FILL
XFILL_0__11085_ vdd gnd FILL
XFILL_0__7672_ vdd gnd FILL
XFILL_2__7608_ vdd gnd FILL
XFILL_2__13734_ vdd gnd FILL
XFILL_0__10036_ vdd gnd FILL
XFILL_0__14913_ vdd gnd FILL
XFILL_1__12375_ vdd gnd FILL
XFILL_2__10946_ vdd gnd FILL
XFILL_0__9411_ vdd gnd FILL
XFILL_1__14114_ vdd gnd FILL
XFILL_2__7539_ vdd gnd FILL
XFILL_1__11326_ vdd gnd FILL
XFILL_2__13665_ vdd gnd FILL
XFILL_0__14844_ vdd gnd FILL
XFILL_2__10877_ vdd gnd FILL
XFILL_0__9342_ vdd gnd FILL
X_9970_ _9970_/A _9970_/B _9970_/C _9970_/Y vdd gnd NAND3X1
XFILL_1__14045_ vdd gnd FILL
XFILL_1__11257_ vdd gnd FILL
XFILL_0__14775_ vdd gnd FILL
XFILL_2__13596_ vdd gnd FILL
XFILL_0__9273_ vdd gnd FILL
X_8921_ _8921_/A _8921_/Y vdd gnd INVX2
XFILL_0__11987_ vdd gnd FILL
XFILL_1__10208_ vdd gnd FILL
XFILL_0__13726_ vdd gnd FILL
XFILL_0__10938_ vdd gnd FILL
XFILL_0__8224_ vdd gnd FILL
XFILL_1__11188_ vdd gnd FILL
X_8852_ _8852_/D _8852_/CLK _8852_/Q vdd gnd DFFPOSX1
XFILL_1__10139_ vdd gnd FILL
XFILL_0__13657_ vdd gnd FILL
X_7803_ _7803_/A _7803_/B _7803_/C _7803_/Y vdd gnd AOI21X1
XFILL_0__8155_ vdd gnd FILL
XFILL_0__10869_ vdd gnd FILL
X_8783_ _8783_/A _8783_/B _8783_/C _8783_/Y vdd gnd OAI21X1
XFILL_0__7106_ vdd gnd FILL
XFILL_0__13588_ vdd gnd FILL
X_7734_ _7734_/A _7734_/B _7734_/C _7734_/Y vdd gnd AOI21X1
XFILL_0__8086_ vdd gnd FILL
X_7665_ _7665_/A _7665_/B _7665_/Y vdd gnd OR2X2
XFILL_1__13829_ vdd gnd FILL
X_9404_ _9404_/A _9404_/B _9404_/Y vdd gnd NAND2X1
XFILL_1__7850_ vdd gnd FILL
X_7596_ _7596_/A _7596_/B _7596_/C _7596_/Y vdd gnd OAI21X1
X_9335_ _9335_/A _9335_/B _9335_/Y vdd gnd NAND2X1
XFILL_0__8988_ vdd gnd FILL
XFILL_1__7781_ vdd gnd FILL
XFILL_1__9520_ vdd gnd FILL
X_9266_ _9266_/A _9266_/B _9266_/Y vdd gnd NAND2X1
X_8217_ _8217_/A _8217_/Y vdd gnd INVX1
XFILL_1__9451_ vdd gnd FILL
X_9197_ _9197_/A _9197_/B _9197_/C _9197_/Y vdd gnd OAI21X1
XFILL_0__9609_ vdd gnd FILL
XFILL_1__8402_ vdd gnd FILL
X_8148_ _8148_/A _8148_/B _8148_/Y vdd gnd NOR2X1
XFILL_1__9382_ vdd gnd FILL
XFILL_1__8333_ vdd gnd FILL
X_8079_ _8079_/A _8079_/B _8079_/C _8079_/Y vdd gnd OAI21X1
XFILL_1__8264_ vdd gnd FILL
X_10981_ _10981_/A _10981_/B _10981_/Y vdd gnd NAND2X1
XFILL_1__7215_ vdd gnd FILL
XFILL_1__8195_ vdd gnd FILL
X_12720_ _12720_/A _12720_/B _12720_/Y vdd gnd NAND2X1
XFILL_1__7146_ vdd gnd FILL
XFILL_1_BUFX2_insert116 vdd gnd FILL
XFILL_1_BUFX2_insert127 vdd gnd FILL
XFILL_1_BUFX2_insert138 vdd gnd FILL
XFILL_1_BUFX2_insert149 vdd gnd FILL
X_12651_ _12651_/A _12651_/Y vdd gnd INVX1
XFILL_1__7077_ vdd gnd FILL
X_11602_ _11602_/A _11602_/B _11602_/Y vdd gnd NAND2X1
X_12582_ _12582_/D _12582_/CLK _12582_/Q vdd gnd DFFPOSX1
X_14321_ _14321_/A _14321_/B _14321_/Y vdd gnd OR2X2
X_11533_ _11533_/A _11533_/B _11533_/Y vdd gnd NAND2X1
X_14252_ _14252_/A _14252_/Y vdd gnd INVX1
X_11464_ _11464_/A _11464_/B _11464_/C _11464_/Y vdd gnd OAI21X1
XFILL_2__9560_ vdd gnd FILL
X_13203_ _13203_/A _13203_/B _13203_/C _13203_/Y vdd gnd NAND3X1
X_10415_ _10415_/A _10415_/Y vdd gnd INVX1
XFILL_1__9718_ vdd gnd FILL
X_11395_ _11395_/A _11395_/B _11395_/Y vdd gnd AND2X2
X_14183_ _14183_/D _14183_/CLK _14183_/Q vdd gnd DFFPOSX1
XFILL_2__9491_ vdd gnd FILL
XFILL_1__10490_ vdd gnd FILL
X_13134_ _13134_/A _13134_/B _13134_/Y vdd gnd NAND2X1
X_10346_ _10346_/A _10346_/B _10346_/C _10346_/Y vdd gnd AOI21X1
XFILL_1__9649_ vdd gnd FILL
XFILL_2__10800_ vdd gnd FILL
X_13065_ _13065_/A _13065_/B _13065_/C _13065_/D _13065_/Y vdd gnd AOI22X1
X_10277_ _10277_/A _10277_/B _10277_/Y vdd gnd NOR2X1
XFILL_0__11910_ vdd gnd FILL
XFILL_1__12160_ vdd gnd FILL
X_12016_ _12016_/A _12016_/Y vdd gnd INVX1
XFILL_0__12890_ vdd gnd FILL
XFILL_2__7324_ vdd gnd FILL
XFILL_1__11111_ vdd gnd FILL
XFILL_0__11841_ vdd gnd FILL
XFILL_1__12091_ vdd gnd FILL
XFILL_2__12401_ vdd gnd FILL
XFILL_1__11042_ vdd gnd FILL
XFILL_2__7255_ vdd gnd FILL
XFILL_0__14560_ vdd gnd FILL
XFILL_0__11772_ vdd gnd FILL
X_13967_ _13967_/A _13967_/B _13967_/Y vdd gnd NAND2X1
XFILL_2__12332_ vdd gnd FILL
XFILL_2__7186_ vdd gnd FILL
XFILL_0__13511_ vdd gnd FILL
XFILL_0__14491_ vdd gnd FILL
X_12918_ _12918_/A _12918_/B _12918_/C _12918_/Y vdd gnd OAI21X1
XFILL_1__14801_ vdd gnd FILL
XFILL_2__12263_ vdd gnd FILL
X_13898_ _13898_/A _13898_/B _13898_/C _13898_/Y vdd gnd OAI21X1
XFILL_0__10654_ vdd gnd FILL
XFILL_1__12993_ vdd gnd FILL
X_12849_ _12849_/A _12849_/B _12849_/C _12849_/Y vdd gnd NAND3X1
XFILL_1__14732_ vdd gnd FILL
XFILL_1__11944_ vdd gnd FILL
XFILL_0__13373_ vdd gnd FILL
XFILL_0__10585_ vdd gnd FILL
XFILL_0__9960_ vdd gnd FILL
XFILL_0__12324_ vdd gnd FILL
XFILL_1__14663_ vdd gnd FILL
XFILL_1__11875_ vdd gnd FILL
X_14519_ _14519_/D _14519_/CLK _14519_/Q vdd gnd DFFPOSX1
X_7450_ _7450_/A _7450_/B _7450_/Y vdd gnd NOR2X1
XFILL_0__9891_ vdd gnd FILL
XFILL_1__13614_ vdd gnd FILL
XFILL_1__10826_ vdd gnd FILL
XFILL_1__14594_ vdd gnd FILL
XFILL_0__12255_ vdd gnd FILL
X_7381_ _7381_/A _7381_/B _7381_/C _7381_/Y vdd gnd OAI21X1
XFILL_2__10027_ vdd gnd FILL
XFILL_1__13545_ vdd gnd FILL
XFILL_0__11206_ vdd gnd FILL
XFILL_2__9758_ vdd gnd FILL
X_9120_ _9120_/A _9120_/B _9120_/Y vdd gnd NOR2X1
XFILL_0__12186_ vdd gnd FILL
XFILL_0__8773_ vdd gnd FILL
XFILL_2__9689_ vdd gnd FILL
XFILL_0__11137_ vdd gnd FILL
X_9051_ _9051_/A _9051_/B _9051_/C _9051_/Y vdd gnd OAI21X1
XFILL_0__7724_ vdd gnd FILL
XFILL_1__12427_ vdd gnd FILL
XFILL_0__11068_ vdd gnd FILL
X_8002_ _8002_/A _8002_/B _8002_/Y vdd gnd NOR2X1
XFILL_0__7655_ vdd gnd FILL
XFILL_0__10019_ vdd gnd FILL
XFILL_1__12358_ vdd gnd FILL
XFILL_2__10929_ vdd gnd FILL
XFILL_0__7586_ vdd gnd FILL
XFILL_1__11309_ vdd gnd FILL
XFILL_0__14827_ vdd gnd FILL
XFILL_1__12289_ vdd gnd FILL
XFILL_0__9325_ vdd gnd FILL
X_9953_ _9953_/A _9953_/B _9953_/C _9953_/Y vdd gnd OAI21X1
XFILL_1__14028_ vdd gnd FILL
XFILL_0__14758_ vdd gnd FILL
XFILL_0__9256_ vdd gnd FILL
X_8904_ _8904_/D _8904_/CLK _8904_/Q vdd gnd DFFPOSX1
X_9884_ _9884_/A _9884_/B _9884_/C _9884_/D _9884_/Y vdd gnd AOI22X1
XFILL_0__13709_ vdd gnd FILL
XFILL_0__14689_ vdd gnd FILL
XFILL_0__8207_ vdd gnd FILL
XFILL_0__9187_ vdd gnd FILL
X_8835_ _8835_/A _8835_/B _8835_/C _8835_/Y vdd gnd OAI21X1
XFILL_0__8138_ vdd gnd FILL
X_8766_ _8766_/A _8766_/B _8766_/C _8766_/Y vdd gnd OAI21X1
X_7717_ _7717_/A _7717_/B _7717_/Y vdd gnd NOR2X1
XFILL_0__8069_ vdd gnd FILL
XFILL_1__8951_ vdd gnd FILL
X_8697_ _8697_/A _8697_/B _8697_/Y vdd gnd NAND2X1
XFILL_1__7902_ vdd gnd FILL
X_7648_ _7648_/A _7648_/B _7648_/Y vdd gnd NAND2X1
XFILL_1__7833_ vdd gnd FILL
X_7579_ _7579_/A _7579_/Y vdd gnd INVX1
X_9318_ _9318_/A _9318_/B _9318_/Y vdd gnd NAND2X1
XFILL_1__7764_ vdd gnd FILL
X_10200_ _10200_/A _10200_/Y vdd gnd INVX1
XFILL_1__9503_ vdd gnd FILL
X_11180_ _11180_/A _11180_/B _11180_/C _11180_/Y vdd gnd OAI21X1
X_9249_ _9249_/A _9249_/B _9249_/C _9249_/Y vdd gnd OAI21X1
XFILL_1__7695_ vdd gnd FILL
X_10131_ _10131_/A _10131_/B _10131_/Y vdd gnd NOR2X1
XFILL_1__9434_ vdd gnd FILL
X_10062_ _10062_/A _10062_/B _10062_/C _10062_/Y vdd gnd OAI21X1
XFILL_1__9365_ vdd gnd FILL
X_14870_ _14870_/D _14870_/CLK _14870_/Q vdd gnd DFFPOSX1
XFILL_1__8316_ vdd gnd FILL
XFILL_1__9296_ vdd gnd FILL
X_13821_ _13821_/A _13821_/B _13821_/Y vdd gnd NAND2X1
XFILL_1__8247_ vdd gnd FILL
X_13752_ _13752_/A _13752_/B _13752_/C _13752_/Y vdd gnd NAND3X1
X_10964_ _10964_/A _10964_/B _10964_/Y vdd gnd OR2X2
XFILL_1__8178_ vdd gnd FILL
X_12703_ _12703_/A _12703_/B _12703_/C _12703_/Y vdd gnd NAND3X1
XFILL_1__7129_ vdd gnd FILL
X_13683_ _13683_/A _13683_/B _13683_/Y vdd gnd NOR2X1
X_10895_ _10895_/A _10895_/B _10895_/Y vdd gnd AND2X2
X_12634_ _12634_/A _12634_/B _12634_/C _12634_/Y vdd gnd OAI21X1
XFILL_0__10370_ vdd gnd FILL
XFILL_1_CLKBUF1_insert90 vdd gnd FILL
X_12565_ _12565_/D _12565_/CLK _12565_/Q vdd gnd DFFPOSX1
X_14304_ _14304_/A _14304_/Y vdd gnd INVX1
X_11516_ _11516_/A _11516_/Y vdd gnd INVX1
XFILL_2__9612_ vdd gnd FILL
XFILL_1__10611_ vdd gnd FILL
X_12496_ _12496_/A _12496_/B _12496_/Y vdd gnd NAND2X1
XFILL_2__12950_ vdd gnd FILL
XFILL_0__12040_ vdd gnd FILL
XFILL_1__11591_ vdd gnd FILL
X_14235_ _14235_/A _14235_/B _14235_/Y vdd gnd NAND2X1
X_11447_ _11447_/A _11447_/B _11447_/C _11447_/Y vdd gnd OAI21X1
XFILL_2__9543_ vdd gnd FILL
XFILL_1__13330_ vdd gnd FILL
XFILL_1__10542_ vdd gnd FILL
XFILL_2__12881_ vdd gnd FILL
X_14166_ _14166_/D _14166_/CLK _14166_/Q vdd gnd DFFPOSX1
X_11378_ _11378_/A _11378_/B _11378_/Y vdd gnd AND2X2
XFILL_2__14620_ vdd gnd FILL
XFILL_2__9474_ vdd gnd FILL
XFILL_1__13261_ vdd gnd FILL
XFILL_1__10473_ vdd gnd FILL
X_13117_ _13117_/A _13117_/B _13117_/C _13117_/Y vdd gnd OAI21X1
X_10329_ _10329_/A _10329_/B _10329_/C _10329_/Y vdd gnd OAI21X1
XFILL_0__13991_ vdd gnd FILL
XFILL_1__12212_ vdd gnd FILL
X_14097_ _14097_/A _14097_/B _14097_/C _14097_/Y vdd gnd OAI21X1
XFILL_1__13192_ vdd gnd FILL
XFILL_0__12942_ vdd gnd FILL
XFILL_0__7440_ vdd gnd FILL
X_13048_ _13048_/A _13048_/B _13048_/C _13048_/Y vdd gnd OAI21X1
XFILL_1__12143_ vdd gnd FILL
XFILL_0__12873_ vdd gnd FILL
XFILL_0__7371_ vdd gnd FILL
XFILL_0__14612_ vdd gnd FILL
XFILL_1__12074_ vdd gnd FILL
XFILL_0__11824_ vdd gnd FILL
XFILL_0__9110_ vdd gnd FILL
XFILL_1__11025_ vdd gnd FILL
XFILL_0__11755_ vdd gnd FILL
XFILL_0__9041_ vdd gnd FILL
XFILL_2__12315_ vdd gnd FILL
XFILL_2__7169_ vdd gnd FILL
XFILL256950x86550 vdd gnd FILL
XFILL_0__14474_ vdd gnd FILL
X_8620_ _8620_/A _8620_/B _8620_/C _8620_/Y vdd gnd AOI21X1
XFILL_2__12246_ vdd gnd FILL
XFILL_0__13425_ vdd gnd FILL
XFILL_0__10637_ vdd gnd FILL
XFILL_1__12976_ vdd gnd FILL
X_8551_ _8551_/A _8551_/B _8551_/C _8551_/Y vdd gnd NAND3X1
XFILL_1__14715_ vdd gnd FILL
XFILL_2__12177_ vdd gnd FILL
XFILL_1__11927_ vdd gnd FILL
XFILL_0__13356_ vdd gnd FILL
X_7502_ _7502_/A _7502_/B _7502_/C _7502_/Y vdd gnd AOI21X1
XFILL_0__10568_ vdd gnd FILL
XFILL_0__9943_ vdd gnd FILL
X_8482_ _8482_/A _8482_/Y vdd gnd INVX1
XFILL_0__12307_ vdd gnd FILL
XFILL_1__14646_ vdd gnd FILL
XFILL_1__11858_ vdd gnd FILL
XFILL_0__13287_ vdd gnd FILL
X_7433_ _7433_/A _7433_/B _7433_/Y vdd gnd NAND2X1
XFILL_0__10499_ vdd gnd FILL
XFILL_0__9874_ vdd gnd FILL
XFILL_0__12238_ vdd gnd FILL
XFILL_1__10809_ vdd gnd FILL
XFILL_1__14577_ vdd gnd FILL
XFILL_1__11789_ vdd gnd FILL
XFILL_0__8825_ vdd gnd FILL
X_7364_ _7364_/A _7364_/B _7364_/C _7364_/Y vdd gnd OAI21X1
XFILL_1__13528_ vdd gnd FILL
X_9103_ _9103_/A _9103_/B _9103_/C _9103_/Y vdd gnd OAI21X1
XFILL_0__12169_ vdd gnd FILL
XFILL_0__8756_ vdd gnd FILL
X_7295_ _7295_/A _7295_/B _7295_/Y vdd gnd AND2X2
X_9034_ _9034_/A _9034_/B _9034_/S _9034_/Y vdd gnd MUX2X1
XFILL_0__7707_ vdd gnd FILL
XFILL_1__7480_ vdd gnd FILL
XFILL_0__8687_ vdd gnd FILL
XFILL_0__7638_ vdd gnd FILL
XFILL_1__9150_ vdd gnd FILL
XFILL_0__7569_ vdd gnd FILL
XFILL_0__9308_ vdd gnd FILL
XFILL_1__8101_ vdd gnd FILL
XFILL_1__9081_ vdd gnd FILL
X_9936_ _9936_/A _9936_/B _9936_/Y vdd gnd NAND2X1
XFILL_0__9239_ vdd gnd FILL
XFILL_1__8032_ vdd gnd FILL
X_9867_ _9867_/A _9867_/B _9867_/Y vdd gnd NAND2X1
X_8818_ _8818_/A _8818_/Y vdd gnd INVX1
X_9798_ _9798_/D _9798_/CLK _9798_/Q vdd gnd DFFPOSX1
X_10680_ _10680_/A _10680_/B _10680_/C _10680_/Y vdd gnd OAI21X1
XFILL_1__9983_ vdd gnd FILL
X_8749_ _8749_/A _8749_/B _8749_/Y vdd gnd NAND2X1
XFILL_1__8934_ vdd gnd FILL
X_12350_ _12350_/A _12350_/B _12350_/Y vdd gnd NAND2X1
XFILL_1_CLKBUF1_insert101 vdd gnd FILL
X_11301_ _11301_/A _11301_/B _11301_/C _11301_/Y vdd gnd NAND3X1
X_12281_ _12281_/A _12281_/Y vdd gnd INVX1
XFILL_1__7816_ vdd gnd FILL
XFILL_1__8796_ vdd gnd FILL
X_11232_ _11232_/A _11232_/Y vdd gnd INVX1
X_14020_ _14020_/A _14020_/Y vdd gnd INVX1
XFILL_1__7747_ vdd gnd FILL
X_11163_ _11163_/A _11163_/Y vdd gnd INVX1
XFILL_1__7678_ vdd gnd FILL
X_10114_ _10114_/A _10114_/B _10114_/Y vdd gnd NAND2X1
X_11094_ _11094_/A _11094_/B _11094_/C _11094_/Y vdd gnd NAND3X1
XFILL_1__9417_ vdd gnd FILL
XFILL_2__8210_ vdd gnd FILL
X_10045_ _10045_/A _10045_/B _10045_/Y vdd gnd AND2X2
XFILL_1__9348_ vdd gnd FILL
XFILL_2__8141_ vdd gnd FILL
X_14853_ _14853_/A _14853_/B _14853_/C _14853_/Y vdd gnd AOI21X1
XFILL_2__10430_ vdd gnd FILL
XFILL_1__9279_ vdd gnd FILL
XFILL_2__8072_ vdd gnd FILL
X_13804_ _13804_/A _13804_/B _13804_/Y vdd gnd AND2X2
X_14784_ _14784_/A _14784_/B _14784_/Y vdd gnd OR2X2
XFILL_2__10361_ vdd gnd FILL
X_11996_ _11996_/A _11996_/Y vdd gnd INVX1
XFILL_0__11540_ vdd gnd FILL
X_13735_ _13735_/A _13735_/Y vdd gnd INVX1
X_10947_ _10947_/A _10947_/B _10947_/C _10947_/Y vdd gnd AOI21X1
XFILL_1__12830_ vdd gnd FILL
XFILL_0__11471_ vdd gnd FILL
X_13666_ _13666_/A _13666_/Y vdd gnd INVX1
XFILL_2__12031_ vdd gnd FILL
XFILL_0__13210_ vdd gnd FILL
XFILL256950x18150 vdd gnd FILL
X_10878_ _10878_/A _10878_/Y vdd gnd INVX1
XFILL_0__10422_ vdd gnd FILL
XFILL_2__8974_ vdd gnd FILL
XFILL_1__12761_ vdd gnd FILL
X_12617_ _12617_/A _12617_/B _12617_/Y vdd gnd NOR2X1
X_13597_ _13597_/A _13597_/B _13597_/Y vdd gnd NAND2X1
XFILL_1__11712_ vdd gnd FILL
XFILL_0__13141_ vdd gnd FILL
XFILL_0__10353_ vdd gnd FILL
XFILL_1__12692_ vdd gnd FILL
X_12548_ _12548_/D _12548_/CLK _12548_/Q vdd gnd DFFPOSX1
XFILL_2__7856_ vdd gnd FILL
XFILL_1__14431_ vdd gnd FILL
XFILL_2__13982_ vdd gnd FILL
XFILL_0__13072_ vdd gnd FILL
XFILL_0__10284_ vdd gnd FILL
X_12479_ _12479_/A _12479_/B _12479_/C _12479_/Y vdd gnd OAI21X1
XFILL_1__14362_ vdd gnd FILL
XFILL_0__12023_ vdd gnd FILL
XFILL_2__7787_ vdd gnd FILL
XFILL_1__11574_ vdd gnd FILL
X_14218_ _14218_/A _14218_/B _14218_/C _14218_/Y vdd gnd OAI21X1
XFILL_0__8610_ vdd gnd FILL
XFILL_0__9590_ vdd gnd FILL
XFILL_1__13313_ vdd gnd FILL
XFILL_1__10525_ vdd gnd FILL
XFILL_1__14293_ vdd gnd FILL
XFILL_2__12864_ vdd gnd FILL
XCLKBUF1_insert100 CLKBUF1_insert100/A CLKBUF1_insert100/Y vdd gnd CLKBUF1
XFILL_0__8541_ vdd gnd FILL
X_14149_ _14149_/A _14149_/B _14149_/C _14149_/Y vdd gnd OAI21X1
XFILL_2__14603_ vdd gnd FILL
X_7080_ _7080_/A _7080_/Y vdd gnd INVX2
XFILL_2__11815_ vdd gnd FILL
XFILL_1__13244_ vdd gnd FILL
XFILL_1__10456_ vdd gnd FILL
XFILL_0__13974_ vdd gnd FILL
XFILL_2__12795_ vdd gnd FILL
XFILL_2__8408_ vdd gnd FILL
XFILL_0__8472_ vdd gnd FILL
XFILL_1__13175_ vdd gnd FILL
XFILL_2__9388_ vdd gnd FILL
XFILL_0__12925_ vdd gnd FILL
XFILL_1__10387_ vdd gnd FILL
XFILL_0__7423_ vdd gnd FILL
XFILL_1__12126_ vdd gnd FILL
XFILL_0__12856_ vdd gnd FILL
XFILL_0__7354_ vdd gnd FILL
X_7982_ _7982_/D _7982_/CLK _7982_/Q vdd gnd DFFPOSX1
XFILL_1__12057_ vdd gnd FILL
XFILL_0__11807_ vdd gnd FILL
XFILL_0__12787_ vdd gnd FILL
XFILL_0__7285_ vdd gnd FILL
X_9721_ _9721_/A _9721_/B _9721_/C _9721_/Y vdd gnd OAI21X1
XFILL_1__11008_ vdd gnd FILL
XFILL_0__11738_ vdd gnd FILL
XFILL_0__9024_ vdd gnd FILL
X_9652_ _9652_/A _9652_/B _9652_/C _9652_/Y vdd gnd NAND3X1
XFILL_0__14457_ vdd gnd FILL
X_8603_ _8603_/A _8603_/B _8603_/Y vdd gnd NOR2X1
X_9583_ _9583_/A _9583_/B _9583_/Y vdd gnd NOR2X1
XFILL_2__12229_ vdd gnd FILL
XFILL_0__13408_ vdd gnd FILL
XFILL_0__14388_ vdd gnd FILL
XFILL_1__12959_ vdd gnd FILL
X_8534_ _8534_/A _8534_/B _8534_/C _8534_/Y vdd gnd NAND3X1
XCLKBUF1_insert70 CLKBUF1_insert70/A CLKBUF1_insert70/Y vdd gnd CLKBUF1
XCLKBUF1_insert81 CLKBUF1_insert81/A CLKBUF1_insert81/Y vdd gnd CLKBUF1
XCLKBUF1_insert92 CLKBUF1_insert92/A CLKBUF1_insert92/Y vdd gnd CLKBUF1
XFILL_0__13339_ vdd gnd FILL
XFILL_0__9926_ vdd gnd FILL
X_8465_ _8465_/A _8465_/B _8465_/C _8465_/Y vdd gnd OAI21X1
XFILL_1__14629_ vdd gnd FILL
X_7416_ _7416_/A _7416_/B _7416_/Y vdd gnd OR2X2
XFILL_0__9857_ vdd gnd FILL
XFILL_1__8650_ vdd gnd FILL
X_8396_ _8396_/A _8396_/B _8396_/C _8396_/Y vdd gnd OAI21X1
XFILL_1__7601_ vdd gnd FILL
XFILL_0__8808_ vdd gnd FILL
X_7347_ _7347_/A _7347_/B _7347_/C _7347_/Y vdd gnd OAI21X1
XFILL_1__8581_ vdd gnd FILL
XFILL_1__7532_ vdd gnd FILL
XFILL_0__8739_ vdd gnd FILL
X_7278_ _7278_/A _7278_/B _7278_/C _7278_/D _7278_/Y vdd gnd AOI22X1
X_9017_ _9017_/A _9017_/B _9017_/C _9017_/D _9017_/Y vdd gnd OAI22X1
XFILL_1__7463_ vdd gnd FILL
XFILL_1__9202_ vdd gnd FILL
XFILL_1__7394_ vdd gnd FILL
XFILL_1__9133_ vdd gnd FILL
X_11850_ _11850_/A _11850_/B _11850_/C _11850_/Y vdd gnd OAI21X1
XFILL_1__9064_ vdd gnd FILL
X_9919_ _9919_/A _9919_/B _9919_/S _9919_/Y vdd gnd MUX2X1
X_10801_ _10801_/A _10801_/Y vdd gnd INVX1
XFILL_1__8015_ vdd gnd FILL
X_11781_ _11781_/A _11781_/B _11781_/S _11781_/Y vdd gnd MUX2X1
X_13520_ _13520_/A _13520_/B _13520_/C _13520_/Y vdd gnd OAI21X1
X_10732_ _10732_/D _10732_/CLK _10732_/Q vdd gnd DFFPOSX1
X_13451_ _13451_/D _13451_/CLK _13451_/Q vdd gnd DFFPOSX1
X_10663_ _10663_/A _10663_/B _10663_/C _10663_/Y vdd gnd OAI21X1
XFILL_1__9966_ vdd gnd FILL
X_12402_ _12402_/A _12402_/B _12402_/Y vdd gnd NAND2X1
XFILL_2__7710_ vdd gnd FILL
X_10594_ _10594_/A _10594_/Y vdd gnd INVX1
X_13382_ _13382_/A _13382_/B _13382_/C _13382_/Y vdd gnd OAI21X1
XFILL_1__9897_ vdd gnd FILL
X_12333_ _12333_/A _12333_/B _12333_/Y vdd gnd NAND2X1
XFILL_2__7641_ vdd gnd FILL
X_12264_ _12264_/A _12264_/B _12264_/C _12264_/Y vdd gnd OAI21X1
XFILL_2__7572_ vdd gnd FILL
XFILL_1__8779_ vdd gnd FILL
X_14003_ _14003_/A _14003_/B _14003_/Y vdd gnd NOR2X1
X_11215_ _11215_/A _11215_/B _11215_/Y vdd gnd OR2X2
X_12195_ _12195_/A _12195_/B _12195_/Y vdd gnd NAND2X1
XFILL_1__10310_ vdd gnd FILL
XFILL_1__11290_ vdd gnd FILL
X_11146_ _11146_/A _11146_/B _11146_/Y vdd gnd NOR2X1
XFILL_1__10241_ vdd gnd FILL
XFILL_0__10971_ vdd gnd FILL
X_11077_ _11077_/A _11077_/B _11077_/C _11077_/Y vdd gnd OAI21X1
XFILL_0__12710_ vdd gnd FILL
XFILL_1__10172_ vdd gnd FILL
X_14905_ _14905_/D _14905_/CLK _14905_/Q vdd gnd DFFPOSX1
X_10028_ _10028_/A _10028_/B _10028_/C _10028_/D _10028_/Y vdd gnd AOI22X1
XFILL_0__13690_ vdd gnd FILL
XFILL_2__8124_ vdd gnd FILL
XFILL_0__12641_ vdd gnd FILL
X_14836_ _14836_/A _14836_/B _14836_/Y vdd gnd NAND2X1
XFILL_2__13201_ vdd gnd FILL
XFILL_2__10413_ vdd gnd FILL
XFILL_2__8055_ vdd gnd FILL
XFILL_1__13931_ vdd gnd FILL
X_14767_ _14767_/A _14767_/B _14767_/Y vdd gnd NAND2X1
XFILL_2__10344_ vdd gnd FILL
X_11979_ _11979_/A _11979_/B _11979_/Y vdd gnd NOR2X1
XFILL_0__14311_ vdd gnd FILL
XFILL_0__11523_ vdd gnd FILL
XFILL_1__13862_ vdd gnd FILL
X_13718_ _13718_/A _13718_/B _13718_/C _13718_/Y vdd gnd OAI21X1
X_14698_ _14698_/A _14698_/B _14698_/C _14698_/Y vdd gnd OAI21X1
XFILL_2__10275_ vdd gnd FILL
XFILL_0__14242_ vdd gnd FILL
XFILL_1__12813_ vdd gnd FILL
XFILL_0__11454_ vdd gnd FILL
XFILL_1__13793_ vdd gnd FILL
X_13649_ _13649_/A _13649_/Y vdd gnd INVX1
XFILL_2__8957_ vdd gnd FILL
XFILL_0__10405_ vdd gnd FILL
XFILL_0_BUFX2_insert240 vdd gnd FILL
XFILL_1__12744_ vdd gnd FILL
XFILL_0__11385_ vdd gnd FILL
XFILL_0_BUFX2_insert251 vdd gnd FILL
XFILL_0_BUFX2_insert262 vdd gnd FILL
XFILL_0_BUFX2_insert273 vdd gnd FILL
XFILL_2__7908_ vdd gnd FILL
XFILL_0__13124_ vdd gnd FILL
XFILL_0__10336_ vdd gnd FILL
XFILL_0_BUFX2_insert284 vdd gnd FILL
XFILL_0__9711_ vdd gnd FILL
XFILL_0_BUFX2_insert295 vdd gnd FILL
XFILL_1__12675_ vdd gnd FILL
X_8250_ _8250_/A _8250_/B _8250_/C _8250_/Y vdd gnd OAI21X1
XFILL_2__7839_ vdd gnd FILL
XFILL_1__14414_ vdd gnd FILL
XFILL_0__13055_ vdd gnd FILL
X_7201_ _7201_/A _7201_/B _7201_/Y vdd gnd OR2X2
XFILL_0__10267_ vdd gnd FILL
XFILL_0__9642_ vdd gnd FILL
X_8181_ _8181_/A _8181_/B _8181_/C _8181_/Y vdd gnd AOI21X1
XFILL_0__12006_ vdd gnd FILL
XFILL_1__14345_ vdd gnd FILL
XFILL_1__11557_ vdd gnd FILL
XFILL_2__13896_ vdd gnd FILL
XFILL_2_BUFX2_insert22 vdd gnd FILL
X_7132_ _7132_/A _7132_/Y vdd gnd INVX8
XFILL_0__10198_ vdd gnd FILL
XFILL_0__9573_ vdd gnd FILL
XFILL_1__10508_ vdd gnd FILL
XFILL_1__14276_ vdd gnd FILL
XFILL_1__11488_ vdd gnd FILL
XFILL_0__8524_ vdd gnd FILL
XFILL_1__10439_ vdd gnd FILL
XFILL_1__13227_ vdd gnd FILL
XFILL_0__13957_ vdd gnd FILL
XFILL_0__8455_ vdd gnd FILL
XFILL_1__13158_ vdd gnd FILL
XFILL_2__11729_ vdd gnd FILL
XFILL_0__12908_ vdd gnd FILL
XFILL_0__7406_ vdd gnd FILL
XFILL257250x3750 vdd gnd FILL
XFILL_0__13888_ vdd gnd FILL
XFILL_1__12109_ vdd gnd FILL
XFILL_0__8386_ vdd gnd FILL
XFILL_1__13089_ vdd gnd FILL
XFILL_0__12839_ vdd gnd FILL
XFILL_0__7337_ vdd gnd FILL
X_7965_ _7965_/D _7965_/CLK _7965_/Q vdd gnd DFFPOSX1
X_9704_ _9704_/A _9704_/B _9704_/C _9704_/Y vdd gnd OAI21X1
XFILL_0__7268_ vdd gnd FILL
X_7896_ _7896_/A _7896_/B _7896_/C _7896_/Y vdd gnd OAI21X1
XFILL_0__9007_ vdd gnd FILL
XFILL_0__7199_ vdd gnd FILL
X_9635_ _9635_/A _9635_/B _9635_/Y vdd gnd NOR2X1
X_9566_ _9566_/A _9566_/B _9566_/Y vdd gnd NAND2X1
XFILL_1__9751_ vdd gnd FILL
X_8517_ _8517_/A _8517_/B _8517_/C _8517_/Y vdd gnd AOI21X1
X_9497_ _9497_/A _9497_/B _9497_/Y vdd gnd NAND2X1
XFILL_0__9909_ vdd gnd FILL
XFILL_1__8702_ vdd gnd FILL
XFILL_1__9682_ vdd gnd FILL
X_8448_ _8448_/A _8448_/B _8448_/Y vdd gnd NAND2X1
XFILL_1__8633_ vdd gnd FILL
X_8379_ _8379_/A _8379_/B _8379_/C _8379_/Y vdd gnd OAI21X1
XFILL_1__8564_ vdd gnd FILL
X_11000_ _11000_/A _11000_/B _11000_/C _11000_/Y vdd gnd OAI21X1
XFILL_1__7515_ vdd gnd FILL
XFILL_1__8495_ vdd gnd FILL
XFILL_0_CLKBUF1_insert39 vdd gnd FILL
XFILL_1__7446_ vdd gnd FILL
XFILL_2_BUFX2_insert313 vdd gnd FILL
X_12951_ _12951_/A _12951_/B _12951_/C _12951_/Y vdd gnd OAI21X1
XFILL_1__7377_ vdd gnd FILL
XFILL_2_BUFX2_insert346 vdd gnd FILL
X_11902_ _11902_/A _11902_/B _11902_/Y vdd gnd NAND2X1
XFILL_1__9116_ vdd gnd FILL
XFILL_2_BUFX2_insert368 vdd gnd FILL
X_12882_ _12882_/A _12882_/B _12882_/C _12882_/Y vdd gnd OAI21X1
X_14621_ _14621_/A _14621_/B _14621_/Y vdd gnd AND2X2
X_11833_ _11833_/A _11833_/B _11833_/C _11833_/D _11833_/Y vdd gnd OAI22X1
XFILL_1__9047_ vdd gnd FILL
X_14552_ _14552_/D _14552_/CLK _14552_/Q vdd gnd DFFPOSX1
X_11764_ _11764_/A _11764_/Y vdd gnd INVX1
XBUFX2_insert301 BUFX2_insert301/A BUFX2_insert301/Y vdd gnd BUFX2
XBUFX2_insert312 BUFX2_insert312/A BUFX2_insert312/Y vdd gnd BUFX2
X_13503_ _13503_/A _13503_/B _13503_/Y vdd gnd NOR2X1
X_10715_ _10715_/D _10715_/CLK _10715_/Q vdd gnd DFFPOSX1
XBUFX2_insert323 BUFX2_insert323/A BUFX2_insert323/Y vdd gnd BUFX2
X_14483_ _14483_/A _14483_/B _14483_/C _14483_/Y vdd gnd OAI21X1
XBUFX2_insert334 BUFX2_insert334/A BUFX2_insert334/Y vdd gnd BUFX2
XFILL_2__10060_ vdd gnd FILL
X_11695_ _11695_/A _11695_/Y vdd gnd INVX2
XBUFX2_insert345 BUFX2_insert345/A BUFX2_insert345/Y vdd gnd BUFX2
XBUFX2_insert356 BUFX2_insert356/A BUFX2_insert356/Y vdd gnd BUFX2
XFILL_1__10790_ vdd gnd FILL
XBUFX2_insert367 BUFX2_insert367/A BUFX2_insert367/Y vdd gnd BUFX2
X_13434_ _13434_/D _13434_/CLK _13434_/Q vdd gnd DFFPOSX1
X_10646_ _10646_/A _10646_/B _10646_/Y vdd gnd NAND2X1
XFILL_1__9949_ vdd gnd FILL
XBUFX2_insert378 BUFX2_insert378/A BUFX2_insert378/Y vdd gnd BUFX2
XFILL_0__11170_ vdd gnd FILL
X_13365_ _13365_/A _13365_/B _13365_/C _13365_/Y vdd gnd OAI21X1
X_10577_ _10577_/A _10577_/B _10577_/C _10577_/Y vdd gnd OAI21X1
XFILL_0__10121_ vdd gnd FILL
XFILL_1__12460_ vdd gnd FILL
X_12316_ _12316_/A _12316_/B _12316_/C _12316_/Y vdd gnd AOI21X1
XFILL_1__11411_ vdd gnd FILL
X_13296_ _13296_/A _13296_/B _13296_/Y vdd gnd NAND2X1
XFILL_2__10962_ vdd gnd FILL
XFILL_0__10052_ vdd gnd FILL
XFILL_1__12391_ vdd gnd FILL
X_12247_ _12247_/A _12247_/B _12247_/C _12247_/Y vdd gnd NAND3X1
XFILL_2__7555_ vdd gnd FILL
XFILL_1__11342_ vdd gnd FILL
XFILL_1__14130_ vdd gnd FILL
XFILL_0__14860_ vdd gnd FILL
XFILL_2__10893_ vdd gnd FILL
X_12178_ _12178_/A _12178_/Y vdd gnd INVX1
XFILL_1__14061_ vdd gnd FILL
XFILL_2__7486_ vdd gnd FILL
XFILL_0__13811_ vdd gnd FILL
XFILL_1__11273_ vdd gnd FILL
XFILL_0__14791_ vdd gnd FILL
X_11129_ _11129_/A _11129_/B _11129_/Y vdd gnd NAND2X1
XFILL_1__13012_ vdd gnd FILL
XFILL_1__10224_ vdd gnd FILL
XFILL_0__13742_ vdd gnd FILL
XFILL_0__10954_ vdd gnd FILL
XFILL_0__8240_ vdd gnd FILL
XFILL_1__10155_ vdd gnd FILL
XFILL_2__12494_ vdd gnd FILL
XFILL_0__13673_ vdd gnd FILL
XFILL_0__10885_ vdd gnd FILL
XFILL_2__8107_ vdd gnd FILL
XFILL_0__8171_ vdd gnd FILL
XFILL_0__12624_ vdd gnd FILL
XFILL_1__10086_ vdd gnd FILL
X_14819_ _14819_/A _14819_/B _14819_/C _14819_/Y vdd gnd OAI21X1
XFILL_0__7122_ vdd gnd FILL
X_7750_ _7750_/A _7750_/B _7750_/C _7750_/Y vdd gnd OAI21X1
XFILL_2__8038_ vdd gnd FILL
XFILL_1__13914_ vdd gnd FILL
XFILL_2__13115_ vdd gnd FILL
X_7681_ _7681_/A _7681_/B _7681_/Y vdd gnd NOR2X1
XFILL_2__10327_ vdd gnd FILL
XFILL_0__11506_ vdd gnd FILL
XFILL_1__13845_ vdd gnd FILL
XFILL_0__12486_ vdd gnd FILL
X_9420_ _9420_/A _9420_/Y vdd gnd INVX1
XFILL_2__10258_ vdd gnd FILL
XFILL_0__14225_ vdd gnd FILL
XFILL_2__13046_ vdd gnd FILL
XFILL_0__11437_ vdd gnd FILL
XFILL_1__13776_ vdd gnd FILL
XFILL_1__10988_ vdd gnd FILL
X_9351_ _9351_/A _9351_/B _9351_/Y vdd gnd NOR2X1
XFILL_2__10189_ vdd gnd FILL
XFILL_1__12727_ vdd gnd FILL
XFILL_0__14156_ vdd gnd FILL
XFILL_0__11368_ vdd gnd FILL
X_8302_ _8302_/A _8302_/Y vdd gnd INVX1
X_9282_ _9282_/A _9282_/B _9282_/Y vdd gnd NAND2X1
XFILL_0__13107_ vdd gnd FILL
XFILL_0__10319_ vdd gnd FILL
XFILL_0__14087_ vdd gnd FILL
XFILL_1__12658_ vdd gnd FILL
XFILL_0__11299_ vdd gnd FILL
X_8233_ _8233_/A _8233_/B _8233_/C _8233_/Y vdd gnd NAND3X1
XFILL_0__7886_ vdd gnd FILL
XFILL_1__11609_ vdd gnd FILL
XFILL_0__13038_ vdd gnd FILL
XFILL_0__9625_ vdd gnd FILL
X_8164_ _8164_/A _8164_/B _8164_/Y vdd gnd NAND2X1
XFILL_1__14328_ vdd gnd FILL
X_7115_ _7115_/A _7115_/B _7115_/C _7115_/Y vdd gnd OAI21X1
XFILL_0__9556_ vdd gnd FILL
X_8095_ _8095_/A _8095_/Y vdd gnd INVX8
XFILL_1__14259_ vdd gnd FILL
XFILL_1__7300_ vdd gnd FILL
XFILL_0__8507_ vdd gnd FILL
XFILL_0__9487_ vdd gnd FILL
XFILL_1__8280_ vdd gnd FILL
XFILL_1__7231_ vdd gnd FILL
XFILL_0__8438_ vdd gnd FILL
XFILL_1__7162_ vdd gnd FILL
XFILL_0__8369_ vdd gnd FILL
X_8997_ _8997_/A _8997_/B _8997_/Y vdd gnd NOR2X1
XFILL_1_BUFX2_insert309 vdd gnd FILL
XFILL_1__7093_ vdd gnd FILL
X_7948_ _7948_/D _7948_/CLK _7948_/Q vdd gnd DFFPOSX1
X_7879_ _7879_/A _7879_/B _7879_/C _7879_/Y vdd gnd OAI21X1
X_9618_ _9618_/A _9618_/B _9618_/Y vdd gnd NAND2X1
X_10500_ _10500_/A _10500_/B _10500_/C _10500_/Y vdd gnd OAI21X1
X_11480_ _11480_/A _11480_/B _11480_/Y vdd gnd NAND2X1
X_9549_ _9549_/A _9549_/B _9549_/Y vdd gnd OR2X2
X_10431_ _10431_/A _10431_/B _10431_/C _10431_/Y vdd gnd OAI21X1
XFILL_1__9734_ vdd gnd FILL
X_13150_ _13150_/A _13150_/B _13150_/Y vdd gnd NAND2X1
X_10362_ _10362_/A _10362_/B _10362_/Y vdd gnd AND2X2
XFILL_1__9665_ vdd gnd FILL
X_12101_ _12101_/A _12101_/B _12101_/Y vdd gnd NAND2X1
X_13081_ _13081_/A _13081_/B _13081_/C _13081_/Y vdd gnd OAI21X1
X_10293_ _10293_/A _10293_/B _10293_/C _10293_/Y vdd gnd AOI21X1
XFILL_1__8616_ vdd gnd FILL
XFILL_1__9596_ vdd gnd FILL
X_12032_ _12032_/A _12032_/B _12032_/Y vdd gnd AND2X2
XFILL_1__8547_ vdd gnd FILL
XFILL_1__8478_ vdd gnd FILL
XFILL257550x68550 vdd gnd FILL
X_13983_ _13983_/A _13983_/B _13983_/Y vdd gnd AND2X2
XFILL_1__7429_ vdd gnd FILL
XFILL_2_BUFX2_insert110 vdd gnd FILL
XFILL_2_BUFX2_insert132 vdd gnd FILL
X_12934_ _12934_/A _12934_/B _12934_/C _12934_/Y vdd gnd AOI21X1
XFILL_2_BUFX2_insert165 vdd gnd FILL
XFILL_2_BUFX2_insert187 vdd gnd FILL
XFILL_0__10670_ vdd gnd FILL
XFILL_2_BUFX2_insert198 vdd gnd FILL
X_12865_ _12865_/A _12865_/Y vdd gnd INVX1
X_14604_ _14604_/A _14604_/B _14604_/C _14604_/Y vdd gnd OAI21X1
XFILL_1__11960_ vdd gnd FILL
X_11816_ _11816_/A _11816_/B _11816_/C _11816_/Y vdd gnd AOI21X1
XFILL_2__9912_ vdd gnd FILL
X_12796_ _12796_/A _12796_/Y vdd gnd INVX1
XFILL_0__12340_ vdd gnd FILL
XFILL_1__10911_ vdd gnd FILL
XFILL_1__11891_ vdd gnd FILL
X_14535_ _14535_/D _14535_/CLK _14535_/Q vdd gnd DFFPOSX1
X_11747_ _11747_/A _11747_/B _11747_/C _11747_/Y vdd gnd OAI21X1
XBUFX2_insert120 BUFX2_insert120/A BUFX2_insert120/Y vdd gnd BUFX2
XFILL_1__13630_ vdd gnd FILL
XBUFX2_insert131 BUFX2_insert131/A BUFX2_insert131/Y vdd gnd BUFX2
XFILL_0__12271_ vdd gnd FILL
XFILL_1__10842_ vdd gnd FILL
XBUFX2_insert142 BUFX2_insert142/A BUFX2_insert142/Y vdd gnd BUFX2
X_14466_ _14466_/A _14466_/B _14466_/C _14466_/Y vdd gnd OAI21X1
XBUFX2_insert153 BUFX2_insert153/A BUFX2_insert153/Y vdd gnd BUFX2
XBUFX2_insert164 BUFX2_insert164/A BUFX2_insert164/Y vdd gnd BUFX2
X_11678_ _11678_/D _11678_/CLK _11678_/Q vdd gnd DFFPOSX1
XFILL_0__14010_ vdd gnd FILL
XBUFX2_insert175 BUFX2_insert175/A BUFX2_insert175/Y vdd gnd BUFX2
XFILL_0__11222_ vdd gnd FILL
XBUFX2_insert186 BUFX2_insert186/A BUFX2_insert186/Y vdd gnd BUFX2
XFILL_1__10773_ vdd gnd FILL
XFILL_1__13561_ vdd gnd FILL
X_13417_ _13417_/A _13417_/B _13417_/C _13417_/Y vdd gnd OAI21X1
XBUFX2_insert197 BUFX2_insert197/A BUFX2_insert197/Y vdd gnd BUFX2
X_10629_ _10629_/A _10629_/B _10629_/C _10629_/Y vdd gnd OAI21X1
X_14397_ _14397_/A _14397_/Y vdd gnd INVX1
XFILL_2__8725_ vdd gnd FILL
XFILL_2__14851_ vdd gnd FILL
XFILL_1__12512_ vdd gnd FILL
XFILL_0__11153_ vdd gnd FILL
XFILL_0__7740_ vdd gnd FILL
X_13348_ _13348_/A _13348_/B _13348_/C _13348_/Y vdd gnd OAI21X1
XFILL_0__10104_ vdd gnd FILL
XFILL_2__14782_ vdd gnd FILL
XFILL_1__12443_ vdd gnd FILL
XFILL_0__11084_ vdd gnd FILL
XFILL_0__7671_ vdd gnd FILL
X_13279_ _13279_/A _13279_/B _13279_/Y vdd gnd OR2X2
XFILL_0__10035_ vdd gnd FILL
XFILL_0__14912_ vdd gnd FILL
XFILL_1__12374_ vdd gnd FILL
XFILL_0__9410_ vdd gnd FILL
XFILL_1__14113_ vdd gnd FILL
XFILL_1__11325_ vdd gnd FILL
XFILL_0__14843_ vdd gnd FILL
XFILL_0__9341_ vdd gnd FILL
XFILL_1__14044_ vdd gnd FILL
XFILL_1__11256_ vdd gnd FILL
XFILL_0__14774_ vdd gnd FILL
XFILL_0__11986_ vdd gnd FILL
XFILL_0__9272_ vdd gnd FILL
X_8920_ _8920_/A _8920_/Y vdd gnd INVX1
XFILL_1__10207_ vdd gnd FILL
XFILL_1__11187_ vdd gnd FILL
XFILL_0__10937_ vdd gnd FILL
XFILL_0__13725_ vdd gnd FILL
XFILL_0__8223_ vdd gnd FILL
X_8851_ _8851_/D _8851_/CLK _8851_/Q vdd gnd DFFPOSX1
XFILL_1__10138_ vdd gnd FILL
XFILL_2__12477_ vdd gnd FILL
XFILL_0__13656_ vdd gnd FILL
XFILL_0__10868_ vdd gnd FILL
X_7802_ _7802_/A _7802_/B _7802_/Y vdd gnd NOR2X1
XFILL_0__8154_ vdd gnd FILL
XFILL_2__14216_ vdd gnd FILL
X_8782_ _8782_/A _8782_/B _8782_/C _8782_/Y vdd gnd OAI21X1
XFILL_1__10069_ vdd gnd FILL
XFILL_0__7105_ vdd gnd FILL
XFILL_0__13587_ vdd gnd FILL
XFILL_0__10799_ vdd gnd FILL
X_7733_ _7733_/A _7733_/B _7733_/C _7733_/Y vdd gnd OAI21X1
XFILL_0__8085_ vdd gnd FILL
XFILL_2__14147_ vdd gnd FILL
X_7664_ _7664_/A _7664_/B _7664_/Y vdd gnd NAND2X1
XFILL_2__14078_ vdd gnd FILL
XFILL_1__13828_ vdd gnd FILL
XFILL_0__12469_ vdd gnd FILL
X_9403_ _9403_/A _9403_/B _9403_/C _9403_/Y vdd gnd AOI21X1
X_7595_ _7595_/A _7595_/B _7595_/Y vdd gnd NOR2X1
XFILL_2__13029_ vdd gnd FILL
XFILL_1__13759_ vdd gnd FILL
X_9334_ _9334_/A _9334_/B _9334_/C _9334_/Y vdd gnd AOI21X1
XFILL_0__8987_ vdd gnd FILL
XFILL_1__7780_ vdd gnd FILL
XFILL_0__14139_ vdd gnd FILL
X_9265_ _9265_/A _9265_/B _9265_/C _9265_/D _9265_/Y vdd gnd AOI22X1
XFILL_1__9450_ vdd gnd FILL
X_8216_ _8216_/A _8216_/B _8216_/C _8216_/Y vdd gnd AOI21X1
XFILL_0__7869_ vdd gnd FILL
X_9196_ _9196_/A _9196_/Y vdd gnd INVX1
XFILL_0__9608_ vdd gnd FILL
XFILL_1__8401_ vdd gnd FILL
XFILL_1__9381_ vdd gnd FILL
X_8147_ _8147_/A _8147_/B _8147_/Y vdd gnd OR2X2
XFILL_0__9539_ vdd gnd FILL
XFILL_1__8332_ vdd gnd FILL
X_8078_ _8078_/A _8078_/Y vdd gnd INVX2
XFILL_1__8263_ vdd gnd FILL
XFILL_1__7214_ vdd gnd FILL
X_10980_ _10980_/A _10980_/B _10980_/C _10980_/Y vdd gnd AOI21X1
XFILL_1__8194_ vdd gnd FILL
XFILL_1__7145_ vdd gnd FILL
XFILL_1_BUFX2_insert117 vdd gnd FILL
XFILL_1_BUFX2_insert128 vdd gnd FILL
XFILL_1_BUFX2_insert139 vdd gnd FILL
X_12650_ _12650_/A _12650_/B _12650_/Y vdd gnd NAND2X1
XFILL_1__7076_ vdd gnd FILL
X_11601_ _11601_/A _11601_/B _11601_/C _11601_/Y vdd gnd OAI21X1
X_12581_ _12581_/D _12581_/CLK _12581_/Q vdd gnd DFFPOSX1
X_14320_ _14320_/A _14320_/B _14320_/C _14320_/Y vdd gnd OAI21X1
X_11532_ _11532_/A _11532_/B _11532_/C _11532_/Y vdd gnd OAI21X1
XFILL257550x43350 vdd gnd FILL
X_14251_ _14251_/A _14251_/B _14251_/C _14251_/Y vdd gnd OAI21X1
X_11463_ _11463_/A _11463_/B _11463_/C _11463_/Y vdd gnd OAI21X1
X_13202_ _13202_/A _13202_/B _13202_/Y vdd gnd OR2X2
X_10414_ _10414_/A _10414_/B _10414_/C _10414_/Y vdd gnd OAI21X1
XFILL_1__9717_ vdd gnd FILL
XFILL_2__8510_ vdd gnd FILL
X_14182_ _14182_/D _14182_/CLK _14182_/Q vdd gnd DFFPOSX1
X_11394_ _11394_/A _11394_/B _11394_/C _11394_/Y vdd gnd OAI21X1
X_13133_ _13133_/A _13133_/B _13133_/C _13133_/Y vdd gnd OAI21X1
X_10345_ _10345_/A _10345_/B _10345_/C _10345_/Y vdd gnd NAND3X1
XFILL_1__9648_ vdd gnd FILL
XFILL_2__8441_ vdd gnd FILL
X_13064_ _13064_/A _13064_/B _13064_/Y vdd gnd NAND2X1
X_10276_ _10276_/A _10276_/B _10276_/Y vdd gnd AND2X2
XFILL_1__9579_ vdd gnd FILL
XFILL_2__8372_ vdd gnd FILL
X_12015_ _12015_/A _12015_/B _12015_/C _12015_/Y vdd gnd OAI21X1
XFILL_1__11110_ vdd gnd FILL
XFILL_2__10661_ vdd gnd FILL
XFILL_0__11840_ vdd gnd FILL
XFILL_1__12090_ vdd gnd FILL
XFILL_1__11041_ vdd gnd FILL
XFILL_2__10592_ vdd gnd FILL
XFILL_0__11771_ vdd gnd FILL
X_13966_ _13966_/A _13966_/B _13966_/C _13966_/Y vdd gnd OAI21X1
XFILL_0__13510_ vdd gnd FILL
XFILL_0__14490_ vdd gnd FILL
X_12917_ _12917_/A _12917_/Y vdd gnd INVX1
X_13897_ _13897_/A _13897_/B _13897_/C _13897_/Y vdd gnd AOI21X1
XFILL_1__14800_ vdd gnd FILL
XFILL_0__10653_ vdd gnd FILL
XFILL_1__12992_ vdd gnd FILL
XFILL_2__14001_ vdd gnd FILL
X_12848_ _12848_/A _12848_/B _12848_/Y vdd gnd NAND2X1
XFILL_2__11213_ vdd gnd FILL
XFILL_1__14731_ vdd gnd FILL
XFILL_1__11943_ vdd gnd FILL
XFILL_2__12193_ vdd gnd FILL
XFILL_0__13372_ vdd gnd FILL
XFILL_0__10584_ vdd gnd FILL
X_12779_ _12779_/A _12779_/B _12779_/Y vdd gnd NOR2X1
XFILL_2__11144_ vdd gnd FILL
XFILL_0__12323_ vdd gnd FILL
XFILL_1__14662_ vdd gnd FILL
X_14518_ _14518_/D _14518_/CLK _14518_/Q vdd gnd DFFPOSX1
XFILL_1__11874_ vdd gnd FILL
XFILL_0__9890_ vdd gnd FILL
XFILL_1__13613_ vdd gnd FILL
XFILL_0__12254_ vdd gnd FILL
XFILL_1__10825_ vdd gnd FILL
XFILL_1__14593_ vdd gnd FILL
X_14449_ _14449_/A _14449_/Y vdd gnd INVX1
X_7380_ _7380_/A _7380_/Y vdd gnd INVX1
XFILL_0__11205_ vdd gnd FILL
XFILL_1__13544_ vdd gnd FILL
XFILL_0__12185_ vdd gnd FILL
XFILL_0__8772_ vdd gnd FILL
XFILL_2__14834_ vdd gnd FILL
XFILL_2__8708_ vdd gnd FILL
XFILL_0__11136_ vdd gnd FILL
XFILL_1__10687_ vdd gnd FILL
X_9050_ _9050_/A _9050_/B _9050_/C _9050_/Y vdd gnd AOI21X1
XFILL_0__7723_ vdd gnd FILL
XFILL_2__8639_ vdd gnd FILL
XFILL_2__14765_ vdd gnd FILL
XFILL_1__12426_ vdd gnd FILL
XFILL_0__11067_ vdd gnd FILL
XFILL_2__11977_ vdd gnd FILL
X_8001_ _8001_/A _8001_/Y vdd gnd INVX4
XFILL_0__7654_ vdd gnd FILL
XFILL_0__10018_ vdd gnd FILL
XFILL_2__14696_ vdd gnd FILL
XFILL_1__12357_ vdd gnd FILL
XFILL_0__7585_ vdd gnd FILL
XFILL_1__11308_ vdd gnd FILL
XFILL_0__14826_ vdd gnd FILL
XFILL_0__9324_ vdd gnd FILL
XFILL_1__12288_ vdd gnd FILL
X_9952_ _9952_/A _9952_/B _9952_/Y vdd gnd NAND2X1
XFILL_1__14027_ vdd gnd FILL
XFILL_1__11239_ vdd gnd FILL
XFILL_0__14757_ vdd gnd FILL
XFILL_0__9255_ vdd gnd FILL
XFILL_0__11969_ vdd gnd FILL
X_8903_ _8903_/D _8903_/CLK _8903_/Q vdd gnd DFFPOSX1
X_9883_ _9883_/A _9883_/B _9883_/C _9883_/Y vdd gnd OAI21X1
XFILL_0__13708_ vdd gnd FILL
XFILL_0__8206_ vdd gnd FILL
XFILL_0__14688_ vdd gnd FILL
XFILL_0__9186_ vdd gnd FILL
X_8834_ _8834_/A _8834_/B _8834_/C _8834_/Y vdd gnd OAI21X1
XFILL_0__13639_ vdd gnd FILL
XFILL_0__8137_ vdd gnd FILL
X_8765_ _8765_/A _8765_/B _8765_/C _8765_/Y vdd gnd OAI21X1
XFILL_1__8950_ vdd gnd FILL
X_7716_ _7716_/A _7716_/Y vdd gnd INVX1
XFILL_0__8068_ vdd gnd FILL
X_8696_ _8696_/A _8696_/B _8696_/Y vdd gnd NAND2X1
XFILL_1__7901_ vdd gnd FILL
X_7647_ _7647_/A _7647_/B _7647_/C _7647_/Y vdd gnd NAND3X1
XFILL_1__7832_ vdd gnd FILL
X_7578_ _7578_/A _7578_/B _7578_/C _7578_/Y vdd gnd NOR3X1
X_9317_ _9317_/A _9317_/B _9317_/C _9317_/Y vdd gnd OAI21X1
XFILL_1__7763_ vdd gnd FILL
XFILL_1__9502_ vdd gnd FILL
X_9248_ _9248_/A _9248_/B _9248_/Y vdd gnd NAND2X1
XFILL_1__7694_ vdd gnd FILL
X_10130_ _10130_/A _10130_/B _10130_/C _10130_/Y vdd gnd NAND3X1
XFILL_1__9433_ vdd gnd FILL
X_9179_ _9179_/A _9179_/B _9179_/Y vdd gnd NOR2X1
X_10061_ _10061_/A _10061_/Y vdd gnd INVX1
XFILL_1__9364_ vdd gnd FILL
XFILL_1__8315_ vdd gnd FILL
XFILL_1__9295_ vdd gnd FILL
X_13820_ _13820_/A _13820_/B _13820_/C _13820_/Y vdd gnd NAND3X1
XFILL_1__8246_ vdd gnd FILL
X_13751_ _13751_/A _13751_/B _13751_/Y vdd gnd NAND2X1
X_10963_ _10963_/A _10963_/B _10963_/C _10963_/Y vdd gnd OAI21X1
XFILL_1__8177_ vdd gnd FILL
X_12702_ _12702_/A _12702_/B _12702_/C _12702_/Y vdd gnd AOI21X1
XFILL_1__7128_ vdd gnd FILL
X_13682_ _13682_/A _13682_/B _13682_/Y vdd gnd OR2X2
X_10894_ _10894_/A _10894_/B _10894_/C _10894_/Y vdd gnd NAND3X1
XFILL_2__8990_ vdd gnd FILL
X_12633_ _12633_/A _12633_/Y vdd gnd INVX1
XFILL_1_CLKBUF1_insert80 vdd gnd FILL
XFILL_1_CLKBUF1_insert91 vdd gnd FILL
X_12564_ _12564_/D _12564_/CLK _12564_/Q vdd gnd DFFPOSX1
XFILL_2__7872_ vdd gnd FILL
X_14303_ _14303_/A _14303_/B _14303_/C _14303_/Y vdd gnd NAND3X1
X_11515_ _11515_/A _11515_/B _11515_/C _11515_/Y vdd gnd NAND3X1
X_12495_ _12495_/A _12495_/B _12495_/C _12495_/Y vdd gnd OAI21X1
XFILL_1__10610_ vdd gnd FILL
XFILL_1__11590_ vdd gnd FILL
X_14234_ _14234_/A _14234_/Y vdd gnd INVX1
X_11446_ _11446_/A _11446_/B _11446_/C _11446_/Y vdd gnd OAI21X1
XFILL_2__11900_ vdd gnd FILL
XFILL_1__10541_ vdd gnd FILL
X_14165_ _14165_/D _14165_/CLK _14165_/Q vdd gnd DFFPOSX1
X_11377_ _11377_/A _11377_/B _11377_/Y vdd gnd NOR2X1
XFILL_2__11831_ vdd gnd FILL
XFILL_1__10472_ vdd gnd FILL
XFILL_1__13260_ vdd gnd FILL
X_13116_ _13116_/A _13116_/Y vdd gnd INVX1
X_10328_ _10328_/A _10328_/B _10328_/Y vdd gnd NAND2X1
XFILL_0__13990_ vdd gnd FILL
XFILL_2__8424_ vdd gnd FILL
X_14096_ _14096_/A _14096_/B _14096_/Y vdd gnd AND2X2
XFILL_1__12211_ vdd gnd FILL
XFILL_1__13191_ vdd gnd FILL
XFILL_2__11762_ vdd gnd FILL
XFILL_0__12941_ vdd gnd FILL
X_13047_ _13047_/A _13047_/B _13047_/Y vdd gnd NAND2X1
X_10259_ _10259_/A _10259_/B _10259_/Y vdd gnd NAND2X1
XFILL_2__8355_ vdd gnd FILL
XFILL_1__12142_ vdd gnd FILL
XFILL_2__11693_ vdd gnd FILL
XFILL_0__12872_ vdd gnd FILL
XFILL_0__7370_ vdd gnd FILL
XFILL_0__14611_ vdd gnd FILL
XFILL_2__10644_ vdd gnd FILL
XFILL_2__8286_ vdd gnd FILL
XFILL_1__12073_ vdd gnd FILL
XFILL_0__11823_ vdd gnd FILL
XFILL_1__11024_ vdd gnd FILL
XFILL_2__13363_ vdd gnd FILL
XFILL_2__10575_ vdd gnd FILL
XFILL_0__9040_ vdd gnd FILL
XFILL_0__11754_ vdd gnd FILL
X_13949_ _13949_/A _13949_/B _13949_/C _13949_/Y vdd gnd OAI21X1
XFILL_0__14473_ vdd gnd FILL
XFILL_0__10636_ vdd gnd FILL
XFILL_0__13424_ vdd gnd FILL
XFILL_1__12975_ vdd gnd FILL
X_8550_ _8550_/A _8550_/Y vdd gnd INVX1
XFILL_1__14714_ vdd gnd FILL
XFILL_1__11926_ vdd gnd FILL
XFILL_0__10567_ vdd gnd FILL
XFILL_0__13355_ vdd gnd FILL
X_7501_ _7501_/A _7501_/Y vdd gnd INVX1
XFILL_0__9942_ vdd gnd FILL
X_8481_ _8481_/A _8481_/B _8481_/C _8481_/Y vdd gnd OAI21X1
XFILL_2__11127_ vdd gnd FILL
XFILL_1__14645_ vdd gnd FILL
XFILL_0__12306_ vdd gnd FILL
XFILL_1__11857_ vdd gnd FILL
XFILL_0__13286_ vdd gnd FILL
XFILL_0__10498_ vdd gnd FILL
X_7432_ _7432_/A _7432_/B _7432_/C _7432_/Y vdd gnd OAI21X1
XFILL_0__9873_ vdd gnd FILL
XFILL_2__11058_ vdd gnd FILL
XFILL_0__12237_ vdd gnd FILL
XFILL_1__10808_ vdd gnd FILL
XFILL_1__14576_ vdd gnd FILL
XFILL_0__8824_ vdd gnd FILL
XFILL_1__11788_ vdd gnd FILL
X_7363_ _7363_/A _7363_/B _7363_/C _7363_/Y vdd gnd NAND3X1
XFILL_1__13527_ vdd gnd FILL
XFILL_0__12168_ vdd gnd FILL
X_9102_ _9102_/A _9102_/B _9102_/C _9102_/Y vdd gnd AOI21X1
XFILL_0__8755_ vdd gnd FILL
X_7294_ _7294_/A _7294_/B _7294_/Y vdd gnd NAND2X1
XFILL_2__14817_ vdd gnd FILL
XFILL_0__11119_ vdd gnd FILL
XFILL_0__7706_ vdd gnd FILL
XFILL_0__12099_ vdd gnd FILL
X_9033_ _9033_/A _9033_/B _9033_/S _9033_/Y vdd gnd MUX2X1
XFILL_0__8686_ vdd gnd FILL
XFILL_2__14748_ vdd gnd FILL
XFILL_1__12409_ vdd gnd FILL
XFILL_1__13389_ vdd gnd FILL
XFILL_0__7637_ vdd gnd FILL
XFILL_2__14679_ vdd gnd FILL
XFILL_0__7568_ vdd gnd FILL
XFILL_0__14809_ vdd gnd FILL
XFILL_0__9307_ vdd gnd FILL
XFILL_1__8100_ vdd gnd FILL
XFILL_1__9080_ vdd gnd FILL
X_9935_ _9935_/A _9935_/Y vdd gnd INVX2
XFILL_0__7499_ vdd gnd FILL
XFILL_0__9238_ vdd gnd FILL
XFILL_1__8031_ vdd gnd FILL
X_9866_ _9866_/A _9866_/B _9866_/C _9866_/D _9866_/Y vdd gnd AOI22X1
XFILL_0__9169_ vdd gnd FILL
X_8817_ _8817_/A _8817_/B _8817_/C _8817_/Y vdd gnd OAI21X1
X_9797_ _9797_/D _9797_/CLK _9797_/Q vdd gnd DFFPOSX1
XFILL_1__9982_ vdd gnd FILL
X_8748_ _8748_/A _8748_/B _8748_/Y vdd gnd NAND2X1
XFILL_1__8933_ vdd gnd FILL
X_8679_ _8679_/A _8679_/B _8679_/Y vdd gnd NAND2X1
XFILL_1_CLKBUF1_insert102 vdd gnd FILL
X_11300_ _11300_/A _11300_/B _11300_/C _11300_/Y vdd gnd OAI21X1
XFILL_1__7815_ vdd gnd FILL
X_12280_ _12280_/A _12280_/B _12280_/C _12280_/Y vdd gnd OAI21X1
XFILL_1__8795_ vdd gnd FILL
X_11231_ _11231_/A _11231_/B _11231_/C _11231_/Y vdd gnd OAI21X1
XFILL_1__7746_ vdd gnd FILL
X_11162_ _11162_/A _11162_/B _11162_/C _11162_/Y vdd gnd OAI21X1
XFILL_1__7677_ vdd gnd FILL
X_10113_ _10113_/A _10113_/B _10113_/C _10113_/Y vdd gnd NAND3X1
XFILL_1__9416_ vdd gnd FILL
X_11093_ _11093_/A _11093_/B _11093_/C _11093_/Y vdd gnd AOI21X1
X_10044_ _10044_/A _10044_/B _10044_/Y vdd gnd NOR2X1
XFILL_1__9347_ vdd gnd FILL
XFILL257550x194550 vdd gnd FILL
X_14852_ _14852_/A _14852_/B _14852_/C _14852_/Y vdd gnd OAI21X1
XFILL_1__9278_ vdd gnd FILL
X_13803_ _13803_/A _13803_/B _13803_/Y vdd gnd AND2X2
X_14783_ _14783_/A _14783_/B _14783_/C _14783_/Y vdd gnd NAND3X1
XFILL_1__8229_ vdd gnd FILL
X_11995_ _11995_/A _11995_/B _11995_/C _11995_/Y vdd gnd OAI21X1
X_13734_ _13734_/A _13734_/B _13734_/C _13734_/D _13734_/Y vdd gnd AOI22X1
X_10946_ _10946_/A _10946_/B _10946_/C _10946_/Y vdd gnd NAND3X1
XFILL_2__10291_ vdd gnd FILL
XFILL_0__11470_ vdd gnd FILL
X_13665_ _13665_/A _13665_/B _13665_/C _13665_/Y vdd gnd AOI21X1
X_10877_ _10877_/A _10877_/B _10877_/C _10877_/Y vdd gnd OAI21X1
XFILL_0__10421_ vdd gnd FILL
XFILL_1__12760_ vdd gnd FILL
X_12616_ _12616_/A _12616_/Y vdd gnd INVX2
X_13596_ _13596_/A _13596_/Y vdd gnd INVX1
XFILL_1__11711_ vdd gnd FILL
XFILL_0__13140_ vdd gnd FILL
XFILL_0__10352_ vdd gnd FILL
XFILL_1__12691_ vdd gnd FILL
X_12547_ _12547_/D _12547_/CLK _12547_/Q vdd gnd DFFPOSX1
XFILL_1__14430_ vdd gnd FILL
XFILL_0__13071_ vdd gnd FILL
XFILL_0__10283_ vdd gnd FILL
X_12478_ _12478_/A _12478_/B _12478_/C _12478_/Y vdd gnd OAI21X1
XFILL_0__12022_ vdd gnd FILL
XFILL_1__14361_ vdd gnd FILL
X_14217_ _14217_/A _14217_/B _14217_/Y vdd gnd NAND2X1
XFILL_1__11573_ vdd gnd FILL
X_11429_ _11429_/A _11429_/B _11429_/C _11429_/Y vdd gnd OAI21X1
XFILL_1__13312_ vdd gnd FILL
XFILL_1__10524_ vdd gnd FILL
XFILL_1__14292_ vdd gnd FILL
XFILL_0__8540_ vdd gnd FILL
XCLKBUF1_insert101 CLKBUF1_insert101/A CLKBUF1_insert101/Y vdd gnd CLKBUF1
X_14148_ _14148_/A _14148_/B _14148_/C _14148_/Y vdd gnd OAI21X1
XFILL_1__13243_ vdd gnd FILL
XFILL_1__10455_ vdd gnd FILL
XFILL_0__13973_ vdd gnd FILL
XFILL_0__8471_ vdd gnd FILL
X_14079_ _14079_/A _14079_/B _14079_/Y vdd gnd OR2X2
XFILL_2__11745_ vdd gnd FILL
XFILL_1__13174_ vdd gnd FILL
XFILL_1__10386_ vdd gnd FILL
XFILL_0__12924_ vdd gnd FILL
XFILL_0__7422_ vdd gnd FILL
XFILL_2__8338_ vdd gnd FILL
XFILL_1__12125_ vdd gnd FILL
XFILL_0__12855_ vdd gnd FILL
XFILL_0__7353_ vdd gnd FILL
XFILL_2__13415_ vdd gnd FILL
XFILL_2__10627_ vdd gnd FILL
X_7981_ _7981_/D _7981_/CLK _7981_/Q vdd gnd DFFPOSX1
XFILL_2__8269_ vdd gnd FILL
XFILL_1__12056_ vdd gnd FILL
XFILL_0__11806_ vdd gnd FILL
X_9720_ _9720_/A _9720_/B _9720_/C _9720_/Y vdd gnd OAI21X1
XFILL_0__12786_ vdd gnd FILL
XFILL_0__7284_ vdd gnd FILL
XFILL_1__11007_ vdd gnd FILL
XFILL_2__13346_ vdd gnd FILL
XFILL257550x216150 vdd gnd FILL
XFILL_2__10558_ vdd gnd FILL
XFILL_0__9023_ vdd gnd FILL
XFILL_0__11737_ vdd gnd FILL
X_9651_ _9651_/A _9651_/B _9651_/C _9651_/Y vdd gnd AOI21X1
XFILL_2__13277_ vdd gnd FILL
XFILL_2__10489_ vdd gnd FILL
XFILL_0__14456_ vdd gnd FILL
X_8602_ _8602_/A _8602_/B _8602_/Y vdd gnd NAND2X1
X_9582_ _9582_/A _9582_/B _9582_/C _9582_/Y vdd gnd AOI21X1
XFILL_0__13407_ vdd gnd FILL
XFILL_0__10619_ vdd gnd FILL
XFILL_1__12958_ vdd gnd FILL
XFILL_0__14387_ vdd gnd FILL
XFILL_0__11599_ vdd gnd FILL
XCLKBUF1_insert60 CLKBUF1_insert60/A CLKBUF1_insert60/Y vdd gnd CLKBUF1
X_8533_ _8533_/A _8533_/B _8533_/C _8533_/Y vdd gnd NAND3X1
XFILL_1__11909_ vdd gnd FILL
XCLKBUF1_insert71 CLKBUF1_insert71/A CLKBUF1_insert71/Y vdd gnd CLKBUF1
XCLKBUF1_insert82 CLKBUF1_insert82/A CLKBUF1_insert82/Y vdd gnd CLKBUF1
XFILL_0__13338_ vdd gnd FILL
XCLKBUF1_insert93 CLKBUF1_insert93/A CLKBUF1_insert93/Y vdd gnd CLKBUF1
XFILL_1__12889_ vdd gnd FILL
XFILL_0__9925_ vdd gnd FILL
X_8464_ _8464_/A _8464_/B _8464_/Y vdd gnd NOR2X1
XFILL_1__14628_ vdd gnd FILL
XFILL_0__13269_ vdd gnd FILL
X_7415_ _7415_/A _7415_/B _7415_/C _7415_/Y vdd gnd OAI21X1
XFILL_0__9856_ vdd gnd FILL
X_8395_ _8395_/A _8395_/B _8395_/C _8395_/Y vdd gnd OAI21X1
XFILL_1__14559_ vdd gnd FILL
XFILL_1__7600_ vdd gnd FILL
XFILL_0__8807_ vdd gnd FILL
X_7346_ _7346_/A _7346_/B _7346_/C _7346_/Y vdd gnd OAI21X1
XFILL_1__8580_ vdd gnd FILL
XFILL_1__7531_ vdd gnd FILL
XFILL_0__8738_ vdd gnd FILL
X_7277_ _7277_/A _7277_/B _7277_/C _7277_/Y vdd gnd OAI21X1
X_9016_ _9016_/A _9016_/B _9016_/C _9016_/Y vdd gnd NAND3X1
XFILL_1__7462_ vdd gnd FILL
XFILL_0__8669_ vdd gnd FILL
XFILL_1__9201_ vdd gnd FILL
XFILL_1__7393_ vdd gnd FILL
XFILL_1__9132_ vdd gnd FILL
XFILL_1__9063_ vdd gnd FILL
X_9918_ _9918_/A _9918_/B _9918_/C _9918_/Y vdd gnd OAI21X1
XFILL257550x126150 vdd gnd FILL
X_10800_ _10800_/A _10800_/B _10800_/Y vdd gnd NAND2X1
XFILL_1__8014_ vdd gnd FILL
X_11780_ _11780_/A _11780_/B _11780_/S _11780_/Y vdd gnd MUX2X1
X_9849_ _9849_/A _9849_/Y vdd gnd INVX4
X_10731_ _10731_/D _10731_/CLK _10731_/Q vdd gnd DFFPOSX1
X_13450_ _13450_/D _13450_/CLK _13450_/Q vdd gnd DFFPOSX1
X_10662_ _10662_/A _10662_/B _10662_/Y vdd gnd NAND2X1
XFILL_1__9965_ vdd gnd FILL
X_12401_ _12401_/A _12401_/Y vdd gnd INVX1
X_13381_ _13381_/A _13381_/B _13381_/C _13381_/Y vdd gnd OAI21X1
X_10593_ _10593_/A _10593_/B _10593_/C _10593_/Y vdd gnd AOI21X1
XFILL_1__9896_ vdd gnd FILL
X_12332_ _12332_/A _12332_/B _12332_/S _12332_/Y vdd gnd MUX2X1
X_12263_ _12263_/A _12263_/Y vdd gnd INVX1
XFILL_1__8778_ vdd gnd FILL
X_14002_ _14002_/A _14002_/B _14002_/Y vdd gnd NAND2X1
X_11214_ _11214_/A _11214_/B _11214_/C _11214_/Y vdd gnd OAI21X1
XFILL_2__9310_ vdd gnd FILL
XFILL_1__7729_ vdd gnd FILL
X_12194_ _12194_/A _12194_/B _12194_/C _12194_/Y vdd gnd AOI21X1
X_11145_ _11145_/A _11145_/B _11145_/Y vdd gnd AND2X2
XFILL_2__9241_ vdd gnd FILL
XFILL_1__10240_ vdd gnd FILL
XFILL_0__10970_ vdd gnd FILL
X_11076_ _11076_/A _11076_/Y vdd gnd INVX1
XFILL_2__9172_ vdd gnd FILL
XFILL_2__11530_ vdd gnd FILL
XFILL_1__10171_ vdd gnd FILL
X_14904_ _14904_/D _14904_/CLK _14904_/Q vdd gnd DFFPOSX1
X_10027_ _10027_/A _10027_/B _10027_/C _10027_/Y vdd gnd OAI21X1
XFILL_2__11461_ vdd gnd FILL
XFILL_0__12640_ vdd gnd FILL
X_14835_ _14835_/A _14835_/B _14835_/C _14835_/Y vdd gnd OAI21X1
XFILL_1__13930_ vdd gnd FILL
XFILL_2__13131_ vdd gnd FILL
X_14766_ _14766_/A _14766_/B _14766_/C _14766_/Y vdd gnd OAI21X1
X_11978_ _11978_/A _11978_/B _11978_/C _11978_/Y vdd gnd NAND3X1
XFILL_0__14310_ vdd gnd FILL
XFILL_1__13861_ vdd gnd FILL
XFILL_0__11522_ vdd gnd FILL
X_10929_ _10929_/A _10929_/B _10929_/C _10929_/Y vdd gnd OAI21X1
X_13717_ _13717_/A _13717_/B _13717_/Y vdd gnd NAND2X1
X_14697_ _14697_/A _14697_/B _14697_/Y vdd gnd NAND2X1
XFILL_1__12812_ vdd gnd FILL
XFILL_2__13062_ vdd gnd FILL
XFILL_0__14241_ vdd gnd FILL
XFILL_0__11453_ vdd gnd FILL
XFILL_1__13792_ vdd gnd FILL
X_13648_ _13648_/A _13648_/Y vdd gnd INVX1
XFILL_0__10404_ vdd gnd FILL
XFILL_1__12743_ vdd gnd FILL
XFILL_0_BUFX2_insert230 vdd gnd FILL
XFILL_0__11384_ vdd gnd FILL
XFILL_0_BUFX2_insert241 vdd gnd FILL
XFILL_0_BUFX2_insert252 vdd gnd FILL
X_13579_ _13579_/A _13579_/B _13579_/C _13579_/Y vdd gnd AOI21X1
XFILL_0_BUFX2_insert263 vdd gnd FILL
XFILL_0__13123_ vdd gnd FILL
XFILL_0__10335_ vdd gnd FILL
XFILL_0_BUFX2_insert274 vdd gnd FILL
XFILL_0_BUFX2_insert285 vdd gnd FILL
XFILL_1__12674_ vdd gnd FILL
XFILL_0__9710_ vdd gnd FILL
XFILL_0_BUFX2_insert296 vdd gnd FILL
XFILL_1__14413_ vdd gnd FILL
XFILL_0__13054_ vdd gnd FILL
XFILL_0__10266_ vdd gnd FILL
X_7200_ _7200_/A _7200_/B _7200_/C _7200_/Y vdd gnd OAI21X1
XFILL_0__9641_ vdd gnd FILL
X_8180_ _8180_/A _8180_/B _8180_/C _8180_/D _8180_/Y vdd gnd AOI22X1
XFILL_2__12915_ vdd gnd FILL
XFILL_0__12005_ vdd gnd FILL
XFILL_1__14344_ vdd gnd FILL
XFILL_1__11556_ vdd gnd FILL
XFILL_0__10197_ vdd gnd FILL
X_7131_ _7131_/A _7131_/Y vdd gnd INVX1
XFILL_0__9572_ vdd gnd FILL
XFILL_2__9508_ vdd gnd FILL
XFILL_1__10507_ vdd gnd FILL
XFILL_1__14275_ vdd gnd FILL
XFILL_0__8523_ vdd gnd FILL
XFILL_1__11487_ vdd gnd FILL
XFILL_1__13226_ vdd gnd FILL
XFILL_1__10438_ vdd gnd FILL
XFILL_0__13956_ vdd gnd FILL
XFILL_0__8454_ vdd gnd FILL
XFILL_1__13157_ vdd gnd FILL
XFILL_0__12907_ vdd gnd FILL
XFILL_1__10369_ vdd gnd FILL
XFILL_0__7405_ vdd gnd FILL
XFILL_0__13887_ vdd gnd FILL
XFILL_0__8385_ vdd gnd FILL
XFILL_1__12108_ vdd gnd FILL
XFILL_2__14447_ vdd gnd FILL
XFILL_1__13088_ vdd gnd FILL
XFILL_0__12838_ vdd gnd FILL
XFILL_0__7336_ vdd gnd FILL
X_7964_ _7964_/D _7964_/CLK _7964_/Q vdd gnd DFFPOSX1
XFILL_1__12039_ vdd gnd FILL
XFILL_2__14378_ vdd gnd FILL
X_9703_ _9703_/A _9703_/B _9703_/C _9703_/Y vdd gnd OAI21X1
XFILL_0__12769_ vdd gnd FILL
XFILL_0__7267_ vdd gnd FILL
XFILL_2__13329_ vdd gnd FILL
X_7895_ _7895_/A _7895_/B _7895_/C _7895_/Y vdd gnd OAI21X1
XFILL_0__9006_ vdd gnd FILL
X_9634_ _9634_/A _9634_/B _9634_/Y vdd gnd NAND2X1
XFILL_0__7198_ vdd gnd FILL
XFILL_0__14439_ vdd gnd FILL
X_9565_ _9565_/A _9565_/B _9565_/Y vdd gnd NOR2X1
X_8516_ _8516_/A _8516_/B _8516_/C _8516_/Y vdd gnd NAND3X1
XFILL_1__9750_ vdd gnd FILL
X_9496_ _9496_/A _9496_/B _9496_/Y vdd gnd NAND2X1
XFILL_0__9908_ vdd gnd FILL
XFILL_1__8701_ vdd gnd FILL
XFILL_1__9681_ vdd gnd FILL
X_8447_ _8447_/A _8447_/B _8447_/C _8447_/Y vdd gnd NAND3X1
XFILL_1__8632_ vdd gnd FILL
X_8378_ _8378_/A _8378_/B _8378_/C _8378_/Y vdd gnd OAI21X1
X_7329_ _7329_/A _7329_/B _7329_/C _7329_/Y vdd gnd NAND3X1
XFILL_1__8563_ vdd gnd FILL
XFILL_1__7514_ vdd gnd FILL
XFILL_1__8494_ vdd gnd FILL
XFILL_1__7445_ vdd gnd FILL
XFILL_0_CLKBUF1_insert29 vdd gnd FILL
XFILL_2_BUFX2_insert303 vdd gnd FILL
X_12950_ _12950_/A _12950_/B _12950_/C _12950_/Y vdd gnd NAND3X1
XFILL_1__7376_ vdd gnd FILL
XFILL_2_BUFX2_insert325 vdd gnd FILL
X_11901_ _11901_/A _11901_/B _11901_/C _11901_/Y vdd gnd NAND3X1
XFILL_1__9115_ vdd gnd FILL
XFILL_2_BUFX2_insert358 vdd gnd FILL
X_12881_ _12881_/A _12881_/B _12881_/Y vdd gnd NOR2X1
X_14620_ _14620_/A _14620_/B _14620_/Y vdd gnd NOR2X1
X_11832_ _11832_/A _11832_/B _11832_/Y vdd gnd NAND2X1
XFILL_1__9046_ vdd gnd FILL
X_14551_ _14551_/D _14551_/CLK _14551_/Q vdd gnd DFFPOSX1
X_11763_ _11763_/A _11763_/B _11763_/C _11763_/Y vdd gnd OAI21X1
X_10714_ _10714_/D _10714_/CLK _10714_/Q vdd gnd DFFPOSX1
X_13502_ _13502_/A _13502_/Y vdd gnd INVX2
XBUFX2_insert302 BUFX2_insert302/A BUFX2_insert302/Y vdd gnd BUFX2
XBUFX2_insert313 BUFX2_insert313/A BUFX2_insert313/Y vdd gnd BUFX2
X_14482_ _14482_/A _14482_/B _14482_/Y vdd gnd NAND2X1
XFILL_2__8810_ vdd gnd FILL
X_11694_ _11694_/A _11694_/B _11694_/Y vdd gnd NOR2X1
XBUFX2_insert324 BUFX2_insert324/A BUFX2_insert324/Y vdd gnd BUFX2
XBUFX2_insert335 BUFX2_insert335/A BUFX2_insert335/Y vdd gnd BUFX2
XBUFX2_insert346 BUFX2_insert346/A BUFX2_insert346/Y vdd gnd BUFX2
X_13433_ _13433_/D _13433_/CLK _13433_/Q vdd gnd DFFPOSX1
X_10645_ _10645_/A _10645_/B _10645_/C _10645_/Y vdd gnd OAI21X1
XBUFX2_insert357 BUFX2_insert357/A BUFX2_insert357/Y vdd gnd BUFX2
XBUFX2_insert368 BUFX2_insert368/A BUFX2_insert368/Y vdd gnd BUFX2
XFILL_1__9948_ vdd gnd FILL
XFILL_2__8741_ vdd gnd FILL
XBUFX2_insert379 BUFX2_insert379/A BUFX2_insert379/Y vdd gnd BUFX2
X_13364_ _13364_/A _13364_/B _13364_/Y vdd gnd NAND2X1
X_10576_ _10576_/A _10576_/B _10576_/C _10576_/Y vdd gnd NAND3X1
XFILL_0__10120_ vdd gnd FILL
XFILL_2__8672_ vdd gnd FILL
XFILL_1__9879_ vdd gnd FILL
X_12315_ _12315_/A _12315_/B _12315_/Y vdd gnd NOR2X1
X_13295_ _13295_/A _13295_/B _13295_/C _13295_/Y vdd gnd OAI21X1
XFILL_1__11410_ vdd gnd FILL
XFILL_0__10051_ vdd gnd FILL
XFILL_1__12390_ vdd gnd FILL
X_12246_ _12246_/A _12246_/Y vdd gnd INVX1
XFILL_2__12700_ vdd gnd FILL
XFILL_1__11341_ vdd gnd FILL
XFILL_2__13680_ vdd gnd FILL
X_12177_ _12177_/A _12177_/B _12177_/C _12177_/Y vdd gnd OAI21X1
XFILL_2__12631_ vdd gnd FILL
XFILL_1__14060_ vdd gnd FILL
XFILL_0__13810_ vdd gnd FILL
XFILL_1__11272_ vdd gnd FILL
XFILL_0__14790_ vdd gnd FILL
X_11128_ _11128_/A _11128_/B _11128_/C _11128_/Y vdd gnd OAI21X1
XFILL_2__9224_ vdd gnd FILL
XFILL_1__13011_ vdd gnd FILL
XFILL_1__10223_ vdd gnd FILL
XFILL_0__13741_ vdd gnd FILL
XFILL_0__10953_ vdd gnd FILL
X_11059_ _11059_/A _11059_/B _11059_/C _11059_/Y vdd gnd NAND3X1
XFILL_2__14301_ vdd gnd FILL
XFILL_2__9155_ vdd gnd FILL
XFILL_2__11513_ vdd gnd FILL
XFILL_1__10154_ vdd gnd FILL
XFILL_0__13672_ vdd gnd FILL
XFILL_0__8170_ vdd gnd FILL
XFILL_0__10884_ vdd gnd FILL
XFILL_2__14232_ vdd gnd FILL
XFILL_2__9086_ vdd gnd FILL
XFILL_2__11444_ vdd gnd FILL
XFILL_1__10085_ vdd gnd FILL
XFILL_0__12623_ vdd gnd FILL
XFILL_0__7121_ vdd gnd FILL
X_14818_ _14818_/A _14818_/B _14818_/C _14818_/Y vdd gnd AOI21X1
XFILL_1__13913_ vdd gnd FILL
XFILL_2__11375_ vdd gnd FILL
X_14749_ _14749_/A _14749_/Y vdd gnd INVX1
X_7680_ _7680_/A _7680_/B _7680_/C _7680_/Y vdd gnd AOI21X1
XFILL_0__11505_ vdd gnd FILL
XFILL_1__13844_ vdd gnd FILL
XFILL_2__14094_ vdd gnd FILL
XFILL_0__12485_ vdd gnd FILL
XFILL_0__14224_ vdd gnd FILL
XFILL_2__9988_ vdd gnd FILL
XFILL_0__11436_ vdd gnd FILL
XFILL_1__13775_ vdd gnd FILL
XFILL_1__10987_ vdd gnd FILL
X_9350_ _9350_/A _9350_/B _9350_/C _9350_/Y vdd gnd AOI21X1
XFILL_1__12726_ vdd gnd FILL
XFILL_0__14155_ vdd gnd FILL
X_8301_ _8301_/A _8301_/B _8301_/C _8301_/Y vdd gnd AOI21X1
XFILL_0__11367_ vdd gnd FILL
X_9281_ _9281_/A _9281_/B _9281_/Y vdd gnd NAND2X1
XFILL_0__13106_ vdd gnd FILL
XFILL_1__12657_ vdd gnd FILL
XFILL_0__10318_ vdd gnd FILL
XFILL_0__11298_ vdd gnd FILL
XFILL_0__14086_ vdd gnd FILL
X_8232_ _8232_/A _8232_/B _8232_/Y vdd gnd NAND2X1
XFILL_0__7885_ vdd gnd FILL
XFILL_1__11608_ vdd gnd FILL
XFILL_0__13037_ vdd gnd FILL
XFILL_0__10249_ vdd gnd FILL
XFILL_2__13947_ vdd gnd FILL
XFILL_0__9624_ vdd gnd FILL
X_8163_ _8163_/A _8163_/B _8163_/C _8163_/Y vdd gnd OAI21X1
XFILL_1__14327_ vdd gnd FILL
XFILL_1__11539_ vdd gnd FILL
X_7114_ _7114_/A _7114_/Y vdd gnd INVX1
XFILL_0__9555_ vdd gnd FILL
X_8094_ _8094_/A _8094_/Y vdd gnd INVX1
XFILL_1__14258_ vdd gnd FILL
XFILL_2__12829_ vdd gnd FILL
XFILL_0__8506_ vdd gnd FILL
XFILL_0__9486_ vdd gnd FILL
XFILL_1__13209_ vdd gnd FILL
XFILL_0__13939_ vdd gnd FILL
XFILL_1__7230_ vdd gnd FILL
XFILL_0__8437_ vdd gnd FILL
XFILL_1__7161_ vdd gnd FILL
XFILL_0__8368_ vdd gnd FILL
X_8996_ _8996_/A _8996_/B _8996_/S _8996_/Y vdd gnd MUX2X1
XFILL_0__7319_ vdd gnd FILL
XFILL_1__7092_ vdd gnd FILL
X_7947_ _7947_/D _7947_/CLK _7947_/Q vdd gnd DFFPOSX1
XFILL_0__8299_ vdd gnd FILL
X_7878_ _7878_/A _7878_/B _7878_/Y vdd gnd NAND2X1
X_9617_ _9617_/A _9617_/B _9617_/Y vdd gnd NOR2X1
X_9548_ _9548_/A _9548_/B _9548_/Y vdd gnd OR2X2
X_10430_ _10430_/A _10430_/B _10430_/C _10430_/Y vdd gnd NAND3X1
XFILL_1__9733_ vdd gnd FILL
X_9479_ _9479_/A _9479_/B _9479_/C _9479_/Y vdd gnd NAND3X1
X_10361_ _10361_/A _10361_/B _10361_/Y vdd gnd NOR2X1
XFILL_1__9664_ vdd gnd FILL
X_12100_ _12100_/A _12100_/B _12100_/Y vdd gnd AND2X2
X_13080_ _13080_/A _13080_/B _13080_/Y vdd gnd OR2X2
X_10292_ _10292_/A _10292_/B _10292_/C _10292_/Y vdd gnd OAI21X1
XFILL_1__8615_ vdd gnd FILL
XFILL_1__9595_ vdd gnd FILL
X_12031_ _12031_/A _12031_/B _12031_/C _12031_/Y vdd gnd AOI21X1
XFILL_1__8546_ vdd gnd FILL
XFILL_2__7270_ vdd gnd FILL
XFILL_1__8477_ vdd gnd FILL
XFILL_1__7428_ vdd gnd FILL
X_13982_ _13982_/A _13982_/B _13982_/Y vdd gnd NOR2X1
XFILL_2_BUFX2_insert122 vdd gnd FILL
X_12933_ _12933_/A _12933_/Y vdd gnd INVX1
XFILL_2_BUFX2_insert144 vdd gnd FILL
XFILL_1__7359_ vdd gnd FILL
XFILL_2_BUFX2_insert177 vdd gnd FILL
X_12864_ _12864_/A _12864_/B _12864_/C _12864_/Y vdd gnd AOI21X1
X_14603_ _14603_/A _14603_/B _14603_/Y vdd gnd NAND2X1
XFILL_1__9029_ vdd gnd FILL
X_11815_ _11815_/A _11815_/B _11815_/C _11815_/Y vdd gnd OAI21X1
X_12795_ _12795_/A _12795_/Y vdd gnd INVX1
XFILL_2__11160_ vdd gnd FILL
XFILL_1__10910_ vdd gnd FILL
XFILL_1__11890_ vdd gnd FILL
X_14534_ _14534_/D _14534_/CLK _14534_/Q vdd gnd DFFPOSX1
X_11746_ _11746_/A _11746_/B _11746_/C _11746_/D _11746_/Y vdd gnd AOI22X1
XBUFX2_insert110 BUFX2_insert110/A BUFX2_insert110/Y vdd gnd BUFX2
XFILL_2__11091_ vdd gnd FILL
XBUFX2_insert121 BUFX2_insert121/A BUFX2_insert121/Y vdd gnd BUFX2
XFILL_0__12270_ vdd gnd FILL
XFILL_1__10841_ vdd gnd FILL
XBUFX2_insert132 BUFX2_insert132/A BUFX2_insert132/Y vdd gnd BUFX2
XBUFX2_insert143 BUFX2_insert143/A BUFX2_insert143/Y vdd gnd BUFX2
X_14465_ _14465_/A _14465_/B _14465_/C _14465_/Y vdd gnd OAI21X1
X_11677_ _11677_/D _11677_/CLK _11677_/Q vdd gnd DFFPOSX1
XBUFX2_insert154 BUFX2_insert154/A BUFX2_insert154/Y vdd gnd BUFX2
XBUFX2_insert165 BUFX2_insert165/A BUFX2_insert165/Y vdd gnd BUFX2
XFILL_0__11221_ vdd gnd FILL
XFILL_1__13560_ vdd gnd FILL
XBUFX2_insert176 BUFX2_insert176/A BUFX2_insert176/Y vdd gnd BUFX2
XFILL_1__10772_ vdd gnd FILL
XBUFX2_insert187 BUFX2_insert187/A BUFX2_insert187/Y vdd gnd BUFX2
X_10628_ _10628_/A _10628_/B _10628_/C _10628_/Y vdd gnd OAI21X1
X_13416_ _13416_/A _13416_/B _13416_/Y vdd gnd NAND2X1
XBUFX2_insert198 BUFX2_insert198/A BUFX2_insert198/Y vdd gnd BUFX2
X_14396_ _14396_/A _14396_/B _14396_/C _14396_/Y vdd gnd OAI21X1
XFILL_1__12511_ vdd gnd FILL
XFILL_0__11152_ vdd gnd FILL
X_13347_ _13347_/A _13347_/B _13347_/Y vdd gnd NAND2X1
X_10559_ _10559_/A _10559_/B _10559_/Y vdd gnd NOR2X1
XFILL_0__10103_ vdd gnd FILL
XFILL_2__13801_ vdd gnd FILL
XFILL_2__8655_ vdd gnd FILL
XFILL_1__12442_ vdd gnd FILL
XFILL_0__11083_ vdd gnd FILL
XFILL_2__11993_ vdd gnd FILL
XFILL_0__7670_ vdd gnd FILL
X_13278_ _13278_/A _13278_/B _13278_/Y vdd gnd NAND2X1
XFILL_2__7606_ vdd gnd FILL
XFILL_0__14911_ vdd gnd FILL
XFILL_0__10034_ vdd gnd FILL
XFILL_2__13732_ vdd gnd FILL
XFILL_2__8586_ vdd gnd FILL
XFILL_1__12373_ vdd gnd FILL
X_12229_ _12229_/A _12229_/B _12229_/C _12229_/Y vdd gnd NAND3X1
XFILL_1__14112_ vdd gnd FILL
XFILL_2__13663_ vdd gnd FILL
XFILL_1__11324_ vdd gnd FILL
XFILL_0__14842_ vdd gnd FILL
XFILL_0__9340_ vdd gnd FILL
XFILL_1__14043_ vdd gnd FILL
XFILL_2__13594_ vdd gnd FILL
XFILL_1__11255_ vdd gnd FILL
XFILL_0__14773_ vdd gnd FILL
XFILL_0__9271_ vdd gnd FILL
XFILL_0__11985_ vdd gnd FILL
XFILL_2_CLKBUF1_insert391 vdd gnd FILL
XFILL_2__9207_ vdd gnd FILL
XFILL_1__10206_ vdd gnd FILL
XFILL_0__13724_ vdd gnd FILL
XFILL_1__11186_ vdd gnd FILL
XFILL_0__10936_ vdd gnd FILL
XFILL_0__8222_ vdd gnd FILL
X_8850_ _8850_/D _8850_/CLK _8850_/Q vdd gnd DFFPOSX1
XFILL_2__9138_ vdd gnd FILL
XFILL_1__10137_ vdd gnd FILL
XFILL_0__13655_ vdd gnd FILL
X_7801_ _7801_/A _7801_/B _7801_/C _7801_/Y vdd gnd OAI21X1
XFILL_0__8153_ vdd gnd FILL
XFILL_0__10867_ vdd gnd FILL
XFILL_2__9069_ vdd gnd FILL
X_8781_ _8781_/A _8781_/B _8781_/C _8781_/Y vdd gnd OAI21X1
XFILL_2__11427_ vdd gnd FILL
XFILL_0__7104_ vdd gnd FILL
XFILL_1__10068_ vdd gnd FILL
XFILL_0__13586_ vdd gnd FILL
X_7732_ _7732_/A _7732_/B _7732_/Y vdd gnd NOR2X1
XFILL_0__8084_ vdd gnd FILL
XFILL_0__10798_ vdd gnd FILL
XFILL_2__11358_ vdd gnd FILL
X_7663_ _7663_/A _7663_/B _7663_/C _7663_/Y vdd gnd OAI21X1
XFILL_1__13827_ vdd gnd FILL
XFILL_2__11289_ vdd gnd FILL
X_9402_ _9402_/A _9402_/B _9402_/Y vdd gnd NOR2X1
XFILL_0__12468_ vdd gnd FILL
X_7594_ _7594_/A _7594_/B _7594_/C _7594_/Y vdd gnd OAI21X1
XFILL_0__11419_ vdd gnd FILL
XFILL_1__13758_ vdd gnd FILL
X_9333_ _9333_/A _9333_/B _9333_/Y vdd gnd NAND2X1
XFILL_0__12399_ vdd gnd FILL
XFILL_1__12709_ vdd gnd FILL
XFILL_0__8986_ vdd gnd FILL
XFILL_0__14138_ vdd gnd FILL
XFILL_1__13689_ vdd gnd FILL
X_9264_ _9264_/A _9264_/B _9264_/Y vdd gnd OR2X2
XFILL_0__14069_ vdd gnd FILL
X_8215_ _8215_/A _8215_/B _8215_/C _8215_/Y vdd gnd NAND3X1
XFILL_0__7868_ vdd gnd FILL
X_9195_ _9195_/A _9195_/B _9195_/C _9195_/Y vdd gnd OAI21X1
XFILL_0__9607_ vdd gnd FILL
XFILL_1__8400_ vdd gnd FILL
XFILL_1__9380_ vdd gnd FILL
X_8146_ _8146_/A _8146_/Y vdd gnd INVX1
XFILL_0__7799_ vdd gnd FILL
XFILL_1__8331_ vdd gnd FILL
XFILL_0__9538_ vdd gnd FILL
X_8077_ _8077_/A _8077_/B _8077_/C _8077_/Y vdd gnd OAI21X1
XFILL_1__8262_ vdd gnd FILL
XFILL_0__9469_ vdd gnd FILL
XFILL_1__7213_ vdd gnd FILL
XFILL_1__8193_ vdd gnd FILL
XFILL_1__7144_ vdd gnd FILL
X_8979_ _8979_/A _8979_/Y vdd gnd INVX1
XFILL_1_BUFX2_insert118 vdd gnd FILL
XFILL_1_BUFX2_insert129 vdd gnd FILL
XFILL_1__7075_ vdd gnd FILL
X_11600_ _11600_/A _11600_/B _11600_/Y vdd gnd NAND2X1
X_12580_ _12580_/D _12580_/CLK _12580_/Q vdd gnd DFFPOSX1
X_11531_ _11531_/A _11531_/B _11531_/Y vdd gnd NAND2X1
X_14250_ _14250_/A _14250_/B _14250_/Y vdd gnd NAND2X1
X_11462_ _11462_/A _11462_/Y vdd gnd INVX1
X_13201_ _13201_/A _13201_/B _13201_/Y vdd gnd NAND2X1
X_10413_ _10413_/A _10413_/B _10413_/Y vdd gnd NOR2X1
X_14181_ _14181_/D _14181_/CLK _14181_/Q vdd gnd DFFPOSX1
XFILL_1__9716_ vdd gnd FILL
X_11393_ _11393_/A _11393_/B _11393_/Y vdd gnd NOR2X1
X_13132_ _13132_/A _13132_/B _13132_/Y vdd gnd NOR2X1
X_10344_ _10344_/A _10344_/Y vdd gnd INVX1
XFILL_1__9647_ vdd gnd FILL
X_13063_ _13063_/A _13063_/B _13063_/Y vdd gnd NAND2X1
X_10275_ _10275_/A _10275_/B _10275_/Y vdd gnd NOR2X1
XFILL_1__9578_ vdd gnd FILL
X_12014_ _12014_/A _12014_/Y vdd gnd INVX1
XFILL256950x7350 vdd gnd FILL
XFILL_2__7322_ vdd gnd FILL
XFILL_1__8529_ vdd gnd FILL
XFILL_2__7253_ vdd gnd FILL
XFILL_1__11040_ vdd gnd FILL
XFILL_0__11770_ vdd gnd FILL
X_13965_ _13965_/A _13965_/Y vdd gnd INVX1
XFILL_2__7184_ vdd gnd FILL
X_12916_ _12916_/A _12916_/B _12916_/C _12916_/Y vdd gnd NOR3X1
X_13896_ _13896_/A _13896_/B _13896_/Y vdd gnd OR2X2
XFILL_0__10652_ vdd gnd FILL
XFILL_1__12991_ vdd gnd FILL
X_12847_ _12847_/A _12847_/B _12847_/C _12847_/Y vdd gnd NAND3X1
XFILL_1__14730_ vdd gnd FILL
XFILL_1__11942_ vdd gnd FILL
XFILL_0__13371_ vdd gnd FILL
XFILL_0__10583_ vdd gnd FILL
X_12778_ _12778_/A _12778_/B _12778_/C _12778_/Y vdd gnd OAI21X1
XFILL_1__14661_ vdd gnd FILL
XFILL_0__12322_ vdd gnd FILL
XFILL256950x46950 vdd gnd FILL
XFILL_1__11873_ vdd gnd FILL
X_14517_ _14517_/D _14517_/CLK _14517_/Q vdd gnd DFFPOSX1
X_11729_ _11729_/A _11729_/B _11729_/Y vdd gnd NAND2X1
XFILL_1__13612_ vdd gnd FILL
XFILL_2__11074_ vdd gnd FILL
XFILL_1__10824_ vdd gnd FILL
XFILL_1__14592_ vdd gnd FILL
XFILL_0__12253_ vdd gnd FILL
X_14448_ _14448_/A _14448_/B _14448_/C _14448_/Y vdd gnd OAI21X1
XFILL_2__10025_ vdd gnd FILL
XFILL_1__13543_ vdd gnd FILL
XFILL_0__11204_ vdd gnd FILL
XFILL_0__12184_ vdd gnd FILL
XFILL_0__8771_ vdd gnd FILL
X_14379_ _14379_/A _14379_/B _14379_/Y vdd gnd OR2X2
XFILL_0__11135_ vdd gnd FILL
XFILL_1__10686_ vdd gnd FILL
XFILL_0__7722_ vdd gnd FILL
XFILL_1__12425_ vdd gnd FILL
XFILL_0__11066_ vdd gnd FILL
X_8000_ _8000_/A _8000_/B _8000_/Y vdd gnd NOR2X1
XFILL_0__7653_ vdd gnd FILL
XFILL_2__10927_ vdd gnd FILL
XFILL_2__13715_ vdd gnd FILL
XFILL_0__10017_ vdd gnd FILL
XFILL_1__12356_ vdd gnd FILL
XFILL_0__7584_ vdd gnd FILL
XFILL_1__11307_ vdd gnd FILL
XFILL_0__14825_ vdd gnd FILL
XFILL_2__13646_ vdd gnd FILL
XFILL_2__10858_ vdd gnd FILL
XFILL_1__12287_ vdd gnd FILL
XFILL_0__9323_ vdd gnd FILL
X_9951_ _9951_/A _9951_/Y vdd gnd INVX1
XFILL_1__14026_ vdd gnd FILL
XFILL_2__13577_ vdd gnd FILL
XFILL_1__11238_ vdd gnd FILL
XFILL_0__14756_ vdd gnd FILL
XFILL_0__9254_ vdd gnd FILL
X_8902_ _8902_/D _8902_/CLK _8902_/Q vdd gnd DFFPOSX1
XFILL_0__11968_ vdd gnd FILL
X_9882_ _9882_/A _9882_/B _9882_/C _9882_/Y vdd gnd OAI21X1
XFILL_0__13707_ vdd gnd FILL
XFILL_0__8205_ vdd gnd FILL
XFILL_0__10919_ vdd gnd FILL
XFILL_1__11169_ vdd gnd FILL
XFILL_0__14687_ vdd gnd FILL
XFILL_0__9185_ vdd gnd FILL
XFILL_0__11899_ vdd gnd FILL
X_8833_ _8833_/A _8833_/B _8833_/C _8833_/Y vdd gnd OAI21X1
XFILL_0__13638_ vdd gnd FILL
XFILL_0__8136_ vdd gnd FILL
X_8764_ _8764_/A _8764_/B _8764_/Y vdd gnd OR2X2
XFILL_0__13569_ vdd gnd FILL
X_7715_ _7715_/A _7715_/B _7715_/Y vdd gnd NAND2X1
XFILL_0__8067_ vdd gnd FILL
X_8695_ _8695_/A _8695_/B _8695_/C _8695_/Y vdd gnd OAI21X1
XFILL_1__14859_ vdd gnd FILL
XFILL_1__7900_ vdd gnd FILL
X_7646_ _7646_/A _7646_/B _7646_/Y vdd gnd OR2X2
XFILL_1__7831_ vdd gnd FILL
X_7577_ _7577_/A _7577_/B _7577_/C _7577_/Y vdd gnd NAND3X1
X_9316_ _9316_/A _9316_/B _9316_/Y vdd gnd NAND2X1
XFILL_0__8969_ vdd gnd FILL
XFILL_1__7762_ vdd gnd FILL
XFILL_1__9501_ vdd gnd FILL
X_9247_ _9247_/A _9247_/B _9247_/Y vdd gnd NAND2X1
XFILL_1__7693_ vdd gnd FILL
XFILL_1__9432_ vdd gnd FILL
X_9178_ _9178_/A _9178_/Y vdd gnd INVX1
X_10060_ _10060_/A _10060_/B _10060_/C _10060_/Y vdd gnd NOR3X1
X_8129_ _8129_/A _8129_/B _8129_/Y vdd gnd NAND2X1
XFILL_1__9363_ vdd gnd FILL
XFILL_1__8314_ vdd gnd FILL
XFILL_1__9294_ vdd gnd FILL
XFILL_1__8245_ vdd gnd FILL
X_10962_ _10962_/A _10962_/Y vdd gnd INVX2
X_13750_ _13750_/A _13750_/B _13750_/C _13750_/Y vdd gnd OAI21X1
XFILL_1__8176_ vdd gnd FILL
X_12701_ _12701_/A _12701_/B _12701_/Y vdd gnd NAND2X1
XFILL_1__7127_ vdd gnd FILL
X_10893_ _10893_/A _10893_/Y vdd gnd INVX1
X_13681_ _13681_/A _13681_/B _13681_/C _13681_/Y vdd gnd OAI21X1
XFILL257250x180150 vdd gnd FILL
X_12632_ _12632_/A _12632_/B _12632_/Y vdd gnd NAND2X1
XFILL_1_CLKBUF1_insert70 vdd gnd FILL
X_12563_ _12563_/D _12563_/CLK _12563_/Q vdd gnd DFFPOSX1
XFILL_1_CLKBUF1_insert81 vdd gnd FILL
XFILL_1_CLKBUF1_insert92 vdd gnd FILL
X_14302_ _14302_/A _14302_/B _14302_/C _14302_/Y vdd gnd NAND3X1
X_11514_ _11514_/A _11514_/B _11514_/C _11514_/Y vdd gnd OAI21X1
XFILL_2__9610_ vdd gnd FILL
X_12494_ _12494_/A _12494_/B _12494_/Y vdd gnd NAND2X1
X_14233_ _14233_/A _14233_/B _14233_/C _14233_/Y vdd gnd OAI21X1
X_11445_ _11445_/A _11445_/Y vdd gnd INVX1
XFILL_2__9541_ vdd gnd FILL
XFILL_1__10540_ vdd gnd FILL
X_14164_ _14164_/D _14164_/CLK _14164_/Q vdd gnd DFFPOSX1
X_11376_ _11376_/A _11376_/B _11376_/C _11376_/Y vdd gnd AOI21X1
XFILL_2__9472_ vdd gnd FILL
XFILL_1__10471_ vdd gnd FILL
X_13115_ _13115_/A _13115_/B _13115_/C _13115_/Y vdd gnd NOR3X1
X_10327_ _10327_/A _10327_/B _10327_/C _10327_/Y vdd gnd AOI21X1
X_14095_ _14095_/A _14095_/B _14095_/Y vdd gnd NOR2X1
XFILL_1__12210_ vdd gnd FILL
XFILL_1__13190_ vdd gnd FILL
XFILL_0__12940_ vdd gnd FILL
X_13046_ _13046_/A _13046_/Y vdd gnd INVX1
X_10258_ _10258_/A _10258_/B _10258_/C _10258_/Y vdd gnd AOI21X1
XFILL_2__14480_ vdd gnd FILL
XFILL_1__12141_ vdd gnd FILL
XFILL256950x21750 vdd gnd FILL
XFILL_0__12871_ vdd gnd FILL
XFILL_2__7305_ vdd gnd FILL
X_10189_ _10189_/A _10189_/B _10189_/C _10189_/D _10189_/Y vdd gnd AOI22X1
XFILL_0__14610_ vdd gnd FILL
XFILL_0__11822_ vdd gnd FILL
XFILL_1__12072_ vdd gnd FILL
XFILL_2__7236_ vdd gnd FILL
XFILL_1__11023_ vdd gnd FILL
XFILL_0__11753_ vdd gnd FILL
XFILL_2__12313_ vdd gnd FILL
X_13948_ _13948_/A _13948_/B _13948_/Y vdd gnd NAND2X1
XFILL_2__7167_ vdd gnd FILL
XFILL_2__13293_ vdd gnd FILL
XFILL_0__14472_ vdd gnd FILL
XFILL_2__12244_ vdd gnd FILL
X_13879_ _13879_/A _13879_/B _13879_/Y vdd gnd NAND2X1
XFILL_2__7098_ vdd gnd FILL
XFILL_0__13423_ vdd gnd FILL
XFILL_0__10635_ vdd gnd FILL
XFILL_1__12974_ vdd gnd FILL
XFILL_1__14713_ vdd gnd FILL
XFILL_1__11925_ vdd gnd FILL
XFILL_0__13354_ vdd gnd FILL
X_7500_ _7500_/A _7500_/B _7500_/C _7500_/Y vdd gnd NAND3X1
XFILL_0__10566_ vdd gnd FILL
XFILL_0__9941_ vdd gnd FILL
X_8480_ _8480_/A _8480_/B _8480_/Y vdd gnd NAND2X1
XFILL_1__14644_ vdd gnd FILL
XFILL_0__12305_ vdd gnd FILL
XFILL_1__11856_ vdd gnd FILL
XFILL_0__13285_ vdd gnd FILL
X_7431_ _7431_/A _7431_/B _7431_/C _7431_/Y vdd gnd OAI21X1
XFILL_0__10497_ vdd gnd FILL
XFILL_0__9872_ vdd gnd FILL
XFILL_1__10807_ vdd gnd FILL
XFILL_1__14575_ vdd gnd FILL
XFILL_0__12236_ vdd gnd FILL
XFILL_1__11787_ vdd gnd FILL
XFILL_0__8823_ vdd gnd FILL
X_7362_ _7362_/A _7362_/B _7362_/C _7362_/Y vdd gnd NAND3X1
XFILL_2__10008_ vdd gnd FILL
XFILL_2__9739_ vdd gnd FILL
XFILL_1__13526_ vdd gnd FILL
X_9101_ _9101_/A _9101_/B _9101_/Y vdd gnd NAND2X1
XFILL_0__12167_ vdd gnd FILL
XFILL_0__8754_ vdd gnd FILL
X_7293_ _7293_/A _7293_/Y vdd gnd INVX1
XFILL_0__11118_ vdd gnd FILL
XFILL_1__10669_ vdd gnd FILL
X_9032_ _9032_/A _9032_/B _9032_/C _9032_/Y vdd gnd OAI21X1
XFILL_0__7705_ vdd gnd FILL
XFILL_0__12098_ vdd gnd FILL
XFILL_0__8685_ vdd gnd FILL
XFILL_1__12408_ vdd gnd FILL
XFILL_0__11049_ vdd gnd FILL
XFILL_1__13388_ vdd gnd FILL
XFILL_0__7636_ vdd gnd FILL
XFILL_1__12339_ vdd gnd FILL
XFILL_0__7567_ vdd gnd FILL
XFILL_0__14808_ vdd gnd FILL
XFILL_0__9306_ vdd gnd FILL
XFILL_0__7498_ vdd gnd FILL
X_9934_ _9934_/A _9934_/B _9934_/S _9934_/Y vdd gnd MUX2X1
XFILL_1__14009_ vdd gnd FILL
XFILL_0__14739_ vdd gnd FILL
XFILL_1__8030_ vdd gnd FILL
XFILL_0__9237_ vdd gnd FILL
X_9865_ _9865_/A _9865_/B _9865_/C _9865_/Y vdd gnd OAI21X1
XFILL_0__9168_ vdd gnd FILL
X_8816_ _8816_/A _8816_/B _8816_/Y vdd gnd NAND2X1
X_9796_ _9796_/D _9796_/CLK _9796_/Q vdd gnd DFFPOSX1
XFILL_0__8119_ vdd gnd FILL
XFILL_0__9099_ vdd gnd FILL
X_8747_ _8747_/A _8747_/B _8747_/Y vdd gnd NAND2X1
XFILL_1__9981_ vdd gnd FILL
XFILL_1__8932_ vdd gnd FILL
X_8678_ _8678_/A _8678_/B _8678_/Y vdd gnd OR2X2
X_7629_ _7629_/A _7629_/B _7629_/Y vdd gnd NAND2X1
XFILL_1_CLKBUF1_insert103 vdd gnd FILL
XFILL_1__7814_ vdd gnd FILL
XFILL_1__8794_ vdd gnd FILL
X_11230_ _11230_/A _11230_/B _11230_/Y vdd gnd NAND2X1
XFILL_1__7745_ vdd gnd FILL
X_11161_ _11161_/A _11161_/B _11161_/Y vdd gnd NAND2X1
XFILL_1__7676_ vdd gnd FILL
X_10112_ _10112_/A _10112_/B _10112_/Y vdd gnd NAND2X1
X_11092_ _11092_/A _11092_/Y vdd gnd INVX1
XFILL_1__9415_ vdd gnd FILL
X_14920_ _14920_/A _14920_/Y vdd gnd BUFX2
X_10043_ _10043_/A _10043_/B _10043_/C _10043_/Y vdd gnd NAND3X1
XFILL_1__9346_ vdd gnd FILL
X_14851_ _14851_/A _14851_/B _14851_/C _14851_/Y vdd gnd AOI21X1
XFILL_1__9277_ vdd gnd FILL
X_13802_ _13802_/A _13802_/B _13802_/C _13802_/Y vdd gnd NAND3X1
X_14782_ _14782_/A _14782_/B _14782_/Y vdd gnd NOR2X1
XFILL_1__8228_ vdd gnd FILL
X_11994_ _11994_/A _11994_/B _11994_/C _11994_/Y vdd gnd NAND3X1
X_13733_ _13733_/A _13733_/B _13733_/C _13733_/Y vdd gnd OAI21X1
X_10945_ _10945_/A _10945_/B _10945_/C _10945_/Y vdd gnd OAI21X1
XFILL_1__8159_ vdd gnd FILL
X_13664_ _13664_/A _13664_/B _13664_/C _13664_/Y vdd gnd NAND3X1
X_10876_ _10876_/A _10876_/B _10876_/Y vdd gnd NAND2X1
XFILL_0__10420_ vdd gnd FILL
X_12615_ _12615_/D _12615_/CLK _12615_/Q vdd gnd DFFPOSX1
X_13595_ _13595_/A _13595_/B _13595_/C _13595_/Y vdd gnd OAI21X1
XFILL_1__11710_ vdd gnd FILL
XFILL_1__12690_ vdd gnd FILL
XFILL_0__10351_ vdd gnd FILL
X_12546_ _12546_/D _12546_/CLK _12546_/Q vdd gnd DFFPOSX1
XFILL_2__13980_ vdd gnd FILL
XFILL_0__10282_ vdd gnd FILL
XFILL_0__13070_ vdd gnd FILL
X_12477_ _12477_/A _12477_/B _12477_/C _12477_/Y vdd gnd OAI21X1
XFILL_0__12021_ vdd gnd FILL
XFILL_1__14360_ vdd gnd FILL
XFILL_2__12931_ vdd gnd FILL
XFILL_1__11572_ vdd gnd FILL
X_14216_ _14216_/A _14216_/Y vdd gnd INVX1
X_11428_ _11428_/A _11428_/B _11428_/Y vdd gnd NOR2X1
XFILL_2__9524_ vdd gnd FILL
XFILL_1__13311_ vdd gnd FILL
XFILL_1__10523_ vdd gnd FILL
XFILL_1__14291_ vdd gnd FILL
XFILL_2__12862_ vdd gnd FILL
X_11359_ _11359_/A _11359_/B _11359_/C _11359_/Y vdd gnd OAI21X1
X_14147_ _14147_/A _14147_/B _14147_/Y vdd gnd NAND2X1
XFILL_2__14601_ vdd gnd FILL
XCLKBUF1_insert102 CLKBUF1_insert102/A CLKBUF1_insert102/Y vdd gnd CLKBUF1
XFILL_2__9455_ vdd gnd FILL
XFILL_1__13242_ vdd gnd FILL
XFILL_1__10454_ vdd gnd FILL
XFILL_2__12793_ vdd gnd FILL
XFILL_0__13972_ vdd gnd FILL
XFILL_0__8470_ vdd gnd FILL
X_14078_ _14078_/A _14078_/B _14078_/Y vdd gnd NAND2X1
XFILL_1__13173_ vdd gnd FILL
XFILL_2__9386_ vdd gnd FILL
XFILL_0__12923_ vdd gnd FILL
XFILL_1__10385_ vdd gnd FILL
XFILL_0__7421_ vdd gnd FILL
X_13029_ _13029_/A _13029_/B _13029_/Y vdd gnd NAND2X1
XFILL_1__12124_ vdd gnd FILL
XFILL_2__14463_ vdd gnd FILL
XFILL_0__12854_ vdd gnd FILL
XFILL_0__7352_ vdd gnd FILL
X_7980_ _7980_/D _7980_/CLK _7980_/Q vdd gnd DFFPOSX1
XFILL_1__12055_ vdd gnd FILL
XFILL_0__11805_ vdd gnd FILL
XFILL256050x64950 vdd gnd FILL
XFILL_2__14394_ vdd gnd FILL
XFILL_0__12785_ vdd gnd FILL
XFILL_0__7283_ vdd gnd FILL
XFILL_1__11006_ vdd gnd FILL
XFILL_2__7219_ vdd gnd FILL
XFILL_0__9022_ vdd gnd FILL
XFILL_0__11736_ vdd gnd FILL
X_9650_ _9650_/A _9650_/B _9650_/Y vdd gnd NOR2X1
XFILL_0__14455_ vdd gnd FILL
X_8601_ _8601_/A _8601_/B _8601_/C _8601_/Y vdd gnd AOI21X1
X_9581_ _9581_/A _9581_/B _9581_/C _9581_/Y vdd gnd OAI21X1
XFILL_2__12227_ vdd gnd FILL
XFILL_0__13406_ vdd gnd FILL
XFILL_0__10618_ vdd gnd FILL
XFILL_0__14386_ vdd gnd FILL
XFILL_1__12957_ vdd gnd FILL
X_8532_ _8532_/A _8532_/B _8532_/Y vdd gnd NAND2X1
XFILL_0__11598_ vdd gnd FILL
XFILL_1_BUFX2_insert290 vdd gnd FILL
XCLKBUF1_insert50 CLKBUF1_insert50/A CLKBUF1_insert50/Y vdd gnd CLKBUF1
XCLKBUF1_insert61 CLKBUF1_insert61/A CLKBUF1_insert61/Y vdd gnd CLKBUF1
XFILL_2__12158_ vdd gnd FILL
XCLKBUF1_insert72 CLKBUF1_insert72/A CLKBUF1_insert72/Y vdd gnd CLKBUF1
XFILL_1__11908_ vdd gnd FILL
XFILL_0__13337_ vdd gnd FILL
XFILL_1__12888_ vdd gnd FILL
XCLKBUF1_insert83 CLKBUF1_insert83/A CLKBUF1_insert83/Y vdd gnd CLKBUF1
XFILL_0__10549_ vdd gnd FILL
XFILL_0__9924_ vdd gnd FILL
XCLKBUF1_insert94 CLKBUF1_insert94/A CLKBUF1_insert94/Y vdd gnd CLKBUF1
X_8463_ _8463_/A _8463_/B _8463_/Y vdd gnd OR2X2
XFILL_1__14627_ vdd gnd FILL
XFILL_2__12089_ vdd gnd FILL
XFILL_1__11839_ vdd gnd FILL
XFILL_0__13268_ vdd gnd FILL
X_7414_ _7414_/A _7414_/B _7414_/C _7414_/Y vdd gnd OAI21X1
XFILL_0__9855_ vdd gnd FILL
X_8394_ _8394_/A _8394_/B _8394_/Y vdd gnd NAND2X1
XFILL_0__12219_ vdd gnd FILL
XFILL_1__14558_ vdd gnd FILL
XFILL_0__13199_ vdd gnd FILL
XFILL_0__8806_ vdd gnd FILL
X_7345_ _7345_/A _7345_/B _7345_/C _7345_/Y vdd gnd OAI21X1
XFILL_1__13509_ vdd gnd FILL
XFILL_1__14489_ vdd gnd FILL
XFILL_1__7530_ vdd gnd FILL
XFILL_0__8737_ vdd gnd FILL
X_7276_ _7276_/A _7276_/B _7276_/C _7276_/Y vdd gnd AOI21X1
X_9015_ _9015_/A _9015_/B _9015_/C _9015_/Y vdd gnd NAND3X1
XFILL_1__7461_ vdd gnd FILL
XFILL_0__8668_ vdd gnd FILL
XFILL_1__9200_ vdd gnd FILL
XFILL_0__7619_ vdd gnd FILL
XFILL_1__7392_ vdd gnd FILL
XFILL_0__8599_ vdd gnd FILL
XFILL_1__9131_ vdd gnd FILL
XFILL_1__9062_ vdd gnd FILL
X_9917_ _9917_/A _9917_/B _9917_/Y vdd gnd NAND2X1
XFILL_1__8013_ vdd gnd FILL
X_9848_ _9848_/A _9848_/B _9848_/Y vdd gnd NOR2X1
X_10730_ _10730_/D _10730_/CLK _10730_/Q vdd gnd DFFPOSX1
X_9779_ _9779_/D _9779_/CLK _9779_/Q vdd gnd DFFPOSX1
X_10661_ _10661_/A _10661_/B _10661_/C _10661_/Y vdd gnd OAI21X1
XFILL_1__9964_ vdd gnd FILL
X_12400_ _12400_/A _12400_/B _12400_/C _12400_/Y vdd gnd OAI21X1
X_13380_ _13380_/A _13380_/Y vdd gnd INVX1
X_10592_ _10592_/A _10592_/Y vdd gnd INVX1
XFILL_1__9895_ vdd gnd FILL
X_12331_ _12331_/A _12331_/B _12331_/C _12331_/Y vdd gnd OAI21X1
X_12262_ _12262_/A _12262_/B _12262_/C _12262_/Y vdd gnd OAI21X1
XFILL_2__7570_ vdd gnd FILL
XFILL_1__8777_ vdd gnd FILL
X_14001_ _14001_/A _14001_/B _14001_/C _14001_/Y vdd gnd OAI21X1
X_11213_ _11213_/A _11213_/B _11213_/Y vdd gnd OR2X2
X_12193_ _12193_/A _12193_/B _12193_/C _12193_/Y vdd gnd NAND3X1
XFILL_1__7728_ vdd gnd FILL
X_11144_ _11144_/A _11144_/B _11144_/Y vdd gnd NAND2X1
XFILL_1__7659_ vdd gnd FILL
X_11075_ _11075_/A _11075_/B _11075_/C _11075_/Y vdd gnd NOR3X1
XFILL_1__10170_ vdd gnd FILL
X_14903_ _14903_/D _14903_/CLK _14903_/Q vdd gnd DFFPOSX1
X_10026_ _10026_/A _10026_/B _10026_/C _10026_/Y vdd gnd AOI21X1
XFILL_1__9329_ vdd gnd FILL
XFILL_2__8122_ vdd gnd FILL
X_14834_ _14834_/A _14834_/Y vdd gnd INVX1
XFILL_2__10411_ vdd gnd FILL
XFILL_2__8053_ vdd gnd FILL
XFILL_2__11391_ vdd gnd FILL
X_14765_ _14765_/A _14765_/B _14765_/Y vdd gnd OR2X2
X_11977_ _11977_/A _11977_/B _11977_/C _11977_/Y vdd gnd OAI21X1
XFILL_0__11521_ vdd gnd FILL
XFILL_1__13860_ vdd gnd FILL
X_13716_ _13716_/A _13716_/B _13716_/C _13716_/Y vdd gnd AOI21X1
X_10928_ _10928_/A _10928_/Y vdd gnd INVX2
X_14696_ _14696_/A _14696_/B _14696_/Y vdd gnd NAND2X1
XFILL_0__14240_ vdd gnd FILL
XFILL_1__12811_ vdd gnd FILL
XFILL_0__11452_ vdd gnd FILL
XFILL_1__13791_ vdd gnd FILL
X_13647_ _13647_/A _13647_/B _13647_/C _13647_/Y vdd gnd OAI21X1
XFILL_2__12012_ vdd gnd FILL
X_10859_ _10859_/A _10859_/Y vdd gnd INVX2
XFILL_2__8955_ vdd gnd FILL
XFILL_0__10403_ vdd gnd FILL
XFILL_1__12742_ vdd gnd FILL
XFILL_0_BUFX2_insert220 vdd gnd FILL
XFILL_0_BUFX2_insert231 vdd gnd FILL
XFILL_0__11383_ vdd gnd FILL
XFILL_0_BUFX2_insert242 vdd gnd FILL
XFILL_2__7906_ vdd gnd FILL
XFILL_0_BUFX2_insert253 vdd gnd FILL
X_13578_ _13578_/A _13578_/B _13578_/Y vdd gnd NAND2X1
XFILL_0__13122_ vdd gnd FILL
XFILL_0_BUFX2_insert264 vdd gnd FILL
XFILL_0__10334_ vdd gnd FILL
XFILL_1__12673_ vdd gnd FILL
XFILL256650x43350 vdd gnd FILL
XFILL_0_BUFX2_insert275 vdd gnd FILL
X_12529_ _12529_/A _12529_/B _12529_/C _12529_/Y vdd gnd OAI21X1
XFILL_0_BUFX2_insert286 vdd gnd FILL
XFILL_0_BUFX2_insert297 vdd gnd FILL
XFILL_2__7837_ vdd gnd FILL
XFILL_1__14412_ vdd gnd FILL
XFILL_2__13963_ vdd gnd FILL
XFILL_0__13053_ vdd gnd FILL
XFILL_0__10265_ vdd gnd FILL
XFILL_0__9640_ vdd gnd FILL
XFILL_0__12004_ vdd gnd FILL
XFILL_1__14343_ vdd gnd FILL
XFILL_2__7768_ vdd gnd FILL
XFILL_1__11555_ vdd gnd FILL
XFILL_2__13894_ vdd gnd FILL
XFILL_2_BUFX2_insert13 vdd gnd FILL
X_7130_ _7130_/A _7130_/Y vdd gnd INVX1
XFILL_0__10196_ vdd gnd FILL
XFILL_0__9571_ vdd gnd FILL
XFILL_1__10506_ vdd gnd FILL
XFILL_1__14274_ vdd gnd FILL
XFILL_2__12845_ vdd gnd FILL
XFILL_1__11486_ vdd gnd FILL
XFILL_0__8522_ vdd gnd FILL
XFILL_2__9438_ vdd gnd FILL
XFILL_1__13225_ vdd gnd FILL
XFILL_1__10437_ vdd gnd FILL
XFILL_0__13955_ vdd gnd FILL
XFILL_2__12776_ vdd gnd FILL
XFILL_0__8453_ vdd gnd FILL
.ends

