VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO phase_accumulator
  CLASS BLOCK ;
  FOREIGN phase_accumulator ;
  ORIGIN 6.000 6.000 ;
  SIZE 777.000 BY 735.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 765.300 686.700 774.300 722.700 ;
        RECT 0.600 684.300 774.300 686.700 ;
        RECT 765.300 614.700 774.300 684.300 ;
        RECT 0.600 612.300 774.300 614.700 ;
        RECT 765.300 542.700 774.300 612.300 ;
        RECT 0.600 540.300 774.300 542.700 ;
        RECT 765.300 470.700 774.300 540.300 ;
        RECT 0.600 468.300 774.300 470.700 ;
        RECT 765.300 398.700 774.300 468.300 ;
        RECT 0.600 396.300 774.300 398.700 ;
        RECT 765.300 326.700 774.300 396.300 ;
        RECT 0.600 324.300 774.300 326.700 ;
        RECT 765.300 254.700 774.300 324.300 ;
        RECT 0.600 252.300 774.300 254.700 ;
        RECT 765.300 182.700 774.300 252.300 ;
        RECT 0.600 180.300 774.300 182.700 ;
        RECT 765.300 110.700 774.300 180.300 ;
        RECT 0.600 108.300 774.300 110.700 ;
        RECT 765.300 38.700 774.300 108.300 ;
        RECT 0.600 36.300 774.300 38.700 ;
        RECT 765.300 0.300 774.300 36.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.300 720.300 764.400 722.700 ;
        RECT -9.300 650.700 -0.300 720.300 ;
        RECT -9.300 648.300 764.400 650.700 ;
        RECT -9.300 578.700 -0.300 648.300 ;
        RECT -9.300 576.300 764.400 578.700 ;
        RECT -9.300 506.700 -0.300 576.300 ;
        RECT -9.300 504.300 764.400 506.700 ;
        RECT -9.300 434.700 -0.300 504.300 ;
        RECT -9.300 432.300 764.400 434.700 ;
        RECT -9.300 362.700 -0.300 432.300 ;
        RECT -9.300 360.300 764.400 362.700 ;
        RECT -9.300 290.700 -0.300 360.300 ;
        RECT -9.300 288.300 764.400 290.700 ;
        RECT -9.300 218.700 -0.300 288.300 ;
        RECT -9.300 216.300 764.400 218.700 ;
        RECT -9.300 146.700 -0.300 216.300 ;
        RECT -9.300 144.300 764.400 146.700 ;
        RECT -9.300 74.700 -0.300 144.300 ;
        RECT -9.300 72.300 764.400 74.700 ;
        RECT -9.300 2.700 -0.300 72.300 ;
        RECT -9.300 0.300 764.400 2.700 ;
    END
  END vdd
  PIN Aout[1]
    PORT
      LAYER metal2 ;
        RECT 659.400 721.050 660.450 729.450 ;
        RECT 433.950 718.950 436.050 721.050 ;
        RECT 658.950 718.950 661.050 721.050 ;
        RECT 430.950 699.450 433.050 700.050 ;
        RECT 434.400 699.450 435.450 718.950 ;
        RECT 430.950 698.400 435.450 699.450 ;
        RECT 430.950 697.950 433.050 698.400 ;
      LAYER metal3 ;
        RECT 433.950 720.600 436.050 721.050 ;
        RECT 658.950 720.600 661.050 721.050 ;
        RECT 433.950 719.400 661.050 720.600 ;
        RECT 433.950 718.950 436.050 719.400 ;
        RECT 658.950 718.950 661.050 719.400 ;
    END
  END Aout[1]
  PIN Aout[0]
    PORT
      LAYER metal2 ;
        RECT 653.400 724.050 654.450 729.450 ;
        RECT 643.950 721.950 646.050 724.050 ;
        RECT 652.950 721.950 655.050 724.050 ;
        RECT 644.400 520.050 645.450 721.950 ;
        RECT 529.950 517.950 532.050 520.050 ;
        RECT 643.950 517.950 646.050 520.050 ;
        RECT 526.950 339.450 529.050 340.050 ;
        RECT 530.400 339.450 531.450 517.950 ;
        RECT 526.950 338.400 531.450 339.450 ;
        RECT 526.950 337.950 529.050 338.400 ;
      LAYER metal3 ;
        RECT 643.950 723.600 646.050 724.050 ;
        RECT 652.950 723.600 655.050 724.050 ;
        RECT 643.950 722.400 655.050 723.600 ;
        RECT 643.950 721.950 646.050 722.400 ;
        RECT 652.950 721.950 655.050 722.400 ;
        RECT 529.950 519.600 532.050 520.050 ;
        RECT 643.950 519.600 646.050 520.050 ;
        RECT 529.950 518.400 646.050 519.600 ;
        RECT 529.950 517.950 532.050 518.400 ;
        RECT 643.950 517.950 646.050 518.400 ;
    END
  END Aout[0]
  PIN En
    PORT
      LAYER metal2 ;
        RECT 187.950 481.950 190.050 484.050 ;
        RECT 188.400 405.450 189.450 481.950 ;
        RECT 185.400 404.400 189.450 405.450 ;
        RECT 1.950 349.950 4.050 352.050 ;
        RECT 2.400 322.050 3.450 349.950 ;
        RECT 185.400 322.050 186.450 404.400 ;
        RECT 361.950 382.950 364.050 385.050 ;
        RECT 376.950 382.950 379.050 385.050 ;
        RECT 362.400 322.050 363.450 382.950 ;
        RECT 1.950 319.950 4.050 322.050 ;
        RECT 151.950 319.950 154.050 322.050 ;
        RECT 184.950 319.950 187.050 322.050 ;
        RECT 361.950 319.950 364.050 322.050 ;
        RECT 152.400 313.050 153.450 319.950 ;
        RECT 151.950 310.950 154.050 313.050 ;
        RECT 362.400 196.050 363.450 319.950 ;
        RECT 337.950 193.950 340.050 196.050 ;
        RECT 361.950 193.950 364.050 196.050 ;
        RECT 376.950 193.950 379.050 196.050 ;
      LAYER metal3 ;
        RECT 361.950 384.600 364.050 385.050 ;
        RECT 376.950 384.600 379.050 385.050 ;
        RECT 361.950 383.400 379.050 384.600 ;
        RECT 361.950 382.950 364.050 383.400 ;
        RECT 376.950 382.950 379.050 383.400 ;
        RECT 1.950 351.600 4.050 352.050 ;
        RECT -3.600 350.400 4.050 351.600 ;
        RECT 1.950 349.950 4.050 350.400 ;
        RECT 1.950 321.600 4.050 322.050 ;
        RECT 151.950 321.600 154.050 322.050 ;
        RECT 184.950 321.600 187.050 322.050 ;
        RECT 361.950 321.600 364.050 322.050 ;
        RECT 1.950 320.400 364.050 321.600 ;
        RECT 1.950 319.950 4.050 320.400 ;
        RECT 151.950 319.950 154.050 320.400 ;
        RECT 184.950 319.950 187.050 320.400 ;
        RECT 361.950 319.950 364.050 320.400 ;
        RECT 337.950 195.600 340.050 196.050 ;
        RECT 361.950 195.600 364.050 196.050 ;
        RECT 376.950 195.600 379.050 196.050 ;
        RECT 337.950 194.400 379.050 195.600 ;
        RECT 337.950 193.950 340.050 194.400 ;
        RECT 361.950 193.950 364.050 194.400 ;
        RECT 376.950 193.950 379.050 194.400 ;
    END
  END En
  PIN FCW[19]
    PORT
      LAYER metal2 ;
        RECT 695.400 728.400 699.450 729.450 ;
        RECT 698.400 706.050 699.450 728.400 ;
        RECT 697.950 703.950 700.050 706.050 ;
        RECT 727.950 703.950 730.050 706.050 ;
        RECT 728.400 700.050 729.450 703.950 ;
        RECT 727.950 697.950 730.050 700.050 ;
        RECT 733.950 697.950 736.050 700.050 ;
      LAYER metal3 ;
        RECT 697.950 705.600 700.050 706.050 ;
        RECT 727.950 705.600 730.050 706.050 ;
        RECT 697.950 704.400 730.050 705.600 ;
        RECT 697.950 703.950 700.050 704.400 ;
        RECT 727.950 703.950 730.050 704.400 ;
        RECT 727.950 699.600 730.050 700.050 ;
        RECT 733.950 699.600 736.050 700.050 ;
        RECT 727.950 698.400 736.050 699.600 ;
        RECT 727.950 697.950 730.050 698.400 ;
        RECT 733.950 697.950 736.050 698.400 ;
    END
  END FCW[19]
  PIN FCW[18]
    PORT
      LAYER metal2 ;
        RECT 734.400 728.400 738.450 729.450 ;
        RECT 737.400 663.450 738.450 728.400 ;
        RECT 737.400 662.400 741.450 663.450 ;
        RECT 736.950 624.450 739.050 625.050 ;
        RECT 740.400 624.450 741.450 662.400 ;
        RECT 736.950 623.400 741.450 624.450 ;
        RECT 736.950 622.950 739.050 623.400 ;
        RECT 737.400 561.450 738.450 622.950 ;
        RECT 734.400 560.400 738.450 561.450 ;
        RECT 734.400 556.050 735.450 560.400 ;
        RECT 733.950 553.950 736.050 556.050 ;
        RECT 742.950 553.950 745.050 556.050 ;
      LAYER metal3 ;
        RECT 733.950 555.600 736.050 556.050 ;
        RECT 742.950 555.600 745.050 556.050 ;
        RECT 733.950 554.400 745.050 555.600 ;
        RECT 733.950 553.950 736.050 554.400 ;
        RECT 742.950 553.950 745.050 554.400 ;
    END
  END FCW[18]
  PIN FCW[17]
    PORT
      LAYER metal2 ;
        RECT 742.950 240.450 745.050 241.050 ;
        RECT 742.950 239.400 747.450 240.450 ;
        RECT 742.950 238.950 745.050 239.400 ;
        RECT 746.400 235.050 747.450 239.400 ;
        RECT 727.950 232.950 730.050 235.050 ;
        RECT 745.950 232.950 748.050 235.050 ;
        RECT 728.400 202.050 729.450 232.950 ;
        RECT 727.950 199.950 730.050 202.050 ;
      LAYER metal3 ;
        RECT 727.950 234.600 730.050 235.050 ;
        RECT 745.950 234.600 748.050 235.050 ;
        RECT 727.950 233.400 771.600 234.600 ;
        RECT 727.950 232.950 730.050 233.400 ;
        RECT 745.950 232.950 748.050 233.400 ;
    END
  END FCW[17]
  PIN FCW[16]
    PORT
      LAYER metal2 ;
        RECT 697.950 310.950 700.050 313.050 ;
        RECT 733.950 304.950 736.050 307.050 ;
      LAYER metal3 ;
        RECT 697.950 310.950 700.050 313.050 ;
        RECT 698.400 306.600 699.600 310.950 ;
        RECT 733.950 306.600 736.050 307.050 ;
        RECT 698.400 305.400 771.600 306.600 ;
        RECT 733.950 304.950 736.050 305.400 ;
    END
  END FCW[16]
  PIN FCW[15]
    PORT
      LAYER metal2 ;
        RECT 352.950 561.450 355.050 562.050 ;
        RECT 352.950 560.400 357.450 561.450 ;
        RECT 352.950 559.950 355.050 560.400 ;
        RECT 356.400 550.050 357.450 560.400 ;
        RECT 745.950 556.950 748.050 559.050 ;
        RECT 746.400 550.050 747.450 556.950 ;
        RECT 355.950 547.950 358.050 550.050 ;
        RECT 745.950 547.950 748.050 550.050 ;
        RECT 356.400 529.050 357.450 547.950 ;
        RECT 349.950 526.950 352.050 529.050 ;
        RECT 355.950 526.950 358.050 529.050 ;
      LAYER metal3 ;
        RECT 745.950 558.600 748.050 559.050 ;
        RECT 745.950 557.400 771.600 558.600 ;
        RECT 745.950 556.950 748.050 557.400 ;
        RECT 355.950 549.600 358.050 550.050 ;
        RECT 745.950 549.600 748.050 550.050 ;
        RECT 355.950 548.400 748.050 549.600 ;
        RECT 355.950 547.950 358.050 548.400 ;
        RECT 745.950 547.950 748.050 548.400 ;
        RECT 349.950 528.600 352.050 529.050 ;
        RECT 355.950 528.600 358.050 529.050 ;
        RECT 349.950 527.400 358.050 528.600 ;
        RECT 349.950 526.950 352.050 527.400 ;
        RECT 355.950 526.950 358.050 527.400 ;
    END
  END FCW[15]
  PIN FCW[14]
    PORT
      LAYER metal2 ;
        RECT 259.950 703.950 262.050 706.050 ;
        RECT 349.950 703.950 352.050 706.050 ;
        RECT 394.950 703.950 397.050 706.050 ;
        RECT 260.400 634.050 261.450 703.950 ;
        RECT 391.950 699.450 394.050 700.050 ;
        RECT 395.400 699.450 396.450 703.950 ;
        RECT 763.950 700.950 766.050 703.050 ;
        RECT 391.950 698.400 396.450 699.450 ;
        RECT 391.950 697.950 394.050 698.400 ;
        RECT 395.400 694.050 396.450 698.400 ;
        RECT 764.400 694.050 765.450 700.950 ;
        RECT 394.950 691.950 397.050 694.050 ;
        RECT 763.950 691.950 766.050 694.050 ;
        RECT 259.950 631.950 262.050 634.050 ;
      LAYER metal3 ;
        RECT 259.950 705.600 262.050 706.050 ;
        RECT 349.950 705.600 352.050 706.050 ;
        RECT 394.950 705.600 397.050 706.050 ;
        RECT 259.950 704.400 397.050 705.600 ;
        RECT 259.950 703.950 262.050 704.400 ;
        RECT 349.950 703.950 352.050 704.400 ;
        RECT 394.950 703.950 397.050 704.400 ;
        RECT 763.950 702.600 766.050 703.050 ;
        RECT 763.950 701.400 771.600 702.600 ;
        RECT 763.950 700.950 766.050 701.400 ;
        RECT 394.950 693.600 397.050 694.050 ;
        RECT 763.950 693.600 766.050 694.050 ;
        RECT 394.950 692.400 766.050 693.600 ;
        RECT 394.950 691.950 397.050 692.400 ;
        RECT 763.950 691.950 766.050 692.400 ;
    END
  END FCW[14]
  PIN FCW[13]
    PORT
      LAYER metal2 ;
        RECT 589.950 706.950 592.050 709.050 ;
        RECT 590.400 706.050 591.450 706.950 ;
        RECT 469.950 703.950 472.050 706.050 ;
        RECT 508.950 703.950 511.050 706.050 ;
        RECT 589.950 703.950 592.050 706.050 ;
        RECT 470.400 699.450 471.450 703.950 ;
        RECT 472.950 699.450 475.050 700.050 ;
        RECT 470.400 698.400 475.050 699.450 ;
        RECT 472.950 697.950 475.050 698.400 ;
        RECT 586.950 699.450 589.050 700.050 ;
        RECT 590.400 699.450 591.450 703.950 ;
        RECT 586.950 698.400 591.450 699.450 ;
        RECT 586.950 697.950 589.050 698.400 ;
      LAYER metal3 ;
        RECT 589.950 708.600 592.050 709.050 ;
        RECT 589.950 707.400 771.600 708.600 ;
        RECT 589.950 706.950 592.050 707.400 ;
        RECT 469.950 705.600 472.050 706.050 ;
        RECT 508.950 705.600 511.050 706.050 ;
        RECT 589.950 705.600 592.050 706.050 ;
        RECT 469.950 704.400 592.050 705.600 ;
        RECT 469.950 703.950 472.050 704.400 ;
        RECT 508.950 703.950 511.050 704.400 ;
        RECT 589.950 703.950 592.050 704.400 ;
    END
  END FCW[13]
  PIN FCW[12]
    PORT
      LAYER metal2 ;
        RECT 700.950 712.950 703.050 715.050 ;
        RECT 701.400 712.050 702.450 712.950 ;
        RECT 622.950 709.950 625.050 712.050 ;
        RECT 700.950 709.950 703.050 712.050 ;
        RECT 623.400 706.050 624.450 709.950 ;
        RECT 622.950 703.950 625.050 706.050 ;
        RECT 701.400 673.050 702.450 709.950 ;
        RECT 700.950 670.950 703.050 673.050 ;
      LAYER metal3 ;
        RECT 700.950 714.600 703.050 715.050 ;
        RECT 700.950 713.400 771.600 714.600 ;
        RECT 700.950 712.950 703.050 713.400 ;
        RECT 622.950 711.600 625.050 712.050 ;
        RECT 700.950 711.600 703.050 712.050 ;
        RECT 622.950 710.400 703.050 711.600 ;
        RECT 622.950 709.950 625.050 710.400 ;
        RECT 700.950 709.950 703.050 710.400 ;
    END
  END FCW[12]
  PIN FCW[11]
    PORT
      LAYER metal2 ;
        RECT 751.950 718.950 754.050 721.050 ;
        RECT 752.400 268.050 753.450 718.950 ;
        RECT 697.950 265.950 700.050 268.050 ;
        RECT 712.950 265.950 715.050 268.050 ;
        RECT 751.950 265.950 754.050 268.050 ;
        RECT 713.400 235.050 714.450 265.950 ;
        RECT 700.950 232.950 703.050 235.050 ;
        RECT 712.950 232.950 715.050 235.050 ;
      LAYER metal3 ;
        RECT 751.950 720.600 754.050 721.050 ;
        RECT 751.950 719.400 771.600 720.600 ;
        RECT 751.950 718.950 754.050 719.400 ;
        RECT 697.950 267.600 700.050 268.050 ;
        RECT 712.950 267.600 715.050 268.050 ;
        RECT 751.950 267.600 754.050 268.050 ;
        RECT 697.950 266.400 754.050 267.600 ;
        RECT 697.950 265.950 700.050 266.400 ;
        RECT 712.950 265.950 715.050 266.400 ;
        RECT 751.950 265.950 754.050 266.400 ;
        RECT 700.950 234.600 703.050 235.050 ;
        RECT 712.950 234.600 715.050 235.050 ;
        RECT 700.950 233.400 715.050 234.600 ;
        RECT 700.950 232.950 703.050 233.400 ;
        RECT 712.950 232.950 715.050 233.400 ;
    END
  END FCW[11]
  PIN FCW[10]
    PORT
      LAYER metal1 ;
        RECT 730.950 99.450 733.050 100.050 ;
        RECT 736.950 99.450 739.050 100.050 ;
        RECT 730.950 98.550 739.050 99.450 ;
        RECT 730.950 97.950 733.050 98.550 ;
        RECT 736.950 97.950 739.050 98.550 ;
      LAYER metal2 ;
        RECT 730.950 160.950 733.050 163.050 ;
        RECT 731.400 132.450 732.450 160.950 ;
        RECT 731.400 131.400 735.450 132.450 ;
        RECT 734.400 130.050 735.450 131.400 ;
        RECT 733.950 129.450 736.050 130.050 ;
        RECT 733.950 128.400 738.450 129.450 ;
        RECT 733.950 127.950 736.050 128.400 ;
        RECT 737.400 100.050 738.450 128.400 ;
        RECT 730.950 97.950 733.050 100.050 ;
        RECT 736.950 97.950 739.050 100.050 ;
        RECT 731.400 52.050 732.450 97.950 ;
        RECT 730.950 49.950 733.050 52.050 ;
        RECT 742.950 49.950 745.050 52.050 ;
        RECT 743.400 4.050 744.450 49.950 ;
        RECT 730.950 1.950 733.050 4.050 ;
        RECT 742.950 1.950 745.050 4.050 ;
        RECT 731.400 -3.600 732.450 1.950 ;
      LAYER metal3 ;
        RECT 730.950 51.600 733.050 52.050 ;
        RECT 742.950 51.600 745.050 52.050 ;
        RECT 730.950 50.400 745.050 51.600 ;
        RECT 730.950 49.950 733.050 50.400 ;
        RECT 742.950 49.950 745.050 50.400 ;
        RECT 730.950 3.600 733.050 4.050 ;
        RECT 742.950 3.600 745.050 4.050 ;
        RECT 730.950 2.400 745.050 3.600 ;
        RECT 730.950 1.950 733.050 2.400 ;
        RECT 742.950 1.950 745.050 2.400 ;
    END
  END FCW[10]
  PIN FCW[9]
    PORT
      LAYER metal2 ;
        RECT 571.950 28.950 574.050 31.050 ;
        RECT 658.950 28.950 661.050 31.050 ;
        RECT 572.400 25.050 573.450 28.950 ;
        RECT 659.400 28.050 660.450 28.950 ;
        RECT 658.950 25.950 661.050 28.050 ;
        RECT 502.950 22.950 505.050 25.050 ;
        RECT 571.950 22.950 574.050 25.050 ;
        RECT 572.400 4.050 573.450 22.950 ;
        RECT 583.950 16.950 586.050 19.050 ;
        RECT 584.400 4.050 585.450 16.950 ;
        RECT 571.950 1.950 574.050 4.050 ;
        RECT 583.950 1.950 586.050 4.050 ;
        RECT 572.400 -3.600 573.450 1.950 ;
      LAYER metal3 ;
        RECT 571.950 30.600 574.050 31.050 ;
        RECT 658.950 30.600 661.050 31.050 ;
        RECT 571.950 29.400 661.050 30.600 ;
        RECT 571.950 28.950 574.050 29.400 ;
        RECT 658.950 28.950 661.050 29.400 ;
        RECT 502.950 24.600 505.050 25.050 ;
        RECT 571.950 24.600 574.050 25.050 ;
        RECT 502.950 23.400 574.050 24.600 ;
        RECT 502.950 22.950 505.050 23.400 ;
        RECT 571.950 22.950 574.050 23.400 ;
        RECT 571.950 3.600 574.050 4.050 ;
        RECT 583.950 3.600 586.050 4.050 ;
        RECT 571.950 2.400 586.050 3.600 ;
        RECT 571.950 1.950 574.050 2.400 ;
        RECT 583.950 1.950 586.050 2.400 ;
    END
  END FCW[9]
  PIN FCW[8]
    PORT
      LAYER metal2 ;
        RECT 421.950 55.950 424.050 58.050 ;
        RECT 439.950 55.950 442.050 58.050 ;
        RECT 440.400 52.050 441.450 55.950 ;
        RECT 439.950 49.950 442.050 52.050 ;
        RECT 448.950 49.950 451.050 52.050 ;
        RECT 460.950 49.950 463.050 52.050 ;
        RECT 449.400 -3.600 450.450 49.950 ;
      LAYER metal3 ;
        RECT 421.950 57.600 424.050 58.050 ;
        RECT 439.950 57.600 442.050 58.050 ;
        RECT 421.950 56.400 442.050 57.600 ;
        RECT 421.950 55.950 424.050 56.400 ;
        RECT 439.950 55.950 442.050 56.400 ;
        RECT 439.950 51.600 442.050 52.050 ;
        RECT 448.950 51.600 451.050 52.050 ;
        RECT 460.950 51.600 463.050 52.050 ;
        RECT 439.950 50.400 463.050 51.600 ;
        RECT 439.950 49.950 442.050 50.400 ;
        RECT 448.950 49.950 451.050 50.400 ;
        RECT 460.950 49.950 463.050 50.400 ;
    END
  END FCW[8]
  PIN FCW[7]
    PORT
      LAYER metal2 ;
        RECT 226.950 57.450 229.050 58.050 ;
        RECT 224.400 56.400 229.050 57.450 ;
        RECT 224.400 25.050 225.450 56.400 ;
        RECT 226.950 55.950 229.050 56.400 ;
        RECT 121.950 22.950 124.050 25.050 ;
        RECT 151.950 22.950 154.050 25.050 ;
        RECT 187.950 22.950 190.050 25.050 ;
        RECT 223.950 22.950 226.050 25.050 ;
        RECT 122.400 19.050 123.450 22.950 ;
        RECT 73.950 16.950 76.050 19.050 ;
        RECT 121.950 16.950 124.050 19.050 ;
        RECT 74.400 -3.600 75.450 16.950 ;
      LAYER metal3 ;
        RECT 121.950 24.600 124.050 25.050 ;
        RECT 151.950 24.600 154.050 25.050 ;
        RECT 187.950 24.600 190.050 25.050 ;
        RECT 223.950 24.600 226.050 25.050 ;
        RECT 121.950 23.400 226.050 24.600 ;
        RECT 121.950 22.950 124.050 23.400 ;
        RECT 151.950 22.950 154.050 23.400 ;
        RECT 187.950 22.950 190.050 23.400 ;
        RECT 223.950 22.950 226.050 23.400 ;
        RECT 73.950 18.600 76.050 19.050 ;
        RECT 121.950 18.600 124.050 19.050 ;
        RECT 73.950 17.400 124.050 18.600 ;
        RECT 73.950 16.950 76.050 17.400 ;
        RECT 121.950 16.950 124.050 17.400 ;
    END
  END FCW[7]
  PIN FCW[6]
    PORT
      LAYER metal2 ;
        RECT 109.950 49.950 112.050 52.050 ;
        RECT 31.950 16.950 34.050 19.050 ;
        RECT 32.400 16.050 33.450 16.950 ;
        RECT 110.400 16.050 111.450 49.950 ;
        RECT 31.950 13.950 34.050 16.050 ;
        RECT 109.950 13.950 112.050 16.050 ;
        RECT 32.400 -2.550 33.450 13.950 ;
        RECT 32.400 -3.600 36.450 -2.550 ;
      LAYER metal3 ;
        RECT 31.950 15.600 34.050 16.050 ;
        RECT 109.950 15.600 112.050 16.050 ;
        RECT 31.950 14.400 112.050 15.600 ;
        RECT 31.950 13.950 34.050 14.400 ;
        RECT 109.950 13.950 112.050 14.400 ;
    END
  END FCW[6]
  PIN FCW[5]
    PORT
      LAYER metal2 ;
        RECT 31.950 88.950 34.050 91.050 ;
        RECT 32.400 57.450 33.450 88.950 ;
        RECT 29.400 56.400 33.450 57.450 ;
        RECT 29.400 51.450 30.450 56.400 ;
        RECT 31.950 51.450 34.050 52.050 ;
        RECT 29.400 50.400 34.050 51.450 ;
        RECT 29.400 -3.600 30.450 50.400 ;
        RECT 31.950 49.950 34.050 50.400 ;
    END
  END FCW[5]
  PIN FCW[4]
    PORT
      LAYER metal2 ;
        RECT 28.950 193.950 31.050 196.050 ;
        RECT 29.400 163.050 30.450 193.950 ;
        RECT 22.950 160.950 25.050 163.050 ;
        RECT 28.950 160.950 31.050 163.050 ;
        RECT 34.950 160.950 37.050 163.050 ;
        RECT 23.400 -3.600 24.450 160.950 ;
      LAYER metal3 ;
        RECT 22.950 162.600 25.050 163.050 ;
        RECT 28.950 162.600 31.050 163.050 ;
        RECT 34.950 162.600 37.050 163.050 ;
        RECT 22.950 161.400 37.050 162.600 ;
        RECT 22.950 160.950 25.050 161.400 ;
        RECT 28.950 160.950 31.050 161.400 ;
        RECT 34.950 160.950 37.050 161.400 ;
    END
  END FCW[4]
  PIN FCW[3]
    PORT
      LAYER metal2 ;
        RECT 4.950 679.950 7.050 682.050 ;
        RECT 5.400 490.050 6.450 679.950 ;
        RECT 4.950 487.950 7.050 490.050 ;
        RECT 31.950 489.450 34.050 490.050 ;
        RECT 34.950 489.450 37.050 490.050 ;
        RECT 31.950 488.400 37.050 489.450 ;
        RECT 31.950 487.950 34.050 488.400 ;
        RECT 34.950 487.950 37.050 488.400 ;
        RECT 32.400 462.450 33.450 487.950 ;
        RECT 32.400 461.400 36.450 462.450 ;
        RECT 35.400 457.050 36.450 461.400 ;
        RECT 34.950 454.950 37.050 457.050 ;
      LAYER metal3 ;
        RECT 4.950 681.600 7.050 682.050 ;
        RECT -3.600 680.400 7.050 681.600 ;
        RECT 4.950 679.950 7.050 680.400 ;
        RECT 4.950 489.600 7.050 490.050 ;
        RECT 31.950 489.600 34.050 490.050 ;
        RECT 4.950 488.400 34.050 489.600 ;
        RECT 4.950 487.950 7.050 488.400 ;
        RECT 31.950 487.950 34.050 488.400 ;
    END
  END FCW[3]
  PIN FCW[2]
    PORT
      LAYER metal2 ;
        RECT 1.950 673.950 4.050 676.050 ;
        RECT 2.400 601.050 3.450 673.950 ;
        RECT 1.950 598.950 4.050 601.050 ;
        RECT 31.950 598.950 34.050 601.050 ;
        RECT 34.950 595.950 37.050 598.050 ;
        RECT 35.400 562.050 36.450 595.950 ;
        RECT 34.950 559.950 37.050 562.050 ;
      LAYER metal3 ;
        RECT 1.950 675.600 4.050 676.050 ;
        RECT -3.600 674.400 4.050 675.600 ;
        RECT 1.950 673.950 4.050 674.400 ;
        RECT 1.950 600.600 4.050 601.050 ;
        RECT 31.950 600.600 34.050 601.050 ;
        RECT 1.950 599.400 34.050 600.600 ;
        RECT 1.950 598.950 4.050 599.400 ;
        RECT 31.950 598.950 34.050 599.400 ;
        RECT 32.400 597.600 33.600 598.950 ;
        RECT 34.950 597.600 37.050 598.050 ;
        RECT 32.400 596.400 37.050 597.600 ;
        RECT 34.950 595.950 37.050 596.400 ;
    END
  END FCW[2]
  PIN FCW[1]
    PORT
      LAYER metal2 ;
        RECT 31.950 697.950 34.050 700.050 ;
        RECT 32.400 697.050 33.450 697.950 ;
        RECT 25.950 694.950 28.050 697.050 ;
        RECT 31.950 694.950 34.050 697.050 ;
        RECT 26.400 667.050 27.450 694.950 ;
        RECT 25.950 664.950 28.050 667.050 ;
        RECT 28.950 664.950 31.050 667.050 ;
      LAYER metal3 ;
        RECT 25.950 696.600 28.050 697.050 ;
        RECT 31.950 696.600 34.050 697.050 ;
        RECT 25.950 695.400 34.050 696.600 ;
        RECT 25.950 694.950 28.050 695.400 ;
        RECT 31.950 694.950 34.050 695.400 ;
        RECT -3.600 666.600 -2.400 669.600 ;
        RECT 25.950 666.600 28.050 667.050 ;
        RECT 28.950 666.600 31.050 667.050 ;
        RECT -3.600 665.400 31.050 666.600 ;
        RECT 25.950 664.950 28.050 665.400 ;
        RECT 28.950 664.950 31.050 665.400 ;
    END
  END FCW[1]
  PIN FCW[0]
    PORT
      LAYER metal2 ;
        RECT 109.950 631.950 112.050 634.050 ;
        RECT 178.950 631.950 181.050 634.050 ;
      LAYER metal3 ;
        RECT 109.950 633.600 112.050 634.050 ;
        RECT 178.950 633.600 181.050 634.050 ;
        RECT -3.600 632.400 181.050 633.600 ;
        RECT -3.600 629.400 -2.400 632.400 ;
        RECT 109.950 631.950 112.050 632.400 ;
        RECT 178.950 631.950 181.050 632.400 ;
    END
  END FCW[0]
  PIN ISout
    PORT
      LAYER metal2 ;
        RECT 647.400 700.050 648.450 729.450 ;
        RECT 646.950 697.950 649.050 700.050 ;
        RECT 658.950 697.950 661.050 700.050 ;
      LAYER metal3 ;
        RECT 646.950 699.600 649.050 700.050 ;
        RECT 658.950 699.600 661.050 700.050 ;
        RECT 646.950 698.400 661.050 699.600 ;
        RECT 646.950 697.950 649.050 698.400 ;
        RECT 658.950 697.950 661.050 698.400 ;
    END
  END ISout
  PIN Vld
    PORT
      LAYER metal2 ;
        RECT 308.400 699.450 309.450 729.450 ;
        RECT 310.950 699.450 313.050 700.050 ;
        RECT 308.400 698.400 313.050 699.450 ;
        RECT 310.950 697.950 313.050 698.400 ;
    END
  END Vld
  PIN clk
    PORT
      LAYER metal2 ;
        RECT 193.950 558.450 196.050 559.050 ;
        RECT 292.950 558.450 295.050 559.050 ;
        RECT 193.950 557.400 198.450 558.450 ;
        RECT 193.950 556.950 196.050 557.400 ;
        RECT 197.400 553.050 198.450 557.400 ;
        RECT 290.400 557.400 295.050 558.450 ;
        RECT 290.400 553.050 291.450 557.400 ;
        RECT 292.950 556.950 295.050 557.400 ;
        RECT 196.950 550.950 199.050 553.050 ;
        RECT 289.950 550.950 292.050 553.050 ;
        RECT 197.400 454.050 198.450 550.950 ;
        RECT 190.950 451.950 193.050 454.050 ;
        RECT 196.950 451.950 199.050 454.050 ;
        RECT 197.400 349.050 198.450 451.950 ;
        RECT 28.950 346.950 31.050 349.050 ;
        RECT 196.950 346.950 199.050 349.050 ;
        RECT 292.950 346.950 295.050 349.050 ;
        RECT 29.400 346.050 30.450 346.950 ;
        RECT 28.950 343.950 31.050 346.050 ;
        RECT 29.400 343.050 30.450 343.950 ;
        RECT 28.950 340.950 31.050 343.050 ;
        RECT 293.400 238.050 294.450 346.950 ;
        RECT 289.950 237.450 292.050 238.050 ;
        RECT 292.950 237.450 295.050 238.050 ;
        RECT 289.950 236.400 295.050 237.450 ;
        RECT 289.950 235.950 292.050 236.400 ;
        RECT 292.950 235.950 295.050 236.400 ;
        RECT 325.950 235.950 328.050 238.050 ;
      LAYER metal3 ;
        RECT 196.950 552.600 199.050 553.050 ;
        RECT 289.950 552.600 292.050 553.050 ;
        RECT 196.950 551.400 292.050 552.600 ;
        RECT 196.950 550.950 199.050 551.400 ;
        RECT 289.950 550.950 292.050 551.400 ;
        RECT 190.950 453.600 193.050 454.050 ;
        RECT 196.950 453.600 199.050 454.050 ;
        RECT 190.950 452.400 199.050 453.600 ;
        RECT 190.950 451.950 193.050 452.400 ;
        RECT 196.950 451.950 199.050 452.400 ;
        RECT 28.950 348.600 31.050 349.050 ;
        RECT 196.950 348.600 199.050 349.050 ;
        RECT 292.950 348.600 295.050 349.050 ;
        RECT 28.950 347.400 295.050 348.600 ;
        RECT 28.950 346.950 31.050 347.400 ;
        RECT 196.950 346.950 199.050 347.400 ;
        RECT 292.950 346.950 295.050 347.400 ;
        RECT 28.950 345.600 31.050 346.050 ;
        RECT -3.600 344.400 31.050 345.600 ;
        RECT 28.950 343.950 31.050 344.400 ;
        RECT 292.950 237.600 295.050 238.050 ;
        RECT 325.950 237.600 328.050 238.050 ;
        RECT 292.950 236.400 328.050 237.600 ;
        RECT 292.950 235.950 295.050 236.400 ;
        RECT 325.950 235.950 328.050 236.400 ;
    END
  END clk
  OBS
      LAYER metal1 ;
        RECT 33.450 707.400 35.250 719.250 ;
        RECT 37.650 707.400 39.450 719.250 ;
        RECT 71.400 713.400 73.200 719.250 ;
        RECT 74.700 707.400 76.500 719.250 ;
        RECT 78.900 707.400 80.700 719.250 ;
        RECT 110.550 713.400 112.350 719.250 ;
        RECT 113.550 713.400 115.350 719.250 ;
        RECT 146.550 713.400 148.350 719.250 ;
        RECT 149.550 713.400 151.350 719.250 ;
        RECT 152.550 713.400 154.350 719.250 ;
        RECT 33.450 706.350 36.000 707.400 ;
        RECT 32.100 702.150 33.900 703.950 ;
        RECT 31.950 700.050 34.050 702.150 ;
        RECT 34.950 699.150 36.000 706.350 ;
        RECT 71.250 705.150 73.050 706.950 ;
        RECT 38.100 702.150 39.900 703.950 ;
        RECT 70.950 703.050 73.050 705.150 ;
        RECT 74.850 702.150 76.050 707.400 ;
        RECT 80.100 702.150 81.900 703.950 ;
        RECT 37.950 700.050 40.050 702.150 ;
        RECT 73.950 700.050 76.050 702.150 ;
        RECT 34.950 697.050 37.050 699.150 ;
        RECT 34.950 690.600 36.000 697.050 ;
        RECT 73.950 696.750 75.150 700.050 ;
        RECT 76.950 698.850 79.050 700.950 ;
        RECT 79.950 700.050 82.050 702.150 ;
        RECT 113.400 700.950 114.600 713.400 ;
        RECT 149.550 705.150 150.750 713.400 ;
        RECT 186.300 707.400 188.100 719.250 ;
        RECT 190.500 707.400 192.300 719.250 ;
        RECT 193.800 713.400 195.600 719.250 ;
        RECT 224.550 708.300 226.350 719.250 ;
        RECT 227.550 709.200 229.350 719.250 ;
        RECT 230.550 708.300 232.350 719.250 ;
        RECT 224.550 707.400 232.350 708.300 ;
        RECT 233.550 707.400 235.350 719.250 ;
        RECT 267.300 707.400 269.100 719.250 ;
        RECT 271.500 707.400 273.300 719.250 ;
        RECT 274.800 713.400 276.600 719.250 ;
        RECT 305.550 713.400 307.350 719.250 ;
        RECT 145.950 701.850 148.050 703.950 ;
        RECT 148.950 703.050 151.050 705.150 ;
        RECT 110.100 699.150 111.900 700.950 ;
        RECT 77.100 697.050 78.900 698.850 ;
        RECT 109.950 697.050 112.050 699.150 ;
        RECT 112.950 698.850 115.050 700.950 ;
        RECT 146.100 700.050 147.900 701.850 ;
        RECT 71.250 695.700 75.000 696.750 ;
        RECT 71.250 693.600 72.450 695.700 ;
        RECT 31.650 687.750 33.450 690.600 ;
        RECT 34.650 687.750 36.450 690.600 ;
        RECT 37.650 687.750 39.450 690.600 ;
        RECT 70.650 687.750 72.450 693.600 ;
        RECT 73.650 692.700 81.450 694.050 ;
        RECT 73.650 687.750 75.450 692.700 ;
        RECT 76.650 687.750 78.450 691.800 ;
        RECT 79.650 687.750 81.450 692.700 ;
        RECT 113.400 690.600 114.600 698.850 ;
        RECT 149.550 695.700 150.750 703.050 ;
        RECT 151.950 701.850 154.050 703.950 ;
        RECT 185.100 702.150 186.900 703.950 ;
        RECT 190.950 702.150 192.150 707.400 ;
        RECT 193.950 705.150 195.750 706.950 ;
        RECT 193.950 703.050 196.050 705.150 ;
        RECT 196.950 702.450 199.050 703.050 ;
        RECT 202.950 702.450 205.050 703.050 ;
        RECT 152.100 700.050 153.900 701.850 ;
        RECT 184.950 700.050 187.050 702.150 ;
        RECT 187.950 698.850 190.050 700.950 ;
        RECT 190.950 700.050 193.050 702.150 ;
        RECT 196.950 701.550 205.050 702.450 ;
        RECT 233.700 702.150 234.900 707.400 ;
        RECT 266.100 702.150 267.900 703.950 ;
        RECT 271.950 702.150 273.150 707.400 ;
        RECT 274.950 705.150 276.750 706.950 ;
        RECT 305.550 706.500 306.750 713.400 ;
        RECT 308.850 707.400 310.650 719.250 ;
        RECT 311.850 707.400 313.650 719.250 ;
        RECT 344.550 713.400 346.350 719.250 ;
        RECT 347.550 713.400 349.350 719.250 ;
        RECT 305.550 705.600 311.250 706.500 ;
        RECT 274.950 703.050 277.050 705.150 ;
        RECT 309.000 704.700 311.250 705.600 ;
        RECT 305.100 702.150 306.900 703.950 ;
        RECT 196.950 700.950 199.050 701.550 ;
        RECT 202.950 700.950 205.050 701.550 ;
        RECT 188.100 697.050 189.900 698.850 ;
        RECT 191.850 696.750 193.050 700.050 ;
        RECT 193.950 699.450 196.050 700.050 ;
        RECT 220.950 699.450 223.050 700.050 ;
        RECT 193.950 698.550 223.050 699.450 ;
        RECT 223.950 698.850 226.050 700.950 ;
        RECT 227.100 699.150 228.900 700.950 ;
        RECT 193.950 697.950 196.050 698.550 ;
        RECT 220.950 697.950 223.050 698.550 ;
        RECT 224.100 697.050 225.900 698.850 ;
        RECT 226.950 697.050 229.050 699.150 ;
        RECT 229.950 698.850 232.050 700.950 ;
        RECT 232.950 700.050 235.050 702.150 ;
        RECT 265.950 700.050 268.050 702.150 ;
        RECT 230.100 697.050 231.900 698.850 ;
        RECT 192.000 695.700 195.750 696.750 ;
        RECT 149.550 694.800 153.150 695.700 ;
        RECT 110.550 687.750 112.350 690.600 ;
        RECT 113.550 687.750 115.350 690.600 ;
        RECT 146.850 687.750 148.650 693.600 ;
        RECT 151.350 687.750 153.150 694.800 ;
        RECT 185.550 692.700 193.350 694.050 ;
        RECT 185.550 687.750 187.350 692.700 ;
        RECT 188.550 687.750 190.350 691.800 ;
        RECT 191.550 687.750 193.350 692.700 ;
        RECT 194.550 693.600 195.750 695.700 ;
        RECT 233.700 693.600 234.900 700.050 ;
        RECT 268.950 698.850 271.050 700.950 ;
        RECT 271.950 700.050 274.050 702.150 ;
        RECT 304.950 700.050 307.050 702.150 ;
        RECT 269.100 697.050 270.900 698.850 ;
        RECT 272.850 696.750 274.050 700.050 ;
        RECT 273.000 695.700 276.750 696.750 ;
        RECT 194.550 687.750 196.350 693.600 ;
        RECT 225.000 687.750 226.800 693.600 ;
        RECT 229.200 691.950 234.900 693.600 ;
        RECT 266.550 692.700 274.350 694.050 ;
        RECT 229.200 687.750 231.000 691.950 ;
        RECT 232.500 687.750 234.300 690.600 ;
        RECT 266.550 687.750 268.350 692.700 ;
        RECT 269.550 687.750 271.350 691.800 ;
        RECT 272.550 687.750 274.350 692.700 ;
        RECT 275.550 693.600 276.750 695.700 ;
        RECT 309.000 696.300 310.050 704.700 ;
        RECT 312.150 702.150 313.350 707.400 ;
        RECT 344.100 702.150 345.900 703.950 ;
        RECT 310.950 700.050 313.350 702.150 ;
        RECT 343.950 700.050 346.050 702.150 ;
        RECT 309.000 695.400 311.250 696.300 ;
        RECT 306.150 694.500 311.250 695.400 ;
        RECT 275.550 687.750 277.350 693.600 ;
        RECT 306.150 690.600 307.350 694.500 ;
        RECT 312.150 693.600 313.350 700.050 ;
        RECT 347.700 696.300 348.900 713.400 ;
        RECT 351.150 707.400 352.950 719.250 ;
        RECT 354.150 707.400 355.950 719.250 ;
        RECT 386.550 707.400 388.350 719.250 ;
        RECT 390.750 707.400 392.550 719.250 ;
        RECT 349.950 701.850 352.050 703.950 ;
        RECT 354.150 702.150 355.350 707.400 ;
        RECT 390.000 706.350 392.550 707.400 ;
        RECT 425.550 713.400 427.350 719.250 ;
        RECT 425.550 706.500 426.750 713.400 ;
        RECT 428.850 707.400 430.650 719.250 ;
        RECT 431.850 707.400 433.650 719.250 ;
        RECT 468.150 708.900 469.950 719.250 ;
        RECT 467.550 707.550 469.950 708.900 ;
        RECT 471.150 707.550 472.950 719.250 ;
        RECT 386.100 702.150 387.900 703.950 ;
        RECT 350.100 700.050 351.900 701.850 ;
        RECT 352.950 700.050 355.350 702.150 ;
        RECT 385.950 700.050 388.050 702.150 ;
        RECT 344.550 695.100 352.050 696.300 ;
        RECT 305.550 687.750 307.350 690.600 ;
        RECT 308.850 687.750 310.650 693.600 ;
        RECT 311.850 687.750 313.650 693.600 ;
        RECT 344.550 687.750 346.350 695.100 ;
        RECT 350.250 694.500 352.050 695.100 ;
        RECT 354.150 693.600 355.350 700.050 ;
        RECT 390.000 699.150 391.050 706.350 ;
        RECT 425.550 705.600 431.250 706.500 ;
        RECT 429.000 704.700 431.250 705.600 ;
        RECT 392.100 702.150 393.900 703.950 ;
        RECT 425.100 702.150 426.900 703.950 ;
        RECT 391.950 700.050 394.050 702.150 ;
        RECT 424.950 700.050 427.050 702.150 ;
        RECT 388.950 697.050 391.050 699.150 ;
        RECT 349.050 687.750 350.850 693.600 ;
        RECT 352.050 692.100 355.350 693.600 ;
        RECT 352.050 687.750 353.850 692.100 ;
        RECT 390.000 690.600 391.050 697.050 ;
        RECT 429.000 696.300 430.050 704.700 ;
        RECT 432.150 702.150 433.350 707.400 ;
        RECT 430.950 700.050 433.350 702.150 ;
        RECT 467.550 700.950 468.900 707.550 ;
        RECT 475.650 707.400 477.450 719.250 ;
        RECT 503.550 713.400 505.350 719.250 ;
        RECT 506.550 713.400 508.350 719.250 ;
        RECT 509.550 713.400 511.350 719.250 ;
        RECT 542.400 713.400 544.200 719.250 ;
        RECT 470.250 706.200 472.050 706.650 ;
        RECT 476.250 706.200 477.450 707.400 ;
        RECT 470.250 705.000 477.450 706.200 ;
        RECT 506.550 705.150 507.750 713.400 ;
        RECT 545.700 707.400 547.500 719.250 ;
        RECT 549.900 707.400 551.700 719.250 ;
        RECT 581.550 707.400 583.350 719.250 ;
        RECT 585.750 707.400 587.550 719.250 ;
        RECT 617.550 713.400 619.350 719.250 ;
        RECT 620.550 713.400 622.350 719.250 ;
        RECT 623.550 713.400 625.350 719.250 ;
        RECT 542.250 705.150 544.050 706.950 ;
        RECT 470.250 704.850 472.050 705.000 ;
        RECT 429.000 695.400 431.250 696.300 ;
        RECT 426.150 694.500 431.250 695.400 ;
        RECT 426.150 690.600 427.350 694.500 ;
        RECT 432.150 693.600 433.350 700.050 ;
        RECT 466.950 698.850 469.050 700.950 ;
        RECT 466.950 693.600 468.000 698.850 ;
        RECT 470.400 696.600 471.300 704.850 ;
        RECT 473.100 702.150 474.900 703.950 ;
        RECT 472.950 700.050 475.050 702.150 ;
        RECT 502.950 701.850 505.050 703.950 ;
        RECT 505.950 703.050 508.050 705.150 ;
        RECT 476.100 699.150 477.900 700.950 ;
        RECT 503.100 700.050 504.900 701.850 ;
        RECT 475.950 697.050 478.050 699.150 ;
        RECT 470.250 695.700 472.050 696.600 ;
        RECT 506.550 695.700 507.750 703.050 ;
        RECT 508.950 701.850 511.050 703.950 ;
        RECT 541.950 703.050 544.050 705.150 ;
        RECT 545.850 702.150 547.050 707.400 ;
        RECT 585.000 706.350 587.550 707.400 ;
        RECT 551.100 702.150 552.900 703.950 ;
        RECT 581.100 702.150 582.900 703.950 ;
        RECT 509.100 700.050 510.900 701.850 ;
        RECT 544.950 700.050 547.050 702.150 ;
        RECT 544.950 696.750 546.150 700.050 ;
        RECT 547.950 698.850 550.050 700.950 ;
        RECT 550.950 700.050 553.050 702.150 ;
        RECT 580.950 700.050 583.050 702.150 ;
        RECT 585.000 699.150 586.050 706.350 ;
        RECT 620.550 705.150 621.750 713.400 ;
        RECT 658.350 707.400 660.150 719.250 ;
        RECT 661.350 707.400 663.150 719.250 ;
        RECT 664.650 713.400 666.450 719.250 ;
        RECT 692.550 713.400 694.350 719.250 ;
        RECT 695.550 713.400 697.350 719.250 ;
        RECT 698.550 713.400 700.350 719.250 ;
        RECT 587.100 702.150 588.900 703.950 ;
        RECT 586.950 700.050 589.050 702.150 ;
        RECT 616.950 701.850 619.050 703.950 ;
        RECT 619.950 703.050 622.050 705.150 ;
        RECT 617.100 700.050 618.900 701.850 ;
        RECT 548.100 697.050 549.900 698.850 ;
        RECT 583.950 697.050 586.050 699.150 ;
        RECT 542.250 695.700 546.000 696.750 ;
        RECT 470.250 694.800 473.550 695.700 ;
        RECT 506.550 694.800 510.150 695.700 ;
        RECT 386.550 687.750 388.350 690.600 ;
        RECT 389.550 687.750 391.350 690.600 ;
        RECT 392.550 687.750 394.350 690.600 ;
        RECT 425.550 687.750 427.350 690.600 ;
        RECT 428.850 687.750 430.650 693.600 ;
        RECT 431.850 687.750 433.650 693.600 ;
        RECT 466.650 687.750 468.450 693.600 ;
        RECT 472.650 690.600 473.550 694.800 ;
        RECT 469.650 687.750 471.450 690.600 ;
        RECT 472.650 687.750 474.450 690.600 ;
        RECT 475.650 687.750 477.450 690.600 ;
        RECT 503.850 687.750 505.650 693.600 ;
        RECT 508.350 687.750 510.150 694.800 ;
        RECT 542.250 693.600 543.450 695.700 ;
        RECT 541.650 687.750 543.450 693.600 ;
        RECT 544.650 692.700 552.450 694.050 ;
        RECT 544.650 687.750 546.450 692.700 ;
        RECT 547.650 687.750 549.450 691.800 ;
        RECT 550.650 687.750 552.450 692.700 ;
        RECT 585.000 690.600 586.050 697.050 ;
        RECT 620.550 695.700 621.750 703.050 ;
        RECT 622.950 701.850 625.050 703.950 ;
        RECT 658.650 702.150 659.850 707.400 ;
        RECT 665.250 706.500 666.450 713.400 ;
        RECT 660.750 705.600 666.450 706.500 ;
        RECT 660.750 704.700 663.000 705.600 ;
        RECT 695.550 705.150 696.750 713.400 ;
        RECT 731.550 707.400 733.350 719.250 ;
        RECT 736.050 707.550 737.850 719.250 ;
        RECT 739.050 708.900 740.850 719.250 ;
        RECT 739.050 707.550 741.450 708.900 ;
        RECT 731.550 706.200 732.750 707.400 ;
        RECT 736.950 706.200 738.750 706.650 ;
        RECT 623.100 700.050 624.900 701.850 ;
        RECT 658.650 700.050 661.050 702.150 ;
        RECT 620.550 694.800 624.150 695.700 ;
        RECT 581.550 687.750 583.350 690.600 ;
        RECT 584.550 687.750 586.350 690.600 ;
        RECT 587.550 687.750 589.350 690.600 ;
        RECT 617.850 687.750 619.650 693.600 ;
        RECT 622.350 687.750 624.150 694.800 ;
        RECT 658.650 693.600 659.850 700.050 ;
        RECT 661.950 696.300 663.000 704.700 ;
        RECT 665.100 702.150 666.900 703.950 ;
        RECT 664.950 700.050 667.050 702.150 ;
        RECT 691.950 701.850 694.050 703.950 ;
        RECT 694.950 703.050 697.050 705.150 ;
        RECT 731.550 705.000 738.750 706.200 ;
        RECT 736.950 704.850 738.750 705.000 ;
        RECT 692.100 700.050 693.900 701.850 ;
        RECT 660.750 695.400 663.000 696.300 ;
        RECT 695.550 695.700 696.750 703.050 ;
        RECT 697.950 701.850 700.050 703.950 ;
        RECT 734.100 702.150 735.900 703.950 ;
        RECT 698.100 700.050 699.900 701.850 ;
        RECT 731.100 699.150 732.900 700.950 ;
        RECT 733.950 700.050 736.050 702.150 ;
        RECT 730.950 697.050 733.050 699.150 ;
        RECT 737.700 696.600 738.600 704.850 ;
        RECT 740.100 700.950 741.450 707.550 ;
        RECT 739.950 698.850 742.050 700.950 ;
        RECT 736.950 695.700 738.750 696.600 ;
        RECT 660.750 694.500 665.850 695.400 ;
        RECT 695.550 694.800 699.150 695.700 ;
        RECT 658.350 687.750 660.150 693.600 ;
        RECT 661.350 687.750 663.150 693.600 ;
        RECT 664.650 690.600 665.850 694.500 ;
        RECT 664.650 687.750 666.450 690.600 ;
        RECT 692.850 687.750 694.650 693.600 ;
        RECT 697.350 687.750 699.150 694.800 ;
        RECT 735.450 694.800 738.750 695.700 ;
        RECT 735.450 690.600 736.350 694.800 ;
        RECT 741.000 693.600 742.050 698.850 ;
        RECT 731.550 687.750 733.350 690.600 ;
        RECT 734.550 687.750 736.350 690.600 ;
        RECT 737.550 687.750 739.350 690.600 ;
        RECT 740.550 687.750 742.350 693.600 ;
        RECT 29.850 676.200 31.650 683.250 ;
        RECT 34.350 677.400 36.150 683.250 ;
        RECT 67.650 677.400 69.450 683.250 ;
        RECT 70.650 680.400 72.450 683.250 ;
        RECT 73.650 680.400 75.450 683.250 ;
        RECT 76.650 680.400 78.450 683.250 ;
        RECT 106.650 680.400 108.450 683.250 ;
        RECT 109.650 680.400 111.450 683.250 ;
        RECT 112.650 680.400 114.450 683.250 ;
        RECT 29.850 675.300 33.450 676.200 ;
        RECT 29.100 669.150 30.900 670.950 ;
        RECT 28.950 667.050 31.050 669.150 ;
        RECT 32.250 667.950 33.450 675.300 ;
        RECT 67.950 672.150 69.000 677.400 ;
        RECT 73.650 676.200 74.550 680.400 ;
        RECT 71.250 675.300 74.550 676.200 ;
        RECT 71.250 674.400 73.050 675.300 ;
        RECT 35.100 669.150 36.900 670.950 ;
        RECT 67.950 670.050 70.050 672.150 ;
        RECT 31.950 665.850 34.050 667.950 ;
        RECT 34.950 667.050 37.050 669.150 ;
        RECT 32.250 657.600 33.450 665.850 ;
        RECT 68.550 663.450 69.900 670.050 ;
        RECT 71.400 666.150 72.300 674.400 ;
        RECT 109.950 673.950 111.000 680.400 ;
        RECT 116.550 677.400 118.350 683.250 ;
        RECT 119.850 680.400 121.650 683.250 ;
        RECT 124.350 680.400 126.150 683.250 ;
        RECT 128.550 680.400 130.350 683.250 ;
        RECT 132.450 680.400 134.250 683.250 ;
        RECT 135.750 680.400 137.550 683.250 ;
        RECT 140.250 681.300 142.050 683.250 ;
        RECT 140.250 680.400 144.000 681.300 ;
        RECT 145.050 680.400 146.850 683.250 ;
        RECT 124.650 679.500 125.700 680.400 ;
        RECT 121.950 678.300 125.700 679.500 ;
        RECT 133.200 678.600 134.250 680.400 ;
        RECT 142.950 679.500 144.000 680.400 ;
        RECT 121.950 677.400 124.050 678.300 ;
        RECT 116.550 675.150 117.750 677.400 ;
        RECT 129.150 676.200 130.950 678.000 ;
        RECT 133.200 677.550 138.150 678.600 ;
        RECT 136.350 676.800 138.150 677.550 ;
        RECT 139.650 676.800 141.450 678.600 ;
        RECT 142.950 677.400 145.050 679.500 ;
        RECT 148.050 677.400 149.850 683.250 ;
        RECT 182.700 680.400 184.500 683.250 ;
        RECT 186.000 679.050 187.800 683.250 ;
        RECT 130.050 675.900 130.950 676.200 ;
        RECT 140.100 675.900 141.150 676.800 ;
        RECT 76.950 671.850 79.050 673.950 ;
        RECT 109.950 671.850 112.050 673.950 ;
        RECT 116.550 673.050 121.050 675.150 ;
        RECT 130.050 675.000 141.150 675.900 ;
        RECT 73.950 668.850 76.050 670.950 ;
        RECT 77.100 670.050 78.900 671.850 ;
        RECT 106.950 668.850 109.050 670.950 ;
        RECT 74.100 667.050 75.900 668.850 ;
        RECT 107.100 667.050 108.900 668.850 ;
        RECT 71.250 666.000 73.050 666.150 ;
        RECT 71.250 664.800 78.450 666.000 ;
        RECT 71.250 664.350 73.050 664.800 ;
        RECT 77.250 663.600 78.450 664.800 ;
        RECT 109.950 664.650 111.000 671.850 ;
        RECT 112.950 668.850 115.050 670.950 ;
        RECT 113.100 667.050 114.900 668.850 ;
        RECT 68.550 662.100 70.950 663.450 ;
        RECT 28.650 651.750 30.450 657.600 ;
        RECT 31.650 651.750 33.450 657.600 ;
        RECT 34.650 651.750 36.450 657.600 ;
        RECT 69.150 651.750 70.950 662.100 ;
        RECT 72.150 651.750 73.950 663.450 ;
        RECT 76.650 651.750 78.450 663.600 ;
        RECT 108.450 663.600 111.000 664.650 ;
        RECT 116.550 663.600 117.750 673.050 ;
        RECT 118.950 671.250 122.850 673.050 ;
        RECT 118.950 670.950 121.050 671.250 ;
        RECT 130.050 670.950 130.950 675.000 ;
        RECT 140.100 673.800 141.150 675.000 ;
        RECT 140.100 672.600 147.000 673.800 ;
        RECT 140.100 672.000 141.900 672.600 ;
        RECT 146.100 671.850 147.000 672.600 ;
        RECT 143.100 670.950 144.900 671.700 ;
        RECT 130.050 668.850 133.050 670.950 ;
        RECT 136.950 669.900 144.900 670.950 ;
        RECT 146.100 670.050 147.900 671.850 ;
        RECT 136.950 668.850 139.050 669.900 ;
        RECT 118.950 665.400 120.750 667.200 ;
        RECT 119.850 664.200 124.050 665.400 ;
        RECT 130.050 664.200 130.950 668.850 ;
        RECT 138.750 665.100 140.550 665.400 ;
        RECT 108.450 651.750 110.250 663.600 ;
        RECT 112.650 651.750 114.450 663.600 ;
        RECT 116.550 651.750 118.350 663.600 ;
        RECT 121.950 663.300 124.050 664.200 ;
        RECT 124.950 663.300 130.950 664.200 ;
        RECT 132.150 664.800 140.550 665.100 ;
        RECT 148.950 664.800 149.850 677.400 ;
        RECT 182.100 677.400 187.800 679.050 ;
        RECT 190.200 677.400 192.000 683.250 ;
        RECT 221.550 678.300 223.350 683.250 ;
        RECT 224.550 679.200 226.350 683.250 ;
        RECT 227.550 678.300 229.350 683.250 ;
        RECT 182.100 670.950 183.300 677.400 ;
        RECT 221.550 676.950 229.350 678.300 ;
        RECT 230.550 677.400 232.350 683.250 ;
        RECT 236.550 677.400 238.350 683.250 ;
        RECT 239.850 680.400 241.650 683.250 ;
        RECT 244.350 680.400 246.150 683.250 ;
        RECT 248.550 680.400 250.350 683.250 ;
        RECT 252.450 680.400 254.250 683.250 ;
        RECT 255.750 680.400 257.550 683.250 ;
        RECT 260.250 681.300 262.050 683.250 ;
        RECT 260.250 680.400 264.000 681.300 ;
        RECT 265.050 680.400 266.850 683.250 ;
        RECT 244.650 679.500 245.700 680.400 ;
        RECT 241.950 678.300 245.700 679.500 ;
        RECT 253.200 678.600 254.250 680.400 ;
        RECT 262.950 679.500 264.000 680.400 ;
        RECT 241.950 677.400 244.050 678.300 ;
        RECT 230.550 675.300 231.750 677.400 ;
        RECT 228.000 674.250 231.750 675.300 ;
        RECT 236.550 675.150 237.750 677.400 ;
        RECT 249.150 676.200 250.950 678.000 ;
        RECT 253.200 677.550 258.150 678.600 ;
        RECT 256.350 676.800 258.150 677.550 ;
        RECT 259.650 676.800 261.450 678.600 ;
        RECT 262.950 677.400 265.050 679.500 ;
        RECT 268.050 677.400 269.850 683.250 ;
        RECT 250.050 675.900 250.950 676.200 ;
        RECT 260.100 675.900 261.150 676.800 ;
        RECT 185.100 672.150 186.900 673.950 ;
        RECT 181.950 668.850 184.050 670.950 ;
        RECT 184.950 670.050 187.050 672.150 ;
        RECT 187.950 671.850 190.050 673.950 ;
        RECT 191.100 672.150 192.900 673.950 ;
        RECT 224.100 672.150 225.900 673.950 ;
        RECT 188.100 670.050 189.900 671.850 ;
        RECT 190.950 670.050 193.050 672.150 ;
        RECT 220.950 668.850 223.050 670.950 ;
        RECT 223.950 670.050 226.050 672.150 ;
        RECT 227.850 670.950 229.050 674.250 ;
        RECT 226.950 668.850 229.050 670.950 ;
        RECT 236.550 673.050 241.050 675.150 ;
        RECT 250.050 675.000 261.150 675.900 ;
        RECT 132.150 664.200 149.850 664.800 ;
        RECT 124.950 662.400 125.850 663.300 ;
        RECT 123.150 660.600 125.850 662.400 ;
        RECT 126.750 662.100 128.550 662.400 ;
        RECT 132.150 662.100 133.050 664.200 ;
        RECT 138.750 663.600 149.850 664.200 ;
        RECT 182.100 663.600 183.300 668.850 ;
        RECT 221.100 667.050 222.900 668.850 ;
        RECT 190.950 666.450 193.050 667.050 ;
        RECT 217.950 666.450 220.050 667.050 ;
        RECT 190.950 665.550 220.050 666.450 ;
        RECT 190.950 664.950 193.050 665.550 ;
        RECT 217.950 664.950 220.050 665.550 ;
        RECT 226.950 663.600 228.150 668.850 ;
        RECT 229.950 665.850 232.050 667.950 ;
        RECT 229.950 664.050 231.750 665.850 ;
        RECT 236.550 663.600 237.750 673.050 ;
        RECT 238.950 671.250 242.850 673.050 ;
        RECT 238.950 670.950 241.050 671.250 ;
        RECT 250.050 670.950 250.950 675.000 ;
        RECT 260.100 673.800 261.150 675.000 ;
        RECT 260.100 672.600 267.000 673.800 ;
        RECT 260.100 672.000 261.900 672.600 ;
        RECT 266.100 671.850 267.000 672.600 ;
        RECT 263.100 670.950 264.900 671.700 ;
        RECT 250.050 668.850 253.050 670.950 ;
        RECT 256.950 669.900 264.900 670.950 ;
        RECT 266.100 670.050 267.900 671.850 ;
        RECT 256.950 668.850 259.050 669.900 ;
        RECT 238.950 665.400 240.750 667.200 ;
        RECT 239.850 664.200 244.050 665.400 ;
        RECT 250.050 664.200 250.950 668.850 ;
        RECT 258.750 665.100 260.550 665.400 ;
        RECT 126.750 661.200 133.050 662.100 ;
        RECT 133.950 662.700 135.750 663.300 ;
        RECT 133.950 661.500 141.450 662.700 ;
        RECT 126.750 660.600 128.550 661.200 ;
        RECT 140.250 660.600 141.450 661.500 ;
        RECT 121.950 657.600 125.850 659.700 ;
        RECT 130.950 658.500 137.850 660.300 ;
        RECT 140.250 658.500 145.050 660.600 ;
        RECT 119.550 651.750 121.350 654.600 ;
        RECT 124.050 651.750 125.850 657.600 ;
        RECT 128.250 651.750 130.050 657.600 ;
        RECT 132.150 651.750 133.950 658.500 ;
        RECT 140.250 657.600 141.450 658.500 ;
        RECT 135.150 651.750 136.950 657.600 ;
        RECT 139.950 651.750 141.750 657.600 ;
        RECT 145.050 651.750 146.850 657.600 ;
        RECT 148.050 651.750 149.850 663.600 ;
        RECT 181.650 651.750 183.450 663.600 ;
        RECT 184.650 662.700 192.450 663.600 ;
        RECT 184.650 651.750 186.450 662.700 ;
        RECT 187.650 651.750 189.450 661.800 ;
        RECT 190.650 651.750 192.450 662.700 ;
        RECT 222.300 651.750 224.100 663.600 ;
        RECT 226.500 651.750 228.300 663.600 ;
        RECT 229.800 651.750 231.600 657.600 ;
        RECT 236.550 651.750 238.350 663.600 ;
        RECT 241.950 663.300 244.050 664.200 ;
        RECT 244.950 663.300 250.950 664.200 ;
        RECT 252.150 664.800 260.550 665.100 ;
        RECT 268.950 664.800 269.850 677.400 ;
        RECT 252.150 664.200 269.850 664.800 ;
        RECT 244.950 662.400 245.850 663.300 ;
        RECT 243.150 660.600 245.850 662.400 ;
        RECT 246.750 662.100 248.550 662.400 ;
        RECT 252.150 662.100 253.050 664.200 ;
        RECT 258.750 663.600 269.850 664.200 ;
        RECT 246.750 661.200 253.050 662.100 ;
        RECT 253.950 662.700 255.750 663.300 ;
        RECT 253.950 661.500 261.450 662.700 ;
        RECT 246.750 660.600 248.550 661.200 ;
        RECT 260.250 660.600 261.450 661.500 ;
        RECT 241.950 657.600 245.850 659.700 ;
        RECT 250.950 658.500 257.850 660.300 ;
        RECT 260.250 658.500 265.050 660.600 ;
        RECT 239.550 651.750 241.350 654.600 ;
        RECT 244.050 651.750 245.850 657.600 ;
        RECT 248.250 651.750 250.050 657.600 ;
        RECT 252.150 651.750 253.950 658.500 ;
        RECT 260.250 657.600 261.450 658.500 ;
        RECT 255.150 651.750 256.950 657.600 ;
        RECT 259.950 651.750 261.750 657.600 ;
        RECT 265.050 651.750 266.850 657.600 ;
        RECT 268.050 651.750 269.850 663.600 ;
        RECT 272.550 677.400 274.350 683.250 ;
        RECT 275.850 680.400 277.650 683.250 ;
        RECT 280.350 680.400 282.150 683.250 ;
        RECT 284.550 680.400 286.350 683.250 ;
        RECT 288.450 680.400 290.250 683.250 ;
        RECT 291.750 680.400 293.550 683.250 ;
        RECT 296.250 681.300 298.050 683.250 ;
        RECT 296.250 680.400 300.000 681.300 ;
        RECT 301.050 680.400 302.850 683.250 ;
        RECT 280.650 679.500 281.700 680.400 ;
        RECT 277.950 678.300 281.700 679.500 ;
        RECT 289.200 678.600 290.250 680.400 ;
        RECT 298.950 679.500 300.000 680.400 ;
        RECT 277.950 677.400 280.050 678.300 ;
        RECT 272.550 675.150 273.750 677.400 ;
        RECT 285.150 676.200 286.950 678.000 ;
        RECT 289.200 677.550 294.150 678.600 ;
        RECT 292.350 676.800 294.150 677.550 ;
        RECT 295.650 676.800 297.450 678.600 ;
        RECT 298.950 677.400 301.050 679.500 ;
        RECT 304.050 677.400 305.850 683.250 ;
        RECT 338.700 680.400 340.500 683.250 ;
        RECT 342.000 679.050 343.800 683.250 ;
        RECT 286.050 675.900 286.950 676.200 ;
        RECT 296.100 675.900 297.150 676.800 ;
        RECT 272.550 673.050 277.050 675.150 ;
        RECT 286.050 675.000 297.150 675.900 ;
        RECT 272.550 663.600 273.750 673.050 ;
        RECT 274.950 671.250 278.850 673.050 ;
        RECT 274.950 670.950 277.050 671.250 ;
        RECT 286.050 670.950 286.950 675.000 ;
        RECT 296.100 673.800 297.150 675.000 ;
        RECT 296.100 672.600 303.000 673.800 ;
        RECT 296.100 672.000 297.900 672.600 ;
        RECT 302.100 671.850 303.000 672.600 ;
        RECT 299.100 670.950 300.900 671.700 ;
        RECT 286.050 668.850 289.050 670.950 ;
        RECT 292.950 669.900 300.900 670.950 ;
        RECT 302.100 670.050 303.900 671.850 ;
        RECT 292.950 668.850 295.050 669.900 ;
        RECT 274.950 665.400 276.750 667.200 ;
        RECT 275.850 664.200 280.050 665.400 ;
        RECT 286.050 664.200 286.950 668.850 ;
        RECT 294.750 665.100 296.550 665.400 ;
        RECT 272.550 651.750 274.350 663.600 ;
        RECT 277.950 663.300 280.050 664.200 ;
        RECT 280.950 663.300 286.950 664.200 ;
        RECT 288.150 664.800 296.550 665.100 ;
        RECT 304.950 664.800 305.850 677.400 ;
        RECT 338.100 677.400 343.800 679.050 ;
        RECT 346.200 677.400 348.000 683.250 ;
        RECT 338.100 670.950 339.300 677.400 ;
        RECT 380.850 676.200 382.650 683.250 ;
        RECT 385.350 677.400 387.150 683.250 ;
        RECT 418.650 677.400 420.450 683.250 ;
        RECT 380.850 675.300 384.450 676.200 ;
        RECT 341.100 672.150 342.900 673.950 ;
        RECT 337.950 668.850 340.050 670.950 ;
        RECT 340.950 670.050 343.050 672.150 ;
        RECT 343.950 671.850 346.050 673.950 ;
        RECT 347.100 672.150 348.900 673.950 ;
        RECT 344.100 670.050 345.900 671.850 ;
        RECT 346.950 670.050 349.050 672.150 ;
        RECT 380.100 669.150 381.900 670.950 ;
        RECT 288.150 664.200 305.850 664.800 ;
        RECT 280.950 662.400 281.850 663.300 ;
        RECT 279.150 660.600 281.850 662.400 ;
        RECT 282.750 662.100 284.550 662.400 ;
        RECT 288.150 662.100 289.050 664.200 ;
        RECT 294.750 663.600 305.850 664.200 ;
        RECT 338.100 663.600 339.300 668.850 ;
        RECT 379.950 667.050 382.050 669.150 ;
        RECT 383.250 667.950 384.450 675.300 ;
        RECT 419.250 675.300 420.450 677.400 ;
        RECT 421.650 678.300 423.450 683.250 ;
        RECT 424.650 679.200 426.450 683.250 ;
        RECT 427.650 678.300 429.450 683.250 ;
        RECT 421.650 676.950 429.450 678.300 ;
        RECT 460.650 677.400 462.450 683.250 ;
        RECT 463.650 680.400 465.450 683.250 ;
        RECT 466.650 680.400 468.450 683.250 ;
        RECT 469.650 680.400 471.450 683.250 ;
        RECT 500.550 680.400 502.350 683.250 ;
        RECT 503.550 680.400 505.350 683.250 ;
        RECT 506.550 680.400 508.350 683.250 ;
        RECT 419.250 674.250 423.000 675.300 ;
        RECT 418.950 672.450 421.050 673.050 ;
        RECT 416.550 671.550 421.050 672.450 ;
        RECT 386.100 669.150 387.900 670.950 ;
        RECT 382.950 665.850 385.050 667.950 ;
        RECT 385.950 667.050 388.050 669.150 ;
        RECT 282.750 661.200 289.050 662.100 ;
        RECT 289.950 662.700 291.750 663.300 ;
        RECT 289.950 661.500 297.450 662.700 ;
        RECT 282.750 660.600 284.550 661.200 ;
        RECT 296.250 660.600 297.450 661.500 ;
        RECT 277.950 657.600 281.850 659.700 ;
        RECT 286.950 658.500 293.850 660.300 ;
        RECT 296.250 658.500 301.050 660.600 ;
        RECT 275.550 651.750 277.350 654.600 ;
        RECT 280.050 651.750 281.850 657.600 ;
        RECT 284.250 651.750 286.050 657.600 ;
        RECT 288.150 651.750 289.950 658.500 ;
        RECT 296.250 657.600 297.450 658.500 ;
        RECT 291.150 651.750 292.950 657.600 ;
        RECT 295.950 651.750 297.750 657.600 ;
        RECT 301.050 651.750 302.850 657.600 ;
        RECT 304.050 651.750 305.850 663.600 ;
        RECT 337.650 651.750 339.450 663.600 ;
        RECT 340.650 662.700 348.450 663.600 ;
        RECT 340.650 651.750 342.450 662.700 ;
        RECT 343.650 651.750 345.450 661.800 ;
        RECT 346.650 651.750 348.450 662.700 ;
        RECT 383.250 657.600 384.450 665.850 ;
        RECT 416.550 660.450 417.450 671.550 ;
        RECT 418.950 670.950 421.050 671.550 ;
        RECT 421.950 670.950 423.150 674.250 ;
        RECT 425.100 672.150 426.900 673.950 ;
        RECT 460.950 672.150 462.000 677.400 ;
        RECT 466.650 676.200 467.550 680.400 ;
        RECT 464.250 675.300 467.550 676.200 ;
        RECT 464.250 674.400 466.050 675.300 ;
        RECT 421.950 668.850 424.050 670.950 ;
        RECT 424.950 670.050 427.050 672.150 ;
        RECT 427.950 668.850 430.050 670.950 ;
        RECT 460.950 670.050 463.050 672.150 ;
        RECT 418.950 665.850 421.050 667.950 ;
        RECT 419.250 664.050 421.050 665.850 ;
        RECT 422.850 663.600 424.050 668.850 ;
        RECT 428.100 667.050 429.900 668.850 ;
        RECT 418.950 660.450 421.050 661.050 ;
        RECT 416.550 659.550 421.050 660.450 ;
        RECT 418.950 658.950 421.050 659.550 ;
        RECT 379.650 651.750 381.450 657.600 ;
        RECT 382.650 651.750 384.450 657.600 ;
        RECT 385.650 651.750 387.450 657.600 ;
        RECT 419.400 651.750 421.200 657.600 ;
        RECT 422.700 651.750 424.500 663.600 ;
        RECT 426.900 651.750 428.700 663.600 ;
        RECT 461.550 663.450 462.900 670.050 ;
        RECT 464.400 666.150 465.300 674.400 ;
        RECT 504.000 673.950 505.050 680.400 ;
        RECT 539.850 677.400 541.650 683.250 ;
        RECT 544.350 676.200 546.150 683.250 ;
        RECT 578.550 678.300 580.350 683.250 ;
        RECT 581.550 679.200 583.350 683.250 ;
        RECT 584.550 678.300 586.350 683.250 ;
        RECT 578.550 676.950 586.350 678.300 ;
        RECT 587.550 677.400 589.350 683.250 ;
        RECT 620.850 677.400 622.650 683.250 ;
        RECT 469.950 671.850 472.050 673.950 ;
        RECT 502.950 671.850 505.050 673.950 ;
        RECT 466.950 668.850 469.050 670.950 ;
        RECT 470.100 670.050 471.900 671.850 ;
        RECT 499.950 668.850 502.050 670.950 ;
        RECT 467.100 667.050 468.900 668.850 ;
        RECT 500.100 667.050 501.900 668.850 ;
        RECT 464.250 666.000 466.050 666.150 ;
        RECT 464.250 664.800 471.450 666.000 ;
        RECT 464.250 664.350 466.050 664.800 ;
        RECT 470.250 663.600 471.450 664.800 ;
        RECT 504.000 664.650 505.050 671.850 ;
        RECT 542.550 675.300 546.150 676.200 ;
        RECT 587.550 675.300 588.750 677.400 ;
        RECT 625.350 676.200 627.150 683.250 ;
        RECT 505.950 668.850 508.050 670.950 ;
        RECT 539.100 669.150 540.900 670.950 ;
        RECT 506.100 667.050 507.900 668.850 ;
        RECT 538.950 667.050 541.050 669.150 ;
        RECT 542.550 667.950 543.750 675.300 ;
        RECT 585.000 674.250 588.750 675.300 ;
        RECT 623.550 675.300 627.150 676.200 ;
        RECT 662.850 676.200 664.650 683.250 ;
        RECT 667.350 677.400 669.150 683.250 ;
        RECT 698.550 680.400 700.350 683.250 ;
        RECT 701.550 680.400 703.350 683.250 ;
        RECT 704.550 680.400 706.350 683.250 ;
        RECT 702.450 676.200 703.350 680.400 ;
        RECT 707.550 677.400 709.350 683.250 ;
        RECT 740.850 677.400 742.650 683.250 ;
        RECT 662.850 675.300 666.450 676.200 ;
        RECT 702.450 675.300 705.750 676.200 ;
        RECT 581.100 672.150 582.900 673.950 ;
        RECT 545.100 669.150 546.900 670.950 ;
        RECT 541.950 665.850 544.050 667.950 ;
        RECT 544.950 667.050 547.050 669.150 ;
        RECT 577.950 668.850 580.050 670.950 ;
        RECT 580.950 670.050 583.050 672.150 ;
        RECT 584.850 670.950 586.050 674.250 ;
        RECT 583.950 668.850 586.050 670.950 ;
        RECT 620.100 669.150 621.900 670.950 ;
        RECT 578.100 667.050 579.900 668.850 ;
        RECT 504.000 663.600 506.550 664.650 ;
        RECT 461.550 662.100 463.950 663.450 ;
        RECT 462.150 651.750 463.950 662.100 ;
        RECT 465.150 651.750 466.950 663.450 ;
        RECT 469.650 651.750 471.450 663.600 ;
        RECT 500.550 651.750 502.350 663.600 ;
        RECT 504.750 651.750 506.550 663.600 ;
        RECT 542.550 657.600 543.750 665.850 ;
        RECT 583.950 663.600 585.150 668.850 ;
        RECT 586.950 665.850 589.050 667.950 ;
        RECT 619.950 667.050 622.050 669.150 ;
        RECT 623.550 667.950 624.750 675.300 ;
        RECT 626.100 669.150 627.900 670.950 ;
        RECT 662.100 669.150 663.900 670.950 ;
        RECT 622.950 665.850 625.050 667.950 ;
        RECT 625.950 667.050 628.050 669.150 ;
        RECT 661.950 667.050 664.050 669.150 ;
        RECT 665.250 667.950 666.450 675.300 ;
        RECT 703.950 674.400 705.750 675.300 ;
        RECT 697.950 671.850 700.050 673.950 ;
        RECT 668.100 669.150 669.900 670.950 ;
        RECT 698.100 670.050 699.900 671.850 ;
        RECT 664.950 665.850 667.050 667.950 ;
        RECT 667.950 667.050 670.050 669.150 ;
        RECT 700.950 668.850 703.050 670.950 ;
        RECT 701.100 667.050 702.900 668.850 ;
        RECT 704.700 666.150 705.600 674.400 ;
        RECT 708.000 672.150 709.050 677.400 ;
        RECT 745.350 676.200 747.150 683.250 ;
        RECT 706.950 670.050 709.050 672.150 ;
        RECT 743.550 675.300 747.150 676.200 ;
        RECT 703.950 666.000 705.750 666.150 ;
        RECT 586.950 664.050 588.750 665.850 ;
        RECT 539.550 651.750 541.350 657.600 ;
        RECT 542.550 651.750 544.350 657.600 ;
        RECT 545.550 651.750 547.350 657.600 ;
        RECT 579.300 651.750 581.100 663.600 ;
        RECT 583.500 651.750 585.300 663.600 ;
        RECT 623.550 657.600 624.750 665.850 ;
        RECT 665.250 657.600 666.450 665.850 ;
        RECT 698.550 664.800 705.750 666.000 ;
        RECT 698.550 663.600 699.750 664.800 ;
        RECT 703.950 664.350 705.750 664.800 ;
        RECT 586.800 651.750 588.600 657.600 ;
        RECT 620.550 651.750 622.350 657.600 ;
        RECT 623.550 651.750 625.350 657.600 ;
        RECT 626.550 651.750 628.350 657.600 ;
        RECT 661.650 651.750 663.450 657.600 ;
        RECT 664.650 651.750 666.450 657.600 ;
        RECT 667.650 651.750 669.450 657.600 ;
        RECT 698.550 651.750 700.350 663.600 ;
        RECT 707.100 663.450 708.450 670.050 ;
        RECT 740.100 669.150 741.900 670.950 ;
        RECT 739.950 667.050 742.050 669.150 ;
        RECT 743.550 667.950 744.750 675.300 ;
        RECT 746.100 669.150 747.900 670.950 ;
        RECT 742.950 665.850 745.050 667.950 ;
        RECT 745.950 667.050 748.050 669.150 ;
        RECT 703.050 651.750 704.850 663.450 ;
        RECT 706.050 662.100 708.450 663.450 ;
        RECT 706.050 651.750 707.850 662.100 ;
        RECT 743.550 657.600 744.750 665.850 ;
        RECT 740.550 651.750 742.350 657.600 ;
        RECT 743.550 651.750 745.350 657.600 ;
        RECT 746.550 651.750 748.350 657.600 ;
        RECT 31.650 641.400 33.450 647.250 ;
        RECT 34.650 641.400 36.450 647.250 ;
        RECT 68.400 641.400 70.200 647.250 ;
        RECT 32.400 628.950 33.600 641.400 ;
        RECT 71.700 635.400 73.500 647.250 ;
        RECT 75.900 635.400 77.700 647.250 ;
        RECT 109.650 641.400 111.450 647.250 ;
        RECT 112.650 641.400 114.450 647.250 ;
        RECT 115.650 641.400 117.450 647.250 ;
        RECT 143.550 641.400 145.350 647.250 ;
        RECT 146.550 641.400 148.350 647.250 ;
        RECT 179.550 641.400 181.350 647.250 ;
        RECT 182.550 641.400 184.350 647.250 ;
        RECT 185.550 641.400 187.350 647.250 ;
        RECT 221.400 641.400 223.200 647.250 ;
        RECT 68.250 633.150 70.050 634.950 ;
        RECT 67.950 631.050 70.050 633.150 ;
        RECT 71.850 630.150 73.050 635.400 ;
        RECT 113.250 633.150 114.450 641.400 ;
        RECT 77.100 630.150 78.900 631.950 ;
        RECT 31.950 626.850 34.050 628.950 ;
        RECT 35.100 627.150 36.900 628.950 ;
        RECT 70.950 628.050 73.050 630.150 ;
        RECT 32.400 618.600 33.600 626.850 ;
        RECT 34.950 625.050 37.050 627.150 ;
        RECT 70.950 624.750 72.150 628.050 ;
        RECT 73.950 626.850 76.050 628.950 ;
        RECT 76.950 628.050 79.050 630.150 ;
        RECT 109.950 629.850 112.050 631.950 ;
        RECT 112.950 631.050 115.050 633.150 ;
        RECT 110.100 628.050 111.900 629.850 ;
        RECT 74.100 625.050 75.900 626.850 ;
        RECT 68.250 623.700 72.000 624.750 ;
        RECT 113.250 623.700 114.450 631.050 ;
        RECT 115.950 629.850 118.050 631.950 ;
        RECT 116.100 628.050 117.900 629.850 ;
        RECT 146.400 628.950 147.600 641.400 ;
        RECT 182.550 633.150 183.750 641.400 ;
        RECT 224.700 635.400 226.500 647.250 ;
        RECT 228.900 635.400 230.700 647.250 ;
        RECT 259.650 641.400 261.450 647.250 ;
        RECT 262.650 641.400 264.450 647.250 ;
        RECT 265.650 641.400 267.450 647.250 ;
        RECT 221.250 633.150 223.050 634.950 ;
        RECT 178.950 629.850 181.050 631.950 ;
        RECT 181.950 631.050 184.050 633.150 ;
        RECT 143.100 627.150 144.900 628.950 ;
        RECT 142.950 625.050 145.050 627.150 ;
        RECT 145.950 626.850 148.050 628.950 ;
        RECT 179.100 628.050 180.900 629.850 ;
        RECT 68.250 621.600 69.450 623.700 ;
        RECT 110.850 622.800 114.450 623.700 ;
        RECT 31.650 615.750 33.450 618.600 ;
        RECT 34.650 615.750 36.450 618.600 ;
        RECT 67.650 615.750 69.450 621.600 ;
        RECT 70.650 620.700 78.450 622.050 ;
        RECT 70.650 615.750 72.450 620.700 ;
        RECT 73.650 615.750 75.450 619.800 ;
        RECT 76.650 615.750 78.450 620.700 ;
        RECT 110.850 615.750 112.650 622.800 ;
        RECT 115.350 615.750 117.150 621.600 ;
        RECT 146.400 618.600 147.600 626.850 ;
        RECT 182.550 623.700 183.750 631.050 ;
        RECT 184.950 629.850 187.050 631.950 ;
        RECT 220.950 631.050 223.050 633.150 ;
        RECT 224.850 630.150 226.050 635.400 ;
        RECT 263.250 633.150 264.450 641.400 ;
        RECT 297.150 636.900 298.950 647.250 ;
        RECT 296.550 635.550 298.950 636.900 ;
        RECT 300.150 635.550 301.950 647.250 ;
        RECT 230.100 630.150 231.900 631.950 ;
        RECT 185.100 628.050 186.900 629.850 ;
        RECT 223.950 628.050 226.050 630.150 ;
        RECT 223.950 624.750 225.150 628.050 ;
        RECT 226.950 626.850 229.050 628.950 ;
        RECT 229.950 628.050 232.050 630.150 ;
        RECT 259.950 629.850 262.050 631.950 ;
        RECT 262.950 631.050 265.050 633.150 ;
        RECT 260.100 628.050 261.900 629.850 ;
        RECT 227.100 625.050 228.900 626.850 ;
        RECT 221.250 623.700 225.000 624.750 ;
        RECT 263.250 623.700 264.450 631.050 ;
        RECT 265.950 629.850 268.050 631.950 ;
        RECT 266.100 628.050 267.900 629.850 ;
        RECT 296.550 628.950 297.900 635.550 ;
        RECT 304.650 635.400 306.450 647.250 ;
        RECT 338.400 641.400 340.200 647.250 ;
        RECT 341.700 635.400 343.500 647.250 ;
        RECT 345.900 635.400 347.700 647.250 ;
        RECT 381.450 635.400 383.250 647.250 ;
        RECT 385.650 635.400 387.450 647.250 ;
        RECT 418.650 635.400 420.450 647.250 ;
        RECT 421.650 636.300 423.450 647.250 ;
        RECT 424.650 637.200 426.450 647.250 ;
        RECT 427.650 636.300 429.450 647.250 ;
        RECT 421.650 635.400 429.450 636.300 ;
        RECT 462.450 635.400 464.250 647.250 ;
        RECT 466.650 635.400 468.450 647.250 ;
        RECT 501.150 636.900 502.950 647.250 ;
        RECT 500.550 635.550 502.950 636.900 ;
        RECT 504.150 635.550 505.950 647.250 ;
        RECT 299.250 634.200 301.050 634.650 ;
        RECT 305.250 634.200 306.450 635.400 ;
        RECT 299.250 633.000 306.450 634.200 ;
        RECT 338.250 633.150 340.050 634.950 ;
        RECT 299.250 632.850 301.050 633.000 ;
        RECT 182.550 622.800 186.150 623.700 ;
        RECT 143.550 615.750 145.350 618.600 ;
        RECT 146.550 615.750 148.350 618.600 ;
        RECT 179.850 615.750 181.650 621.600 ;
        RECT 184.350 615.750 186.150 622.800 ;
        RECT 221.250 621.600 222.450 623.700 ;
        RECT 260.850 622.800 264.450 623.700 ;
        RECT 295.950 626.850 298.050 628.950 ;
        RECT 220.650 615.750 222.450 621.600 ;
        RECT 223.650 620.700 231.450 622.050 ;
        RECT 223.650 615.750 225.450 620.700 ;
        RECT 226.650 615.750 228.450 619.800 ;
        RECT 229.650 615.750 231.450 620.700 ;
        RECT 260.850 615.750 262.650 622.800 ;
        RECT 295.950 621.600 297.000 626.850 ;
        RECT 299.400 624.600 300.300 632.850 ;
        RECT 302.100 630.150 303.900 631.950 ;
        RECT 337.950 631.050 340.050 633.150 ;
        RECT 341.850 630.150 343.050 635.400 ;
        RECT 381.450 634.350 384.000 635.400 ;
        RECT 347.100 630.150 348.900 631.950 ;
        RECT 380.100 630.150 381.900 631.950 ;
        RECT 301.950 628.050 304.050 630.150 ;
        RECT 305.100 627.150 306.900 628.950 ;
        RECT 340.950 628.050 343.050 630.150 ;
        RECT 304.950 625.050 307.050 627.150 ;
        RECT 340.950 624.750 342.150 628.050 ;
        RECT 343.950 626.850 346.050 628.950 ;
        RECT 346.950 628.050 349.050 630.150 ;
        RECT 379.950 628.050 382.050 630.150 ;
        RECT 382.950 627.150 384.000 634.350 ;
        RECT 386.100 630.150 387.900 631.950 ;
        RECT 419.100 630.150 420.300 635.400 ;
        RECT 462.450 634.350 465.000 635.400 ;
        RECT 461.100 630.150 462.900 631.950 ;
        RECT 385.950 628.050 388.050 630.150 ;
        RECT 418.950 628.050 421.050 630.150 ;
        RECT 344.100 625.050 345.900 626.850 ;
        RECT 382.950 625.050 385.050 627.150 ;
        RECT 299.250 623.700 301.050 624.600 ;
        RECT 338.250 623.700 342.000 624.750 ;
        RECT 299.250 622.800 302.550 623.700 ;
        RECT 265.350 615.750 267.150 621.600 ;
        RECT 295.650 615.750 297.450 621.600 ;
        RECT 301.650 618.600 302.550 622.800 ;
        RECT 338.250 621.600 339.450 623.700 ;
        RECT 298.650 615.750 300.450 618.600 ;
        RECT 301.650 615.750 303.450 618.600 ;
        RECT 304.650 615.750 306.450 618.600 ;
        RECT 337.650 615.750 339.450 621.600 ;
        RECT 340.650 620.700 348.450 622.050 ;
        RECT 340.650 615.750 342.450 620.700 ;
        RECT 343.650 615.750 345.450 619.800 ;
        RECT 346.650 615.750 348.450 620.700 ;
        RECT 382.950 618.600 384.000 625.050 ;
        RECT 419.100 621.600 420.300 628.050 ;
        RECT 421.950 626.850 424.050 628.950 ;
        RECT 425.100 627.150 426.900 628.950 ;
        RECT 422.100 625.050 423.900 626.850 ;
        RECT 424.950 625.050 427.050 627.150 ;
        RECT 427.950 626.850 430.050 628.950 ;
        RECT 460.950 628.050 463.050 630.150 ;
        RECT 463.950 627.150 465.000 634.350 ;
        RECT 467.100 630.150 468.900 631.950 ;
        RECT 466.950 628.050 469.050 630.150 ;
        RECT 500.550 628.950 501.900 635.550 ;
        RECT 508.650 635.400 510.450 647.250 ;
        RECT 541.650 635.400 543.450 647.250 ;
        RECT 544.650 636.300 546.450 647.250 ;
        RECT 547.650 637.200 549.450 647.250 ;
        RECT 550.650 636.300 552.450 647.250 ;
        RECT 583.650 641.400 585.450 647.250 ;
        RECT 586.650 641.400 588.450 647.250 ;
        RECT 614.550 641.400 616.350 647.250 ;
        RECT 617.550 641.400 619.350 647.250 ;
        RECT 544.650 635.400 552.450 636.300 ;
        RECT 503.250 634.200 505.050 634.650 ;
        RECT 509.250 634.200 510.450 635.400 ;
        RECT 503.250 633.000 510.450 634.200 ;
        RECT 503.250 632.850 505.050 633.000 ;
        RECT 428.100 625.050 429.900 626.850 ;
        RECT 463.950 625.050 466.050 627.150 ;
        RECT 499.950 626.850 502.050 628.950 ;
        RECT 419.100 619.950 424.800 621.600 ;
        RECT 379.650 615.750 381.450 618.600 ;
        RECT 382.650 615.750 384.450 618.600 ;
        RECT 385.650 615.750 387.450 618.600 ;
        RECT 419.700 615.750 421.500 618.600 ;
        RECT 423.000 615.750 424.800 619.950 ;
        RECT 427.200 615.750 429.000 621.600 ;
        RECT 463.950 618.600 465.000 625.050 ;
        RECT 499.950 621.600 501.000 626.850 ;
        RECT 503.400 624.600 504.300 632.850 ;
        RECT 506.100 630.150 507.900 631.950 ;
        RECT 542.100 630.150 543.300 635.400 ;
        RECT 505.950 628.050 508.050 630.150 ;
        RECT 509.100 627.150 510.900 628.950 ;
        RECT 541.950 628.050 544.050 630.150 ;
        RECT 584.400 628.950 585.600 641.400 ;
        RECT 614.100 630.150 615.900 631.950 ;
        RECT 508.950 625.050 511.050 627.150 ;
        RECT 503.250 623.700 505.050 624.600 ;
        RECT 503.250 622.800 506.550 623.700 ;
        RECT 460.650 615.750 462.450 618.600 ;
        RECT 463.650 615.750 465.450 618.600 ;
        RECT 466.650 615.750 468.450 618.600 ;
        RECT 499.650 615.750 501.450 621.600 ;
        RECT 505.650 618.600 506.550 622.800 ;
        RECT 542.100 621.600 543.300 628.050 ;
        RECT 544.950 626.850 547.050 628.950 ;
        RECT 548.100 627.150 549.900 628.950 ;
        RECT 545.100 625.050 546.900 626.850 ;
        RECT 547.950 625.050 550.050 627.150 ;
        RECT 550.950 626.850 553.050 628.950 ;
        RECT 583.950 626.850 586.050 628.950 ;
        RECT 587.100 627.150 588.900 628.950 ;
        RECT 613.950 628.050 616.050 630.150 ;
        RECT 551.100 625.050 552.900 626.850 ;
        RECT 542.100 619.950 547.800 621.600 ;
        RECT 502.650 615.750 504.450 618.600 ;
        RECT 505.650 615.750 507.450 618.600 ;
        RECT 508.650 615.750 510.450 618.600 ;
        RECT 542.700 615.750 544.500 618.600 ;
        RECT 546.000 615.750 547.800 619.950 ;
        RECT 550.200 615.750 552.000 621.600 ;
        RECT 584.400 618.600 585.600 626.850 ;
        RECT 586.950 625.050 589.050 627.150 ;
        RECT 617.700 624.300 618.900 641.400 ;
        RECT 621.150 635.400 622.950 647.250 ;
        RECT 624.150 635.400 625.950 647.250 ;
        RECT 657.300 635.400 659.100 647.250 ;
        RECT 661.500 635.400 663.300 647.250 ;
        RECT 664.800 641.400 666.600 647.250 ;
        RECT 697.650 641.400 699.450 647.250 ;
        RECT 700.650 641.400 702.450 647.250 ;
        RECT 733.650 641.400 735.450 647.250 ;
        RECT 736.650 641.400 738.450 647.250 ;
        RECT 619.950 629.850 622.050 631.950 ;
        RECT 624.150 630.150 625.350 635.400 ;
        RECT 656.100 630.150 657.900 631.950 ;
        RECT 661.950 630.150 663.150 635.400 ;
        RECT 664.950 633.150 666.750 634.950 ;
        RECT 664.950 631.050 667.050 633.150 ;
        RECT 620.100 628.050 621.900 629.850 ;
        RECT 622.950 628.050 625.350 630.150 ;
        RECT 655.950 628.050 658.050 630.150 ;
        RECT 614.550 623.100 622.050 624.300 ;
        RECT 583.650 615.750 585.450 618.600 ;
        RECT 586.650 615.750 588.450 618.600 ;
        RECT 614.550 615.750 616.350 623.100 ;
        RECT 620.250 622.500 622.050 623.100 ;
        RECT 624.150 621.600 625.350 628.050 ;
        RECT 658.950 626.850 661.050 628.950 ;
        RECT 661.950 628.050 664.050 630.150 ;
        RECT 698.400 628.950 699.600 641.400 ;
        RECT 734.400 628.950 735.600 641.400 ;
        RECT 659.100 625.050 660.900 626.850 ;
        RECT 662.850 624.750 664.050 628.050 ;
        RECT 697.950 626.850 700.050 628.950 ;
        RECT 701.100 627.150 702.900 628.950 ;
        RECT 663.000 623.700 666.750 624.750 ;
        RECT 619.050 615.750 620.850 621.600 ;
        RECT 622.050 620.100 625.350 621.600 ;
        RECT 656.550 620.700 664.350 622.050 ;
        RECT 622.050 615.750 623.850 620.100 ;
        RECT 656.550 615.750 658.350 620.700 ;
        RECT 659.550 615.750 661.350 619.800 ;
        RECT 662.550 615.750 664.350 620.700 ;
        RECT 665.550 621.600 666.750 623.700 ;
        RECT 665.550 615.750 667.350 621.600 ;
        RECT 698.400 618.600 699.600 626.850 ;
        RECT 700.950 625.050 703.050 627.150 ;
        RECT 733.950 626.850 736.050 628.950 ;
        RECT 737.100 627.150 738.900 628.950 ;
        RECT 734.400 618.600 735.600 626.850 ;
        RECT 736.950 625.050 739.050 627.150 ;
        RECT 697.650 615.750 699.450 618.600 ;
        RECT 700.650 615.750 702.450 618.600 ;
        RECT 733.650 615.750 735.450 618.600 ;
        RECT 736.650 615.750 738.450 618.600 ;
        RECT 31.650 608.400 33.450 611.250 ;
        RECT 34.650 608.400 36.450 611.250 ;
        RECT 37.650 608.400 39.450 611.250 ;
        RECT 34.950 601.950 36.000 608.400 ;
        RECT 41.550 605.400 43.350 611.250 ;
        RECT 44.850 608.400 46.650 611.250 ;
        RECT 49.350 608.400 51.150 611.250 ;
        RECT 53.550 608.400 55.350 611.250 ;
        RECT 57.450 608.400 59.250 611.250 ;
        RECT 60.750 608.400 62.550 611.250 ;
        RECT 65.250 609.300 67.050 611.250 ;
        RECT 65.250 608.400 69.000 609.300 ;
        RECT 70.050 608.400 71.850 611.250 ;
        RECT 49.650 607.500 50.700 608.400 ;
        RECT 46.950 606.300 50.700 607.500 ;
        RECT 58.200 606.600 59.250 608.400 ;
        RECT 67.950 607.500 69.000 608.400 ;
        RECT 46.950 605.400 49.050 606.300 ;
        RECT 41.550 603.150 42.750 605.400 ;
        RECT 54.150 604.200 55.950 606.000 ;
        RECT 58.200 605.550 63.150 606.600 ;
        RECT 61.350 604.800 63.150 605.550 ;
        RECT 64.650 604.800 66.450 606.600 ;
        RECT 67.950 605.400 70.050 607.500 ;
        RECT 73.050 605.400 74.850 611.250 ;
        RECT 55.050 603.900 55.950 604.200 ;
        RECT 65.100 603.900 66.150 604.800 ;
        RECT 34.950 599.850 37.050 601.950 ;
        RECT 41.550 601.050 46.050 603.150 ;
        RECT 55.050 603.000 66.150 603.900 ;
        RECT 31.950 596.850 34.050 598.950 ;
        RECT 32.100 595.050 33.900 596.850 ;
        RECT 34.950 592.650 36.000 599.850 ;
        RECT 37.950 596.850 40.050 598.950 ;
        RECT 38.100 595.050 39.900 596.850 ;
        RECT 33.450 591.600 36.000 592.650 ;
        RECT 41.550 591.600 42.750 601.050 ;
        RECT 43.950 599.250 47.850 601.050 ;
        RECT 43.950 598.950 46.050 599.250 ;
        RECT 55.050 598.950 55.950 603.000 ;
        RECT 65.100 601.800 66.150 603.000 ;
        RECT 65.100 600.600 72.000 601.800 ;
        RECT 65.100 600.000 66.900 600.600 ;
        RECT 71.100 599.850 72.000 600.600 ;
        RECT 68.100 598.950 69.900 599.700 ;
        RECT 55.050 596.850 58.050 598.950 ;
        RECT 61.950 597.900 69.900 598.950 ;
        RECT 71.100 598.050 72.900 599.850 ;
        RECT 61.950 596.850 64.050 597.900 ;
        RECT 43.950 593.400 45.750 595.200 ;
        RECT 44.850 592.200 49.050 593.400 ;
        RECT 55.050 592.200 55.950 596.850 ;
        RECT 63.750 593.100 65.550 593.400 ;
        RECT 33.450 579.750 35.250 591.600 ;
        RECT 37.650 579.750 39.450 591.600 ;
        RECT 41.550 579.750 43.350 591.600 ;
        RECT 46.950 591.300 49.050 592.200 ;
        RECT 49.950 591.300 55.950 592.200 ;
        RECT 57.150 592.800 65.550 593.100 ;
        RECT 73.950 592.800 74.850 605.400 ;
        RECT 57.150 592.200 74.850 592.800 ;
        RECT 49.950 590.400 50.850 591.300 ;
        RECT 48.150 588.600 50.850 590.400 ;
        RECT 51.750 590.100 53.550 590.400 ;
        RECT 57.150 590.100 58.050 592.200 ;
        RECT 63.750 591.600 74.850 592.200 ;
        RECT 51.750 589.200 58.050 590.100 ;
        RECT 58.950 590.700 60.750 591.300 ;
        RECT 58.950 589.500 66.450 590.700 ;
        RECT 51.750 588.600 53.550 589.200 ;
        RECT 65.250 588.600 66.450 589.500 ;
        RECT 46.950 585.600 50.850 587.700 ;
        RECT 55.950 586.500 62.850 588.300 ;
        RECT 65.250 586.500 70.050 588.600 ;
        RECT 44.550 579.750 46.350 582.600 ;
        RECT 49.050 579.750 50.850 585.600 ;
        RECT 53.250 579.750 55.050 585.600 ;
        RECT 57.150 579.750 58.950 586.500 ;
        RECT 65.250 585.600 66.450 586.500 ;
        RECT 60.150 579.750 61.950 585.600 ;
        RECT 64.950 579.750 66.750 585.600 ;
        RECT 70.050 579.750 71.850 585.600 ;
        RECT 73.050 579.750 74.850 591.600 ;
        RECT 78.150 605.400 79.950 611.250 ;
        RECT 81.150 608.400 82.950 611.250 ;
        RECT 85.950 609.300 87.750 611.250 ;
        RECT 84.000 608.400 87.750 609.300 ;
        RECT 90.450 608.400 92.250 611.250 ;
        RECT 93.750 608.400 95.550 611.250 ;
        RECT 97.650 608.400 99.450 611.250 ;
        RECT 101.850 608.400 103.650 611.250 ;
        RECT 106.350 608.400 108.150 611.250 ;
        RECT 84.000 607.500 85.050 608.400 ;
        RECT 82.950 605.400 85.050 607.500 ;
        RECT 93.750 606.600 94.800 608.400 ;
        RECT 78.150 592.800 79.050 605.400 ;
        RECT 86.550 604.800 88.350 606.600 ;
        RECT 89.850 605.550 94.800 606.600 ;
        RECT 102.300 607.500 103.350 608.400 ;
        RECT 102.300 606.300 106.050 607.500 ;
        RECT 89.850 604.800 91.650 605.550 ;
        RECT 86.850 603.900 87.900 604.800 ;
        RECT 97.050 604.200 98.850 606.000 ;
        RECT 103.950 605.400 106.050 606.300 ;
        RECT 109.650 605.400 111.450 611.250 ;
        RECT 140.550 608.400 142.350 611.250 ;
        RECT 143.550 608.400 145.350 611.250 ;
        RECT 176.700 608.400 178.500 611.250 ;
        RECT 97.050 603.900 97.950 604.200 ;
        RECT 86.850 603.000 97.950 603.900 ;
        RECT 110.250 603.150 111.450 605.400 ;
        RECT 86.850 601.800 87.900 603.000 ;
        RECT 81.000 600.600 87.900 601.800 ;
        RECT 81.000 599.850 81.900 600.600 ;
        RECT 86.100 600.000 87.900 600.600 ;
        RECT 80.100 598.050 81.900 599.850 ;
        RECT 83.100 598.950 84.900 599.700 ;
        RECT 97.050 598.950 97.950 603.000 ;
        RECT 106.950 601.050 111.450 603.150 ;
        RECT 105.150 599.250 109.050 601.050 ;
        RECT 106.950 598.950 109.050 599.250 ;
        RECT 83.100 597.900 91.050 598.950 ;
        RECT 88.950 596.850 91.050 597.900 ;
        RECT 94.950 596.850 97.950 598.950 ;
        RECT 87.450 593.100 89.250 593.400 ;
        RECT 87.450 592.800 95.850 593.100 ;
        RECT 78.150 592.200 95.850 592.800 ;
        RECT 78.150 591.600 89.250 592.200 ;
        RECT 78.150 579.750 79.950 591.600 ;
        RECT 92.250 590.700 94.050 591.300 ;
        RECT 86.550 589.500 94.050 590.700 ;
        RECT 94.950 590.100 95.850 592.200 ;
        RECT 97.050 592.200 97.950 596.850 ;
        RECT 107.250 593.400 109.050 595.200 ;
        RECT 103.950 592.200 108.150 593.400 ;
        RECT 97.050 591.300 103.050 592.200 ;
        RECT 103.950 591.300 106.050 592.200 ;
        RECT 110.250 591.600 111.450 601.050 ;
        RECT 139.950 599.850 142.050 601.950 ;
        RECT 143.400 600.150 144.600 608.400 ;
        RECT 180.000 607.050 181.800 611.250 ;
        RECT 176.100 605.400 181.800 607.050 ;
        RECT 184.200 605.400 186.000 611.250 ;
        RECT 189.150 605.400 190.950 611.250 ;
        RECT 192.150 608.400 193.950 611.250 ;
        RECT 196.950 609.300 198.750 611.250 ;
        RECT 195.000 608.400 198.750 609.300 ;
        RECT 201.450 608.400 203.250 611.250 ;
        RECT 204.750 608.400 206.550 611.250 ;
        RECT 208.650 608.400 210.450 611.250 ;
        RECT 212.850 608.400 214.650 611.250 ;
        RECT 217.350 608.400 219.150 611.250 ;
        RECT 195.000 607.500 196.050 608.400 ;
        RECT 193.950 605.400 196.050 607.500 ;
        RECT 204.750 606.600 205.800 608.400 ;
        RECT 140.100 598.050 141.900 599.850 ;
        RECT 142.950 598.050 145.050 600.150 ;
        RECT 176.100 598.950 177.300 605.400 ;
        RECT 179.100 600.150 180.900 601.950 ;
        RECT 102.150 590.400 103.050 591.300 ;
        RECT 99.450 590.100 101.250 590.400 ;
        RECT 86.550 588.600 87.750 589.500 ;
        RECT 94.950 589.200 101.250 590.100 ;
        RECT 99.450 588.600 101.250 589.200 ;
        RECT 102.150 588.600 104.850 590.400 ;
        RECT 82.950 586.500 87.750 588.600 ;
        RECT 90.150 586.500 97.050 588.300 ;
        RECT 86.550 585.600 87.750 586.500 ;
        RECT 81.150 579.750 82.950 585.600 ;
        RECT 86.250 579.750 88.050 585.600 ;
        RECT 91.050 579.750 92.850 585.600 ;
        RECT 94.050 579.750 95.850 586.500 ;
        RECT 102.150 585.600 106.050 587.700 ;
        RECT 97.950 579.750 99.750 585.600 ;
        RECT 102.150 579.750 103.950 585.600 ;
        RECT 106.650 579.750 108.450 582.600 ;
        RECT 109.650 579.750 111.450 591.600 ;
        RECT 143.400 585.600 144.600 598.050 ;
        RECT 175.950 596.850 178.050 598.950 ;
        RECT 178.950 598.050 181.050 600.150 ;
        RECT 181.950 599.850 184.050 601.950 ;
        RECT 185.100 600.150 186.900 601.950 ;
        RECT 182.100 598.050 183.900 599.850 ;
        RECT 184.950 598.050 187.050 600.150 ;
        RECT 176.100 591.600 177.300 596.850 ;
        RECT 189.150 592.800 190.050 605.400 ;
        RECT 197.550 604.800 199.350 606.600 ;
        RECT 200.850 605.550 205.800 606.600 ;
        RECT 213.300 607.500 214.350 608.400 ;
        RECT 213.300 606.300 217.050 607.500 ;
        RECT 200.850 604.800 202.650 605.550 ;
        RECT 197.850 603.900 198.900 604.800 ;
        RECT 208.050 604.200 209.850 606.000 ;
        RECT 214.950 605.400 217.050 606.300 ;
        RECT 220.650 605.400 222.450 611.250 ;
        RECT 254.700 608.400 256.500 611.250 ;
        RECT 258.000 607.050 259.800 611.250 ;
        RECT 208.050 603.900 208.950 604.200 ;
        RECT 197.850 603.000 208.950 603.900 ;
        RECT 221.250 603.150 222.450 605.400 ;
        RECT 197.850 601.800 198.900 603.000 ;
        RECT 192.000 600.600 198.900 601.800 ;
        RECT 192.000 599.850 192.900 600.600 ;
        RECT 197.100 600.000 198.900 600.600 ;
        RECT 191.100 598.050 192.900 599.850 ;
        RECT 194.100 598.950 195.900 599.700 ;
        RECT 208.050 598.950 208.950 603.000 ;
        RECT 217.950 601.050 222.450 603.150 ;
        RECT 216.150 599.250 220.050 601.050 ;
        RECT 217.950 598.950 220.050 599.250 ;
        RECT 194.100 597.900 202.050 598.950 ;
        RECT 199.950 596.850 202.050 597.900 ;
        RECT 205.950 596.850 208.950 598.950 ;
        RECT 198.450 593.100 200.250 593.400 ;
        RECT 198.450 592.800 206.850 593.100 ;
        RECT 189.150 592.200 206.850 592.800 ;
        RECT 189.150 591.600 200.250 592.200 ;
        RECT 140.550 579.750 142.350 585.600 ;
        RECT 143.550 579.750 145.350 585.600 ;
        RECT 175.650 579.750 177.450 591.600 ;
        RECT 178.650 590.700 186.450 591.600 ;
        RECT 178.650 579.750 180.450 590.700 ;
        RECT 181.650 579.750 183.450 589.800 ;
        RECT 184.650 579.750 186.450 590.700 ;
        RECT 189.150 579.750 190.950 591.600 ;
        RECT 203.250 590.700 205.050 591.300 ;
        RECT 197.550 589.500 205.050 590.700 ;
        RECT 205.950 590.100 206.850 592.200 ;
        RECT 208.050 592.200 208.950 596.850 ;
        RECT 218.250 593.400 220.050 595.200 ;
        RECT 214.950 592.200 219.150 593.400 ;
        RECT 208.050 591.300 214.050 592.200 ;
        RECT 214.950 591.300 217.050 592.200 ;
        RECT 221.250 591.600 222.450 601.050 ;
        RECT 254.100 605.400 259.800 607.050 ;
        RECT 262.200 605.400 264.000 611.250 ;
        RECT 254.100 598.950 255.300 605.400 ;
        RECT 299.100 603.000 300.900 611.250 ;
        RECT 257.100 600.150 258.900 601.950 ;
        RECT 253.950 596.850 256.050 598.950 ;
        RECT 256.950 598.050 259.050 600.150 ;
        RECT 259.950 599.850 262.050 601.950 ;
        RECT 263.100 600.150 264.900 601.950 ;
        RECT 296.400 601.350 300.900 603.000 ;
        RECT 304.500 602.400 306.300 611.250 ;
        RECT 335.700 608.400 337.500 611.250 ;
        RECT 339.000 607.050 340.800 611.250 ;
        RECT 335.100 605.400 340.800 607.050 ;
        RECT 343.200 605.400 345.000 611.250 ;
        RECT 374.850 605.400 376.650 611.250 ;
        RECT 260.100 598.050 261.900 599.850 ;
        RECT 262.950 598.050 265.050 600.150 ;
        RECT 296.400 597.150 297.600 601.350 ;
        RECT 335.100 598.950 336.300 605.400 ;
        RECT 379.350 604.200 381.150 611.250 ;
        RECT 377.550 603.300 381.150 604.200 ;
        RECT 413.550 603.900 415.350 611.250 ;
        RECT 418.050 605.400 419.850 611.250 ;
        RECT 421.050 606.900 422.850 611.250 ;
        RECT 421.050 605.400 424.350 606.900 ;
        RECT 419.250 603.900 421.050 604.500 ;
        RECT 338.100 600.150 339.900 601.950 ;
        RECT 254.100 591.600 255.300 596.850 ;
        RECT 295.950 595.050 298.050 597.150 ;
        RECT 334.950 596.850 337.050 598.950 ;
        RECT 337.950 598.050 340.050 600.150 ;
        RECT 340.950 599.850 343.050 601.950 ;
        RECT 344.100 600.150 345.900 601.950 ;
        RECT 341.100 598.050 342.900 599.850 ;
        RECT 343.950 598.050 346.050 600.150 ;
        RECT 374.100 597.150 375.900 598.950 ;
        RECT 213.150 590.400 214.050 591.300 ;
        RECT 210.450 590.100 212.250 590.400 ;
        RECT 197.550 588.600 198.750 589.500 ;
        RECT 205.950 589.200 212.250 590.100 ;
        RECT 210.450 588.600 212.250 589.200 ;
        RECT 213.150 588.600 215.850 590.400 ;
        RECT 193.950 586.500 198.750 588.600 ;
        RECT 201.150 586.500 208.050 588.300 ;
        RECT 197.550 585.600 198.750 586.500 ;
        RECT 192.150 579.750 193.950 585.600 ;
        RECT 197.250 579.750 199.050 585.600 ;
        RECT 202.050 579.750 203.850 585.600 ;
        RECT 205.050 579.750 206.850 586.500 ;
        RECT 213.150 585.600 217.050 587.700 ;
        RECT 208.950 579.750 210.750 585.600 ;
        RECT 213.150 579.750 214.950 585.600 ;
        RECT 217.650 579.750 219.450 582.600 ;
        RECT 220.650 579.750 222.450 591.600 ;
        RECT 253.650 579.750 255.450 591.600 ;
        RECT 256.650 590.700 264.450 591.600 ;
        RECT 256.650 579.750 258.450 590.700 ;
        RECT 259.650 579.750 261.450 589.800 ;
        RECT 262.650 579.750 264.450 590.700 ;
        RECT 296.250 586.800 297.300 595.050 ;
        RECT 298.950 593.850 301.050 595.950 ;
        RECT 304.950 593.850 307.050 595.950 ;
        RECT 298.950 592.050 300.750 593.850 ;
        RECT 301.950 590.850 304.050 592.950 ;
        RECT 305.100 592.050 306.900 593.850 ;
        RECT 335.100 591.600 336.300 596.850 ;
        RECT 373.950 595.050 376.050 597.150 ;
        RECT 377.550 595.950 378.750 603.300 ;
        RECT 413.550 602.700 421.050 603.900 ;
        RECT 380.100 597.150 381.900 598.950 ;
        RECT 376.950 593.850 379.050 595.950 ;
        RECT 379.950 595.050 382.050 597.150 ;
        RECT 412.950 596.850 415.050 598.950 ;
        RECT 413.100 595.050 414.900 596.850 ;
        RECT 302.100 589.050 303.900 590.850 ;
        RECT 296.250 585.900 303.300 586.800 ;
        RECT 296.250 585.600 297.450 585.900 ;
        RECT 295.650 579.750 297.450 585.600 ;
        RECT 301.650 585.600 303.300 585.900 ;
        RECT 298.650 579.750 300.450 585.000 ;
        RECT 301.650 579.750 303.450 585.600 ;
        RECT 304.650 579.750 306.450 585.600 ;
        RECT 334.650 579.750 336.450 591.600 ;
        RECT 337.650 590.700 345.450 591.600 ;
        RECT 337.650 579.750 339.450 590.700 ;
        RECT 340.650 579.750 342.450 589.800 ;
        RECT 343.650 579.750 345.450 590.700 ;
        RECT 377.550 585.600 378.750 593.850 ;
        RECT 416.700 585.600 417.900 602.700 ;
        RECT 423.150 598.950 424.350 605.400 ;
        RECT 461.100 603.000 462.900 611.250 ;
        RECT 419.100 597.150 420.900 598.950 ;
        RECT 418.950 595.050 421.050 597.150 ;
        RECT 421.950 596.850 424.350 598.950 ;
        RECT 458.400 601.350 462.900 603.000 ;
        RECT 466.500 602.400 468.300 611.250 ;
        RECT 498.000 605.400 499.800 611.250 ;
        RECT 502.200 607.050 504.000 611.250 ;
        RECT 505.500 608.400 507.300 611.250 ;
        RECT 502.200 605.400 507.900 607.050 ;
        RECT 458.400 597.150 459.600 601.350 ;
        RECT 497.100 600.150 498.900 601.950 ;
        RECT 496.950 598.050 499.050 600.150 ;
        RECT 499.950 599.850 502.050 601.950 ;
        RECT 503.100 600.150 504.900 601.950 ;
        RECT 500.100 598.050 501.900 599.850 ;
        RECT 502.950 598.050 505.050 600.150 ;
        RECT 506.700 598.950 507.900 605.400 ;
        RECT 513.150 605.400 514.950 611.250 ;
        RECT 516.150 608.400 517.950 611.250 ;
        RECT 520.950 609.300 522.750 611.250 ;
        RECT 519.000 608.400 522.750 609.300 ;
        RECT 525.450 608.400 527.250 611.250 ;
        RECT 528.750 608.400 530.550 611.250 ;
        RECT 532.650 608.400 534.450 611.250 ;
        RECT 536.850 608.400 538.650 611.250 ;
        RECT 541.350 608.400 543.150 611.250 ;
        RECT 519.000 607.500 520.050 608.400 ;
        RECT 517.950 605.400 520.050 607.500 ;
        RECT 528.750 606.600 529.800 608.400 ;
        RECT 423.150 591.600 424.350 596.850 ;
        RECT 457.950 595.050 460.050 597.150 ;
        RECT 505.950 596.850 508.050 598.950 ;
        RECT 374.550 579.750 376.350 585.600 ;
        RECT 377.550 579.750 379.350 585.600 ;
        RECT 380.550 579.750 382.350 585.600 ;
        RECT 413.550 579.750 415.350 585.600 ;
        RECT 416.550 579.750 418.350 585.600 ;
        RECT 420.150 579.750 421.950 591.600 ;
        RECT 423.150 579.750 424.950 591.600 ;
        RECT 458.250 586.800 459.300 595.050 ;
        RECT 460.950 593.850 463.050 595.950 ;
        RECT 466.950 593.850 469.050 595.950 ;
        RECT 460.950 592.050 462.750 593.850 ;
        RECT 463.950 590.850 466.050 592.950 ;
        RECT 467.100 592.050 468.900 593.850 ;
        RECT 506.700 591.600 507.900 596.850 ;
        RECT 513.150 592.800 514.050 605.400 ;
        RECT 521.550 604.800 523.350 606.600 ;
        RECT 524.850 605.550 529.800 606.600 ;
        RECT 537.300 607.500 538.350 608.400 ;
        RECT 537.300 606.300 541.050 607.500 ;
        RECT 524.850 604.800 526.650 605.550 ;
        RECT 521.850 603.900 522.900 604.800 ;
        RECT 532.050 604.200 533.850 606.000 ;
        RECT 538.950 605.400 541.050 606.300 ;
        RECT 544.650 605.400 546.450 611.250 ;
        RECT 575.550 608.400 577.350 611.250 ;
        RECT 578.550 608.400 580.350 611.250 ;
        RECT 581.550 608.400 583.350 611.250 ;
        RECT 532.050 603.900 532.950 604.200 ;
        RECT 521.850 603.000 532.950 603.900 ;
        RECT 545.250 603.150 546.450 605.400 ;
        RECT 521.850 601.800 522.900 603.000 ;
        RECT 516.000 600.600 522.900 601.800 ;
        RECT 516.000 599.850 516.900 600.600 ;
        RECT 521.100 600.000 522.900 600.600 ;
        RECT 515.100 598.050 516.900 599.850 ;
        RECT 518.100 598.950 519.900 599.700 ;
        RECT 532.050 598.950 532.950 603.000 ;
        RECT 541.950 601.050 546.450 603.150 ;
        RECT 579.000 601.950 580.050 608.400 ;
        RECT 540.150 599.250 544.050 601.050 ;
        RECT 541.950 598.950 544.050 599.250 ;
        RECT 518.100 597.900 526.050 598.950 ;
        RECT 523.950 596.850 526.050 597.900 ;
        RECT 529.950 596.850 532.950 598.950 ;
        RECT 522.450 593.100 524.250 593.400 ;
        RECT 522.450 592.800 530.850 593.100 ;
        RECT 513.150 592.200 530.850 592.800 ;
        RECT 513.150 591.600 524.250 592.200 ;
        RECT 464.100 589.050 465.900 590.850 ;
        RECT 497.550 590.700 505.350 591.600 ;
        RECT 458.250 585.900 465.300 586.800 ;
        RECT 458.250 585.600 459.450 585.900 ;
        RECT 457.650 579.750 459.450 585.600 ;
        RECT 463.650 585.600 465.300 585.900 ;
        RECT 460.650 579.750 462.450 585.000 ;
        RECT 463.650 579.750 465.450 585.600 ;
        RECT 466.650 579.750 468.450 585.600 ;
        RECT 497.550 579.750 499.350 590.700 ;
        RECT 500.550 579.750 502.350 589.800 ;
        RECT 503.550 579.750 505.350 590.700 ;
        RECT 506.550 579.750 508.350 591.600 ;
        RECT 513.150 579.750 514.950 591.600 ;
        RECT 527.250 590.700 529.050 591.300 ;
        RECT 521.550 589.500 529.050 590.700 ;
        RECT 529.950 590.100 530.850 592.200 ;
        RECT 532.050 592.200 532.950 596.850 ;
        RECT 542.250 593.400 544.050 595.200 ;
        RECT 538.950 592.200 543.150 593.400 ;
        RECT 532.050 591.300 538.050 592.200 ;
        RECT 538.950 591.300 541.050 592.200 ;
        RECT 545.250 591.600 546.450 601.050 ;
        RECT 577.950 599.850 580.050 601.950 ;
        RECT 574.950 596.850 577.050 598.950 ;
        RECT 575.100 595.050 576.900 596.850 ;
        RECT 579.000 592.650 580.050 599.850 ;
        RECT 588.150 605.400 589.950 611.250 ;
        RECT 591.150 608.400 592.950 611.250 ;
        RECT 595.950 609.300 597.750 611.250 ;
        RECT 594.000 608.400 597.750 609.300 ;
        RECT 600.450 608.400 602.250 611.250 ;
        RECT 603.750 608.400 605.550 611.250 ;
        RECT 607.650 608.400 609.450 611.250 ;
        RECT 611.850 608.400 613.650 611.250 ;
        RECT 616.350 608.400 618.150 611.250 ;
        RECT 594.000 607.500 595.050 608.400 ;
        RECT 592.950 605.400 595.050 607.500 ;
        RECT 603.750 606.600 604.800 608.400 ;
        RECT 580.950 596.850 583.050 598.950 ;
        RECT 581.100 595.050 582.900 596.850 ;
        RECT 588.150 592.800 589.050 605.400 ;
        RECT 596.550 604.800 598.350 606.600 ;
        RECT 599.850 605.550 604.800 606.600 ;
        RECT 612.300 607.500 613.350 608.400 ;
        RECT 612.300 606.300 616.050 607.500 ;
        RECT 599.850 604.800 601.650 605.550 ;
        RECT 596.850 603.900 597.900 604.800 ;
        RECT 607.050 604.200 608.850 606.000 ;
        RECT 613.950 605.400 616.050 606.300 ;
        RECT 619.650 605.400 621.450 611.250 ;
        RECT 607.050 603.900 607.950 604.200 ;
        RECT 596.850 603.000 607.950 603.900 ;
        RECT 620.250 603.150 621.450 605.400 ;
        RECT 653.850 604.200 655.650 611.250 ;
        RECT 658.350 605.400 660.150 611.250 ;
        RECT 692.850 604.200 694.650 611.250 ;
        RECT 697.350 605.400 699.150 611.250 ;
        RECT 725.550 608.400 727.350 611.250 ;
        RECT 728.550 608.400 730.350 611.250 ;
        RECT 731.550 608.400 733.350 611.250 ;
        RECT 653.850 603.300 657.450 604.200 ;
        RECT 692.850 603.300 696.450 604.200 ;
        RECT 596.850 601.800 597.900 603.000 ;
        RECT 591.000 600.600 597.900 601.800 ;
        RECT 591.000 599.850 591.900 600.600 ;
        RECT 596.100 600.000 597.900 600.600 ;
        RECT 590.100 598.050 591.900 599.850 ;
        RECT 593.100 598.950 594.900 599.700 ;
        RECT 607.050 598.950 607.950 603.000 ;
        RECT 616.950 601.050 621.450 603.150 ;
        RECT 615.150 599.250 619.050 601.050 ;
        RECT 616.950 598.950 619.050 599.250 ;
        RECT 593.100 597.900 601.050 598.950 ;
        RECT 598.950 596.850 601.050 597.900 ;
        RECT 604.950 596.850 607.950 598.950 ;
        RECT 597.450 593.100 599.250 593.400 ;
        RECT 597.450 592.800 605.850 593.100 ;
        RECT 579.000 591.600 581.550 592.650 ;
        RECT 537.150 590.400 538.050 591.300 ;
        RECT 534.450 590.100 536.250 590.400 ;
        RECT 521.550 588.600 522.750 589.500 ;
        RECT 529.950 589.200 536.250 590.100 ;
        RECT 534.450 588.600 536.250 589.200 ;
        RECT 537.150 588.600 539.850 590.400 ;
        RECT 517.950 586.500 522.750 588.600 ;
        RECT 525.150 586.500 532.050 588.300 ;
        RECT 521.550 585.600 522.750 586.500 ;
        RECT 516.150 579.750 517.950 585.600 ;
        RECT 521.250 579.750 523.050 585.600 ;
        RECT 526.050 579.750 527.850 585.600 ;
        RECT 529.050 579.750 530.850 586.500 ;
        RECT 537.150 585.600 541.050 587.700 ;
        RECT 532.950 579.750 534.750 585.600 ;
        RECT 537.150 579.750 538.950 585.600 ;
        RECT 541.650 579.750 543.450 582.600 ;
        RECT 544.650 579.750 546.450 591.600 ;
        RECT 575.550 579.750 577.350 591.600 ;
        RECT 579.750 579.750 581.550 591.600 ;
        RECT 588.150 592.200 605.850 592.800 ;
        RECT 588.150 591.600 599.250 592.200 ;
        RECT 588.150 579.750 589.950 591.600 ;
        RECT 602.250 590.700 604.050 591.300 ;
        RECT 596.550 589.500 604.050 590.700 ;
        RECT 604.950 590.100 605.850 592.200 ;
        RECT 607.050 592.200 607.950 596.850 ;
        RECT 617.250 593.400 619.050 595.200 ;
        RECT 613.950 592.200 618.150 593.400 ;
        RECT 607.050 591.300 613.050 592.200 ;
        RECT 613.950 591.300 616.050 592.200 ;
        RECT 620.250 591.600 621.450 601.050 ;
        RECT 653.100 597.150 654.900 598.950 ;
        RECT 652.950 595.050 655.050 597.150 ;
        RECT 656.250 595.950 657.450 603.300 ;
        RECT 659.100 597.150 660.900 598.950 ;
        RECT 692.100 597.150 693.900 598.950 ;
        RECT 655.950 593.850 658.050 595.950 ;
        RECT 658.950 595.050 661.050 597.150 ;
        RECT 691.950 595.050 694.050 597.150 ;
        RECT 695.250 595.950 696.450 603.300 ;
        RECT 729.000 601.950 730.050 608.400 ;
        RECT 727.950 599.850 730.050 601.950 ;
        RECT 698.100 597.150 699.900 598.950 ;
        RECT 694.950 593.850 697.050 595.950 ;
        RECT 697.950 595.050 700.050 597.150 ;
        RECT 724.950 596.850 727.050 598.950 ;
        RECT 725.100 595.050 726.900 596.850 ;
        RECT 612.150 590.400 613.050 591.300 ;
        RECT 609.450 590.100 611.250 590.400 ;
        RECT 596.550 588.600 597.750 589.500 ;
        RECT 604.950 589.200 611.250 590.100 ;
        RECT 609.450 588.600 611.250 589.200 ;
        RECT 612.150 588.600 614.850 590.400 ;
        RECT 592.950 586.500 597.750 588.600 ;
        RECT 600.150 586.500 607.050 588.300 ;
        RECT 596.550 585.600 597.750 586.500 ;
        RECT 591.150 579.750 592.950 585.600 ;
        RECT 596.250 579.750 598.050 585.600 ;
        RECT 601.050 579.750 602.850 585.600 ;
        RECT 604.050 579.750 605.850 586.500 ;
        RECT 612.150 585.600 616.050 587.700 ;
        RECT 607.950 579.750 609.750 585.600 ;
        RECT 612.150 579.750 613.950 585.600 ;
        RECT 616.650 579.750 618.450 582.600 ;
        RECT 619.650 579.750 621.450 591.600 ;
        RECT 656.250 585.600 657.450 593.850 ;
        RECT 695.250 585.600 696.450 593.850 ;
        RECT 729.000 592.650 730.050 599.850 ;
        RECT 730.950 596.850 733.050 598.950 ;
        RECT 731.100 595.050 732.900 596.850 ;
        RECT 729.000 591.600 731.550 592.650 ;
        RECT 652.650 579.750 654.450 585.600 ;
        RECT 655.650 579.750 657.450 585.600 ;
        RECT 658.650 579.750 660.450 585.600 ;
        RECT 691.650 579.750 693.450 585.600 ;
        RECT 694.650 579.750 696.450 585.600 ;
        RECT 697.650 579.750 699.450 585.600 ;
        RECT 725.550 579.750 727.350 591.600 ;
        RECT 729.750 579.750 731.550 591.600 ;
        RECT 31.050 563.400 32.850 575.250 ;
        RECT 34.050 563.400 35.850 575.250 ;
        RECT 37.650 569.400 39.450 575.250 ;
        RECT 40.650 569.400 42.450 575.250 ;
        RECT 31.650 558.150 32.850 563.400 ;
        RECT 31.650 556.050 34.050 558.150 ;
        RECT 34.950 557.850 37.050 559.950 ;
        RECT 35.100 556.050 36.900 557.850 ;
        RECT 31.650 549.600 32.850 556.050 ;
        RECT 38.100 552.300 39.300 569.400 ;
        RECT 71.550 563.400 73.350 575.250 ;
        RECT 75.750 563.400 77.550 575.250 ;
        RECT 112.650 563.400 114.450 575.250 ;
        RECT 115.650 564.300 117.450 575.250 ;
        RECT 118.650 565.200 120.450 575.250 ;
        RECT 121.650 564.300 123.450 575.250 ;
        RECT 152.550 569.400 154.350 575.250 ;
        RECT 155.550 569.400 157.350 575.250 ;
        RECT 158.550 569.400 160.350 575.250 ;
        RECT 115.650 563.400 123.450 564.300 ;
        RECT 75.000 562.350 77.550 563.400 ;
        RECT 41.100 558.150 42.900 559.950 ;
        RECT 71.100 558.150 72.900 559.950 ;
        RECT 40.950 556.050 43.050 558.150 ;
        RECT 70.950 556.050 73.050 558.150 ;
        RECT 75.000 555.150 76.050 562.350 ;
        RECT 77.100 558.150 78.900 559.950 ;
        RECT 113.100 558.150 114.300 563.400 ;
        RECT 155.550 561.150 156.750 569.400 ;
        RECT 191.550 563.400 193.350 575.250 ;
        RECT 194.550 562.500 196.350 575.250 ;
        RECT 197.550 563.400 199.350 575.250 ;
        RECT 200.550 562.500 202.350 575.250 ;
        RECT 203.550 563.400 205.350 575.250 ;
        RECT 206.550 562.500 208.350 575.250 ;
        RECT 209.550 563.400 211.350 575.250 ;
        RECT 212.550 562.500 214.350 575.250 ;
        RECT 215.550 563.400 217.350 575.250 ;
        RECT 249.300 563.400 251.100 575.250 ;
        RECT 253.500 563.400 255.300 575.250 ;
        RECT 256.800 569.400 258.600 575.250 ;
        RECT 290.550 563.400 292.350 575.250 ;
        RECT 194.550 561.300 198.450 562.500 ;
        RECT 200.550 561.300 204.300 562.500 ;
        RECT 206.550 561.300 210.300 562.500 ;
        RECT 212.550 561.300 215.250 562.500 ;
        RECT 76.950 556.050 79.050 558.150 ;
        RECT 112.950 556.050 115.050 558.150 ;
        RECT 151.950 557.850 154.050 559.950 ;
        RECT 154.950 559.050 157.050 561.150 ;
        RECT 73.950 553.050 76.050 555.150 ;
        RECT 34.950 551.100 42.450 552.300 ;
        RECT 34.950 550.500 36.750 551.100 ;
        RECT 31.650 548.100 34.950 549.600 ;
        RECT 33.150 543.750 34.950 548.100 ;
        RECT 36.150 543.750 37.950 549.600 ;
        RECT 40.650 543.750 42.450 551.100 ;
        RECT 75.000 546.600 76.050 553.050 ;
        RECT 113.100 549.600 114.300 556.050 ;
        RECT 115.950 554.850 118.050 556.950 ;
        RECT 119.100 555.150 120.900 556.950 ;
        RECT 116.100 553.050 117.900 554.850 ;
        RECT 118.950 553.050 121.050 555.150 ;
        RECT 121.950 554.850 124.050 556.950 ;
        RECT 152.100 556.050 153.900 557.850 ;
        RECT 122.100 553.050 123.900 554.850 ;
        RECT 155.550 551.700 156.750 559.050 ;
        RECT 157.950 557.850 160.050 559.950 ;
        RECT 158.100 556.050 159.900 557.850 ;
        RECT 193.950 554.850 196.050 556.950 ;
        RECT 194.100 553.050 195.900 554.850 ;
        RECT 197.250 554.400 198.450 561.300 ;
        RECT 203.100 554.400 204.300 561.300 ;
        RECT 209.100 554.400 210.300 561.300 ;
        RECT 214.200 556.950 215.250 561.300 ;
        RECT 248.100 558.150 249.900 559.950 ;
        RECT 253.950 558.150 255.150 563.400 ;
        RECT 256.950 561.150 258.750 562.950 ;
        RECT 293.550 562.500 295.350 575.250 ;
        RECT 296.550 563.400 298.350 575.250 ;
        RECT 299.550 562.500 301.350 575.250 ;
        RECT 302.550 563.400 304.350 575.250 ;
        RECT 305.550 562.500 307.350 575.250 ;
        RECT 308.550 563.400 310.350 575.250 ;
        RECT 311.550 562.500 313.350 575.250 ;
        RECT 314.550 563.400 316.350 575.250 ;
        RECT 347.550 569.400 349.350 575.250 ;
        RECT 350.550 569.400 352.350 575.250 ;
        RECT 353.550 569.400 355.350 575.250 ;
        RECT 293.550 561.300 297.450 562.500 ;
        RECT 299.550 561.300 303.300 562.500 ;
        RECT 305.550 561.300 309.300 562.500 ;
        RECT 311.550 561.300 314.250 562.500 ;
        RECT 256.950 559.050 259.050 561.150 ;
        RECT 214.200 554.850 217.050 556.950 ;
        RECT 247.950 556.050 250.050 558.150 ;
        RECT 250.950 554.850 253.050 556.950 ;
        RECT 253.950 556.050 256.050 558.150 ;
        RECT 197.250 552.600 201.300 554.400 ;
        RECT 203.100 552.600 207.300 554.400 ;
        RECT 209.100 552.600 213.300 554.400 ;
        RECT 197.250 551.700 198.450 552.600 ;
        RECT 203.100 551.700 204.300 552.600 ;
        RECT 209.100 551.700 210.300 552.600 ;
        RECT 214.200 551.700 215.250 554.850 ;
        RECT 251.100 553.050 252.900 554.850 ;
        RECT 254.850 552.750 256.050 556.050 ;
        RECT 292.950 554.850 295.050 556.950 ;
        RECT 293.100 553.050 294.900 554.850 ;
        RECT 296.250 554.400 297.450 561.300 ;
        RECT 302.100 554.400 303.300 561.300 ;
        RECT 308.100 554.400 309.300 561.300 ;
        RECT 313.200 556.950 314.250 561.300 ;
        RECT 350.550 561.150 351.750 569.400 ;
        RECT 383.550 563.400 385.350 575.250 ;
        RECT 387.750 563.400 389.550 575.250 ;
        RECT 422.550 569.400 424.350 575.250 ;
        RECT 425.550 569.400 427.350 575.250 ;
        RECT 460.650 569.400 462.450 575.250 ;
        RECT 463.650 570.000 465.450 575.250 ;
        RECT 387.000 562.350 389.550 563.400 ;
        RECT 346.950 557.850 349.050 559.950 ;
        RECT 349.950 559.050 352.050 561.150 ;
        RECT 313.200 554.850 316.050 556.950 ;
        RECT 347.100 556.050 348.900 557.850 ;
        RECT 255.000 551.700 258.750 552.750 ;
        RECT 296.250 552.600 300.300 554.400 ;
        RECT 302.100 552.600 306.300 554.400 ;
        RECT 308.100 552.600 312.300 554.400 ;
        RECT 296.250 551.700 297.450 552.600 ;
        RECT 302.100 551.700 303.300 552.600 ;
        RECT 308.100 551.700 309.300 552.600 ;
        RECT 313.200 551.700 314.250 554.850 ;
        RECT 155.550 550.800 159.150 551.700 ;
        RECT 113.100 547.950 118.800 549.600 ;
        RECT 71.550 543.750 73.350 546.600 ;
        RECT 74.550 543.750 76.350 546.600 ;
        RECT 77.550 543.750 79.350 546.600 ;
        RECT 113.700 543.750 115.500 546.600 ;
        RECT 117.000 543.750 118.800 547.950 ;
        RECT 121.200 543.750 123.000 549.600 ;
        RECT 152.850 543.750 154.650 549.600 ;
        RECT 157.350 543.750 159.150 550.800 ;
        RECT 194.400 550.500 198.450 551.700 ;
        RECT 200.550 550.500 204.300 551.700 ;
        RECT 206.400 550.500 210.300 551.700 ;
        RECT 212.400 550.650 215.250 551.700 ;
        RECT 212.400 550.500 215.100 550.650 ;
        RECT 194.400 549.600 196.200 550.500 ;
        RECT 191.550 543.750 193.350 549.600 ;
        RECT 194.550 543.750 196.350 549.600 ;
        RECT 197.550 543.750 199.350 549.600 ;
        RECT 200.550 543.750 202.350 550.500 ;
        RECT 206.400 549.600 208.200 550.500 ;
        RECT 212.400 549.600 214.200 550.500 ;
        RECT 203.550 543.750 205.350 549.600 ;
        RECT 206.550 543.750 208.350 549.600 ;
        RECT 209.550 543.750 211.350 549.600 ;
        RECT 212.550 543.750 214.350 549.600 ;
        RECT 215.550 543.750 217.350 549.600 ;
        RECT 248.550 548.700 256.350 550.050 ;
        RECT 248.550 543.750 250.350 548.700 ;
        RECT 251.550 543.750 253.350 547.800 ;
        RECT 254.550 543.750 256.350 548.700 ;
        RECT 257.550 549.600 258.750 551.700 ;
        RECT 293.400 550.500 297.450 551.700 ;
        RECT 299.550 550.500 303.300 551.700 ;
        RECT 305.400 550.500 309.300 551.700 ;
        RECT 311.400 550.650 314.250 551.700 ;
        RECT 350.550 551.700 351.750 559.050 ;
        RECT 352.950 557.850 355.050 559.950 ;
        RECT 383.100 558.150 384.900 559.950 ;
        RECT 353.100 556.050 354.900 557.850 ;
        RECT 382.950 556.050 385.050 558.150 ;
        RECT 387.000 555.150 388.050 562.350 ;
        RECT 389.100 558.150 390.900 559.950 ;
        RECT 388.950 556.050 391.050 558.150 ;
        RECT 425.400 556.950 426.600 569.400 ;
        RECT 461.250 569.100 462.450 569.400 ;
        RECT 466.650 569.400 468.450 575.250 ;
        RECT 469.650 569.400 471.450 575.250 ;
        RECT 500.400 569.400 502.200 575.250 ;
        RECT 466.650 569.100 468.300 569.400 ;
        RECT 461.250 568.200 468.300 569.100 ;
        RECT 461.250 559.950 462.300 568.200 ;
        RECT 467.100 564.150 468.900 565.950 ;
        RECT 463.950 561.150 465.750 562.950 ;
        RECT 466.950 562.050 469.050 564.150 ;
        RECT 503.700 563.400 505.500 575.250 ;
        RECT 507.900 563.400 509.700 575.250 ;
        RECT 541.650 569.400 543.450 575.250 ;
        RECT 544.650 569.400 546.450 575.250 ;
        RECT 547.650 569.400 549.450 575.250 ;
        RECT 470.100 561.150 471.900 562.950 ;
        RECT 500.250 561.150 502.050 562.950 ;
        RECT 460.950 557.850 463.050 559.950 ;
        RECT 463.950 559.050 466.050 561.150 ;
        RECT 469.950 559.050 472.050 561.150 ;
        RECT 499.950 559.050 502.050 561.150 ;
        RECT 503.850 558.150 505.050 563.400 ;
        RECT 545.250 561.150 546.450 569.400 ;
        RECT 580.650 563.400 582.450 575.250 ;
        RECT 583.650 564.300 585.450 575.250 ;
        RECT 586.650 565.200 588.450 575.250 ;
        RECT 589.650 564.300 591.450 575.250 ;
        RECT 583.650 563.400 591.450 564.300 ;
        RECT 621.300 563.400 623.100 575.250 ;
        RECT 625.500 563.400 627.300 575.250 ;
        RECT 628.800 569.400 630.600 575.250 ;
        RECT 662.550 569.400 664.350 575.250 ;
        RECT 665.550 569.400 667.350 575.250 ;
        RECT 668.550 569.400 670.350 575.250 ;
        RECT 703.650 569.400 705.450 575.250 ;
        RECT 706.650 569.400 708.450 575.250 ;
        RECT 509.100 558.150 510.900 559.950 ;
        RECT 422.100 555.150 423.900 556.950 ;
        RECT 385.950 553.050 388.050 555.150 ;
        RECT 421.950 553.050 424.050 555.150 ;
        RECT 424.950 554.850 427.050 556.950 ;
        RECT 350.550 550.800 354.150 551.700 ;
        RECT 311.400 550.500 314.100 550.650 ;
        RECT 293.400 549.600 295.200 550.500 ;
        RECT 257.550 543.750 259.350 549.600 ;
        RECT 290.550 543.750 292.350 549.600 ;
        RECT 293.550 543.750 295.350 549.600 ;
        RECT 296.550 543.750 298.350 549.600 ;
        RECT 299.550 543.750 301.350 550.500 ;
        RECT 305.400 549.600 307.200 550.500 ;
        RECT 311.400 549.600 313.200 550.500 ;
        RECT 302.550 543.750 304.350 549.600 ;
        RECT 305.550 543.750 307.350 549.600 ;
        RECT 308.550 543.750 310.350 549.600 ;
        RECT 311.550 543.750 313.350 549.600 ;
        RECT 314.550 543.750 316.350 549.600 ;
        RECT 347.850 543.750 349.650 549.600 ;
        RECT 352.350 543.750 354.150 550.800 ;
        RECT 387.000 546.600 388.050 553.050 ;
        RECT 425.400 546.600 426.600 554.850 ;
        RECT 461.400 553.650 462.600 557.850 ;
        RECT 502.950 556.050 505.050 558.150 ;
        RECT 461.400 552.000 465.900 553.650 ;
        RECT 502.950 552.750 504.150 556.050 ;
        RECT 505.950 554.850 508.050 556.950 ;
        RECT 508.950 556.050 511.050 558.150 ;
        RECT 541.950 557.850 544.050 559.950 ;
        RECT 544.950 559.050 547.050 561.150 ;
        RECT 542.100 556.050 543.900 557.850 ;
        RECT 506.100 553.050 507.900 554.850 ;
        RECT 383.550 543.750 385.350 546.600 ;
        RECT 386.550 543.750 388.350 546.600 ;
        RECT 389.550 543.750 391.350 546.600 ;
        RECT 422.550 543.750 424.350 546.600 ;
        RECT 425.550 543.750 427.350 546.600 ;
        RECT 464.100 543.750 465.900 552.000 ;
        RECT 469.500 543.750 471.300 552.600 ;
        RECT 500.250 551.700 504.000 552.750 ;
        RECT 545.250 551.700 546.450 559.050 ;
        RECT 547.950 557.850 550.050 559.950 ;
        RECT 581.100 558.150 582.300 563.400 ;
        RECT 620.100 558.150 621.900 559.950 ;
        RECT 625.950 558.150 627.150 563.400 ;
        RECT 628.950 561.150 630.750 562.950 ;
        RECT 665.550 561.150 666.750 569.400 ;
        RECT 628.950 559.050 631.050 561.150 ;
        RECT 548.100 556.050 549.900 557.850 ;
        RECT 580.950 556.050 583.050 558.150 ;
        RECT 500.250 549.600 501.450 551.700 ;
        RECT 542.850 550.800 546.450 551.700 ;
        RECT 499.650 543.750 501.450 549.600 ;
        RECT 502.650 548.700 510.450 550.050 ;
        RECT 502.650 543.750 504.450 548.700 ;
        RECT 505.650 543.750 507.450 547.800 ;
        RECT 508.650 543.750 510.450 548.700 ;
        RECT 542.850 543.750 544.650 550.800 ;
        RECT 581.100 549.600 582.300 556.050 ;
        RECT 583.950 554.850 586.050 556.950 ;
        RECT 587.100 555.150 588.900 556.950 ;
        RECT 584.100 553.050 585.900 554.850 ;
        RECT 586.950 553.050 589.050 555.150 ;
        RECT 589.950 554.850 592.050 556.950 ;
        RECT 619.950 556.050 622.050 558.150 ;
        RECT 622.950 554.850 625.050 556.950 ;
        RECT 625.950 556.050 628.050 558.150 ;
        RECT 661.950 557.850 664.050 559.950 ;
        RECT 664.950 559.050 667.050 561.150 ;
        RECT 662.100 556.050 663.900 557.850 ;
        RECT 590.100 553.050 591.900 554.850 ;
        RECT 623.100 553.050 624.900 554.850 ;
        RECT 626.850 552.750 628.050 556.050 ;
        RECT 627.000 551.700 630.750 552.750 ;
        RECT 547.350 543.750 549.150 549.600 ;
        RECT 581.100 547.950 586.800 549.600 ;
        RECT 581.700 543.750 583.500 546.600 ;
        RECT 585.000 543.750 586.800 547.950 ;
        RECT 589.200 543.750 591.000 549.600 ;
        RECT 620.550 548.700 628.350 550.050 ;
        RECT 620.550 543.750 622.350 548.700 ;
        RECT 623.550 543.750 625.350 547.800 ;
        RECT 626.550 543.750 628.350 548.700 ;
        RECT 629.550 549.600 630.750 551.700 ;
        RECT 665.550 551.700 666.750 559.050 ;
        RECT 667.950 557.850 670.050 559.950 ;
        RECT 668.100 556.050 669.900 557.850 ;
        RECT 704.400 556.950 705.600 569.400 ;
        RECT 737.550 563.400 739.350 575.250 ;
        RECT 741.750 563.400 743.550 575.250 ;
        RECT 741.000 562.350 743.550 563.400 ;
        RECT 737.100 558.150 738.900 559.950 ;
        RECT 703.950 554.850 706.050 556.950 ;
        RECT 707.100 555.150 708.900 556.950 ;
        RECT 736.950 556.050 739.050 558.150 ;
        RECT 741.000 555.150 742.050 562.350 ;
        RECT 743.100 558.150 744.900 559.950 ;
        RECT 742.950 556.050 745.050 558.150 ;
        RECT 665.550 550.800 669.150 551.700 ;
        RECT 629.550 543.750 631.350 549.600 ;
        RECT 662.850 543.750 664.650 549.600 ;
        RECT 667.350 543.750 669.150 550.800 ;
        RECT 704.400 546.600 705.600 554.850 ;
        RECT 706.950 553.050 709.050 555.150 ;
        RECT 739.950 553.050 742.050 555.150 ;
        RECT 741.000 546.600 742.050 553.050 ;
        RECT 703.650 543.750 705.450 546.600 ;
        RECT 706.650 543.750 708.450 546.600 ;
        RECT 737.550 543.750 739.350 546.600 ;
        RECT 740.550 543.750 742.350 546.600 ;
        RECT 743.550 543.750 745.350 546.600 ;
        RECT 30.150 534.900 31.950 539.250 ;
        RECT 28.650 533.400 31.950 534.900 ;
        RECT 33.150 533.400 34.950 539.250 ;
        RECT 28.650 526.950 29.850 533.400 ;
        RECT 31.950 531.900 33.750 532.500 ;
        RECT 37.650 531.900 39.450 539.250 ;
        RECT 31.950 530.700 39.450 531.900 ;
        RECT 28.650 524.850 31.050 526.950 ;
        RECT 32.100 525.150 33.900 526.950 ;
        RECT 28.650 519.600 29.850 524.850 ;
        RECT 31.950 523.050 34.050 525.150 ;
        RECT 28.050 507.750 29.850 519.600 ;
        RECT 31.050 507.750 32.850 519.600 ;
        RECT 35.100 513.600 36.300 530.700 ;
        RECT 65.700 530.400 67.500 539.250 ;
        RECT 71.100 531.000 72.900 539.250 ;
        RECT 107.550 534.300 109.350 539.250 ;
        RECT 110.550 535.200 112.350 539.250 ;
        RECT 113.550 534.300 115.350 539.250 ;
        RECT 107.550 532.950 115.350 534.300 ;
        RECT 116.550 533.400 118.350 539.250 ;
        RECT 151.650 536.400 153.450 539.250 ;
        RECT 154.650 536.400 156.450 539.250 ;
        RECT 157.650 536.400 159.450 539.250 ;
        RECT 188.550 536.400 190.350 539.250 ;
        RECT 116.550 531.300 117.750 533.400 ;
        RECT 71.100 529.350 75.600 531.000 ;
        RECT 114.000 530.250 117.750 531.300 ;
        RECT 37.950 524.850 40.050 526.950 ;
        RECT 74.400 525.150 75.600 529.350 ;
        RECT 110.100 528.150 111.900 529.950 ;
        RECT 38.100 523.050 39.900 524.850 ;
        RECT 64.950 521.850 67.050 523.950 ;
        RECT 70.950 521.850 73.050 523.950 ;
        RECT 73.950 523.050 76.050 525.150 ;
        RECT 106.950 524.850 109.050 526.950 ;
        RECT 109.950 526.050 112.050 528.150 ;
        RECT 113.850 526.950 115.050 530.250 ;
        RECT 154.950 529.950 156.000 536.400 ;
        RECT 189.150 532.500 190.350 536.400 ;
        RECT 191.850 533.400 193.650 539.250 ;
        RECT 194.850 533.400 196.650 539.250 ;
        RECT 227.550 536.400 229.350 539.250 ;
        RECT 189.150 531.600 194.250 532.500 ;
        RECT 192.000 530.700 194.250 531.600 ;
        RECT 154.950 527.850 157.050 529.950 ;
        RECT 112.950 524.850 115.050 526.950 ;
        RECT 151.950 524.850 154.050 526.950 ;
        RECT 107.100 523.050 108.900 524.850 ;
        RECT 65.100 520.050 66.900 521.850 ;
        RECT 67.950 518.850 70.050 520.950 ;
        RECT 71.250 520.050 73.050 521.850 ;
        RECT 68.100 517.050 69.900 518.850 ;
        RECT 74.700 514.800 75.750 523.050 ;
        RECT 112.950 519.600 114.150 524.850 ;
        RECT 115.950 521.850 118.050 523.950 ;
        RECT 152.100 523.050 153.900 524.850 ;
        RECT 115.950 520.050 117.750 521.850 ;
        RECT 154.950 520.650 156.000 527.850 ;
        RECT 157.950 524.850 160.050 526.950 ;
        RECT 187.950 524.850 190.050 526.950 ;
        RECT 158.100 523.050 159.900 524.850 ;
        RECT 188.100 523.050 189.900 524.850 ;
        RECT 192.000 522.300 193.050 530.700 ;
        RECT 195.150 526.950 196.350 533.400 ;
        RECT 228.150 532.500 229.350 536.400 ;
        RECT 230.850 533.400 232.650 539.250 ;
        RECT 233.850 533.400 235.650 539.250 ;
        RECT 268.650 533.400 270.450 539.250 ;
        RECT 228.150 531.600 233.250 532.500 ;
        RECT 231.000 530.700 233.250 531.600 ;
        RECT 193.950 524.850 196.350 526.950 ;
        RECT 226.950 524.850 229.050 526.950 ;
        RECT 192.000 521.400 194.250 522.300 ;
        RECT 153.450 519.600 156.000 520.650 ;
        RECT 188.550 520.500 194.250 521.400 ;
        RECT 68.700 513.900 75.750 514.800 ;
        RECT 68.700 513.600 70.350 513.900 ;
        RECT 34.650 507.750 36.450 513.600 ;
        RECT 37.650 507.750 39.450 513.600 ;
        RECT 65.550 507.750 67.350 513.600 ;
        RECT 68.550 507.750 70.350 513.600 ;
        RECT 74.550 513.600 75.750 513.900 ;
        RECT 71.550 507.750 73.350 513.000 ;
        RECT 74.550 507.750 76.350 513.600 ;
        RECT 108.300 507.750 110.100 519.600 ;
        RECT 112.500 507.750 114.300 519.600 ;
        RECT 115.800 507.750 117.600 513.600 ;
        RECT 153.450 507.750 155.250 519.600 ;
        RECT 157.650 507.750 159.450 519.600 ;
        RECT 188.550 513.600 189.750 520.500 ;
        RECT 195.150 519.600 196.350 524.850 ;
        RECT 227.100 523.050 228.900 524.850 ;
        RECT 231.000 522.300 232.050 530.700 ;
        RECT 234.150 526.950 235.350 533.400 ;
        RECT 269.250 531.300 270.450 533.400 ;
        RECT 271.650 534.300 273.450 539.250 ;
        RECT 274.650 535.200 276.450 539.250 ;
        RECT 277.650 534.300 279.450 539.250 ;
        RECT 310.650 536.400 312.450 539.250 ;
        RECT 313.650 536.400 315.450 539.250 ;
        RECT 344.550 536.400 346.350 539.250 ;
        RECT 347.550 536.400 349.350 539.250 ;
        RECT 350.550 536.400 352.350 539.250 ;
        RECT 271.650 532.950 279.450 534.300 ;
        RECT 269.250 530.250 273.000 531.300 ;
        RECT 232.950 524.850 235.350 526.950 ;
        RECT 271.950 526.950 273.150 530.250 ;
        RECT 275.100 528.150 276.900 529.950 ;
        RECT 311.400 528.150 312.600 536.400 ;
        RECT 348.000 529.950 349.050 536.400 ;
        RECT 381.000 533.400 382.800 539.250 ;
        RECT 385.200 535.050 387.000 539.250 ;
        RECT 388.500 536.400 390.300 539.250 ;
        RECT 385.200 533.400 390.900 535.050 ;
        RECT 426.150 534.900 427.950 539.250 ;
        RECT 271.950 524.850 274.050 526.950 ;
        RECT 274.950 526.050 277.050 528.150 ;
        RECT 277.950 524.850 280.050 526.950 ;
        RECT 310.950 526.050 313.050 528.150 ;
        RECT 313.950 527.850 316.050 529.950 ;
        RECT 346.950 527.850 349.050 529.950 ;
        RECT 380.100 528.150 381.900 529.950 ;
        RECT 314.100 526.050 315.900 527.850 ;
        RECT 231.000 521.400 233.250 522.300 ;
        RECT 227.550 520.500 233.250 521.400 ;
        RECT 188.550 507.750 190.350 513.600 ;
        RECT 191.850 507.750 193.650 519.600 ;
        RECT 194.850 507.750 196.650 519.600 ;
        RECT 227.550 513.600 228.750 520.500 ;
        RECT 234.150 519.600 235.350 524.850 ;
        RECT 268.950 521.850 271.050 523.950 ;
        RECT 269.250 520.050 271.050 521.850 ;
        RECT 272.850 519.600 274.050 524.850 ;
        RECT 278.100 523.050 279.900 524.850 ;
        RECT 227.550 507.750 229.350 513.600 ;
        RECT 230.850 507.750 232.650 519.600 ;
        RECT 233.850 507.750 235.650 519.600 ;
        RECT 269.400 507.750 271.200 513.600 ;
        RECT 272.700 507.750 274.500 519.600 ;
        RECT 276.900 507.750 278.700 519.600 ;
        RECT 311.400 513.600 312.600 526.050 ;
        RECT 343.950 524.850 346.050 526.950 ;
        RECT 344.100 523.050 345.900 524.850 ;
        RECT 348.000 520.650 349.050 527.850 ;
        RECT 349.950 524.850 352.050 526.950 ;
        RECT 379.950 526.050 382.050 528.150 ;
        RECT 382.950 527.850 385.050 529.950 ;
        RECT 386.100 528.150 387.900 529.950 ;
        RECT 383.100 526.050 384.900 527.850 ;
        RECT 385.950 526.050 388.050 528.150 ;
        RECT 389.700 526.950 390.900 533.400 ;
        RECT 424.650 533.400 427.950 534.900 ;
        RECT 429.150 533.400 430.950 539.250 ;
        RECT 424.650 526.950 425.850 533.400 ;
        RECT 427.950 531.900 429.750 532.500 ;
        RECT 433.650 531.900 435.450 539.250 ;
        RECT 464.850 533.400 466.650 539.250 ;
        RECT 469.350 532.200 471.150 539.250 ;
        RECT 502.650 533.400 504.450 539.250 ;
        RECT 427.950 530.700 435.450 531.900 ;
        RECT 467.550 531.300 471.150 532.200 ;
        RECT 503.250 531.300 504.450 533.400 ;
        RECT 505.650 534.300 507.450 539.250 ;
        RECT 508.650 535.200 510.450 539.250 ;
        RECT 511.650 534.300 513.450 539.250 ;
        RECT 505.650 532.950 513.450 534.300 ;
        RECT 515.550 533.400 517.350 539.250 ;
        RECT 518.850 536.400 520.650 539.250 ;
        RECT 523.350 536.400 525.150 539.250 ;
        RECT 527.550 536.400 529.350 539.250 ;
        RECT 531.450 536.400 533.250 539.250 ;
        RECT 534.750 536.400 536.550 539.250 ;
        RECT 539.250 537.300 541.050 539.250 ;
        RECT 539.250 536.400 543.000 537.300 ;
        RECT 544.050 536.400 545.850 539.250 ;
        RECT 523.650 535.500 524.700 536.400 ;
        RECT 520.950 534.300 524.700 535.500 ;
        RECT 532.200 534.600 533.250 536.400 ;
        RECT 541.950 535.500 543.000 536.400 ;
        RECT 520.950 533.400 523.050 534.300 ;
        RECT 388.950 524.850 391.050 526.950 ;
        RECT 424.650 524.850 427.050 526.950 ;
        RECT 428.100 525.150 429.900 526.950 ;
        RECT 350.100 523.050 351.900 524.850 ;
        RECT 348.000 519.600 350.550 520.650 ;
        RECT 389.700 519.600 390.900 524.850 ;
        RECT 424.650 519.600 425.850 524.850 ;
        RECT 427.950 523.050 430.050 525.150 ;
        RECT 310.650 507.750 312.450 513.600 ;
        RECT 313.650 507.750 315.450 513.600 ;
        RECT 344.550 507.750 346.350 519.600 ;
        RECT 348.750 507.750 350.550 519.600 ;
        RECT 380.550 518.700 388.350 519.600 ;
        RECT 380.550 507.750 382.350 518.700 ;
        RECT 383.550 507.750 385.350 517.800 ;
        RECT 386.550 507.750 388.350 518.700 ;
        RECT 389.550 507.750 391.350 519.600 ;
        RECT 424.050 507.750 425.850 519.600 ;
        RECT 427.050 507.750 428.850 519.600 ;
        RECT 431.100 513.600 432.300 530.700 ;
        RECT 433.950 524.850 436.050 526.950 ;
        RECT 464.100 525.150 465.900 526.950 ;
        RECT 434.100 523.050 435.900 524.850 ;
        RECT 463.950 523.050 466.050 525.150 ;
        RECT 467.550 523.950 468.750 531.300 ;
        RECT 503.250 530.250 507.000 531.300 ;
        RECT 515.550 531.150 516.750 533.400 ;
        RECT 528.150 532.200 529.950 534.000 ;
        RECT 532.200 533.550 537.150 534.600 ;
        RECT 535.350 532.800 537.150 533.550 ;
        RECT 538.650 532.800 540.450 534.600 ;
        RECT 541.950 533.400 544.050 535.500 ;
        RECT 547.050 533.400 548.850 539.250 ;
        RECT 529.050 531.900 529.950 532.200 ;
        RECT 539.100 531.900 540.150 532.800 ;
        RECT 505.950 526.950 507.150 530.250 ;
        RECT 509.100 528.150 510.900 529.950 ;
        RECT 515.550 529.050 520.050 531.150 ;
        RECT 529.050 531.000 540.150 531.900 ;
        RECT 470.100 525.150 471.900 526.950 ;
        RECT 466.950 521.850 469.050 523.950 ;
        RECT 469.950 523.050 472.050 525.150 ;
        RECT 505.950 524.850 508.050 526.950 ;
        RECT 508.950 526.050 511.050 528.150 ;
        RECT 511.950 524.850 514.050 526.950 ;
        RECT 502.950 521.850 505.050 523.950 ;
        RECT 467.550 513.600 468.750 521.850 ;
        RECT 503.250 520.050 505.050 521.850 ;
        RECT 506.850 519.600 508.050 524.850 ;
        RECT 512.100 523.050 513.900 524.850 ;
        RECT 515.550 519.600 516.750 529.050 ;
        RECT 517.950 527.250 521.850 529.050 ;
        RECT 517.950 526.950 520.050 527.250 ;
        RECT 529.050 526.950 529.950 531.000 ;
        RECT 539.100 529.800 540.150 531.000 ;
        RECT 539.100 528.600 546.000 529.800 ;
        RECT 539.100 528.000 540.900 528.600 ;
        RECT 545.100 527.850 546.000 528.600 ;
        RECT 542.100 526.950 543.900 527.700 ;
        RECT 529.050 524.850 532.050 526.950 ;
        RECT 535.950 525.900 543.900 526.950 ;
        RECT 545.100 526.050 546.900 527.850 ;
        RECT 535.950 524.850 538.050 525.900 ;
        RECT 517.950 521.400 519.750 523.200 ;
        RECT 518.850 520.200 523.050 521.400 ;
        RECT 529.050 520.200 529.950 524.850 ;
        RECT 537.750 521.100 539.550 521.400 ;
        RECT 430.650 507.750 432.450 513.600 ;
        RECT 433.650 507.750 435.450 513.600 ;
        RECT 464.550 507.750 466.350 513.600 ;
        RECT 467.550 507.750 469.350 513.600 ;
        RECT 470.550 507.750 472.350 513.600 ;
        RECT 503.400 507.750 505.200 513.600 ;
        RECT 506.700 507.750 508.500 519.600 ;
        RECT 510.900 507.750 512.700 519.600 ;
        RECT 515.550 507.750 517.350 519.600 ;
        RECT 520.950 519.300 523.050 520.200 ;
        RECT 523.950 519.300 529.950 520.200 ;
        RECT 531.150 520.800 539.550 521.100 ;
        RECT 547.950 520.800 548.850 533.400 ;
        RECT 581.850 532.200 583.650 539.250 ;
        RECT 586.350 533.400 588.150 539.250 ;
        RECT 590.550 533.400 592.350 539.250 ;
        RECT 593.850 536.400 595.650 539.250 ;
        RECT 598.350 536.400 600.150 539.250 ;
        RECT 602.550 536.400 604.350 539.250 ;
        RECT 606.450 536.400 608.250 539.250 ;
        RECT 609.750 536.400 611.550 539.250 ;
        RECT 614.250 537.300 616.050 539.250 ;
        RECT 614.250 536.400 618.000 537.300 ;
        RECT 619.050 536.400 620.850 539.250 ;
        RECT 598.650 535.500 599.700 536.400 ;
        RECT 595.950 534.300 599.700 535.500 ;
        RECT 607.200 534.600 608.250 536.400 ;
        RECT 616.950 535.500 618.000 536.400 ;
        RECT 595.950 533.400 598.050 534.300 ;
        RECT 581.850 531.300 585.450 532.200 ;
        RECT 581.100 525.150 582.900 526.950 ;
        RECT 580.950 523.050 583.050 525.150 ;
        RECT 584.250 523.950 585.450 531.300 ;
        RECT 590.550 531.150 591.750 533.400 ;
        RECT 603.150 532.200 604.950 534.000 ;
        RECT 607.200 533.550 612.150 534.600 ;
        RECT 610.350 532.800 612.150 533.550 ;
        RECT 613.650 532.800 615.450 534.600 ;
        RECT 616.950 533.400 619.050 535.500 ;
        RECT 622.050 533.400 623.850 539.250 ;
        RECT 653.850 533.400 655.650 539.250 ;
        RECT 604.050 531.900 604.950 532.200 ;
        RECT 614.100 531.900 615.150 532.800 ;
        RECT 590.550 529.050 595.050 531.150 ;
        RECT 604.050 531.000 615.150 531.900 ;
        RECT 587.100 525.150 588.900 526.950 ;
        RECT 583.950 521.850 586.050 523.950 ;
        RECT 586.950 523.050 589.050 525.150 ;
        RECT 531.150 520.200 548.850 520.800 ;
        RECT 523.950 518.400 524.850 519.300 ;
        RECT 522.150 516.600 524.850 518.400 ;
        RECT 525.750 518.100 527.550 518.400 ;
        RECT 531.150 518.100 532.050 520.200 ;
        RECT 537.750 519.600 548.850 520.200 ;
        RECT 525.750 517.200 532.050 518.100 ;
        RECT 532.950 518.700 534.750 519.300 ;
        RECT 532.950 517.500 540.450 518.700 ;
        RECT 525.750 516.600 527.550 517.200 ;
        RECT 539.250 516.600 540.450 517.500 ;
        RECT 520.950 513.600 524.850 515.700 ;
        RECT 529.950 514.500 536.850 516.300 ;
        RECT 539.250 514.500 544.050 516.600 ;
        RECT 518.550 507.750 520.350 510.600 ;
        RECT 523.050 507.750 524.850 513.600 ;
        RECT 527.250 507.750 529.050 513.600 ;
        RECT 531.150 507.750 532.950 514.500 ;
        RECT 539.250 513.600 540.450 514.500 ;
        RECT 534.150 507.750 535.950 513.600 ;
        RECT 538.950 507.750 540.750 513.600 ;
        RECT 544.050 507.750 545.850 513.600 ;
        RECT 547.050 507.750 548.850 519.600 ;
        RECT 584.250 513.600 585.450 521.850 ;
        RECT 590.550 519.600 591.750 529.050 ;
        RECT 592.950 527.250 596.850 529.050 ;
        RECT 592.950 526.950 595.050 527.250 ;
        RECT 604.050 526.950 604.950 531.000 ;
        RECT 614.100 529.800 615.150 531.000 ;
        RECT 614.100 528.600 621.000 529.800 ;
        RECT 614.100 528.000 615.900 528.600 ;
        RECT 620.100 527.850 621.000 528.600 ;
        RECT 617.100 526.950 618.900 527.700 ;
        RECT 604.050 524.850 607.050 526.950 ;
        RECT 610.950 525.900 618.900 526.950 ;
        RECT 620.100 526.050 621.900 527.850 ;
        RECT 610.950 524.850 613.050 525.900 ;
        RECT 592.950 521.400 594.750 523.200 ;
        RECT 593.850 520.200 598.050 521.400 ;
        RECT 604.050 520.200 604.950 524.850 ;
        RECT 612.750 521.100 614.550 521.400 ;
        RECT 580.650 507.750 582.450 513.600 ;
        RECT 583.650 507.750 585.450 513.600 ;
        RECT 586.650 507.750 588.450 513.600 ;
        RECT 590.550 507.750 592.350 519.600 ;
        RECT 595.950 519.300 598.050 520.200 ;
        RECT 598.950 519.300 604.950 520.200 ;
        RECT 606.150 520.800 614.550 521.100 ;
        RECT 622.950 520.800 623.850 533.400 ;
        RECT 658.350 532.200 660.150 539.250 ;
        RECT 692.550 536.400 694.350 539.250 ;
        RECT 695.550 536.400 697.350 539.250 ;
        RECT 730.650 536.400 732.450 539.250 ;
        RECT 733.650 536.400 735.450 539.250 ;
        RECT 652.950 531.450 655.050 532.050 ;
        RECT 606.150 520.200 623.850 520.800 ;
        RECT 598.950 518.400 599.850 519.300 ;
        RECT 597.150 516.600 599.850 518.400 ;
        RECT 600.750 518.100 602.550 518.400 ;
        RECT 606.150 518.100 607.050 520.200 ;
        RECT 612.750 519.600 623.850 520.200 ;
        RECT 650.550 530.550 655.050 531.450 ;
        RECT 650.550 520.050 651.450 530.550 ;
        RECT 652.950 529.950 655.050 530.550 ;
        RECT 656.550 531.300 660.150 532.200 ;
        RECT 653.100 525.150 654.900 526.950 ;
        RECT 652.950 523.050 655.050 525.150 ;
        RECT 656.550 523.950 657.750 531.300 ;
        RECT 691.950 527.850 694.050 529.950 ;
        RECT 695.400 528.150 696.600 536.400 ;
        RECT 731.400 528.150 732.600 536.400 ;
        RECT 659.100 525.150 660.900 526.950 ;
        RECT 692.100 526.050 693.900 527.850 ;
        RECT 694.950 526.050 697.050 528.150 ;
        RECT 730.950 526.050 733.050 528.150 ;
        RECT 733.950 527.850 736.050 529.950 ;
        RECT 734.100 526.050 735.900 527.850 ;
        RECT 655.950 521.850 658.050 523.950 ;
        RECT 658.950 523.050 661.050 525.150 ;
        RECT 600.750 517.200 607.050 518.100 ;
        RECT 607.950 518.700 609.750 519.300 ;
        RECT 607.950 517.500 615.450 518.700 ;
        RECT 600.750 516.600 602.550 517.200 ;
        RECT 614.250 516.600 615.450 517.500 ;
        RECT 595.950 513.600 599.850 515.700 ;
        RECT 604.950 514.500 611.850 516.300 ;
        RECT 614.250 514.500 619.050 516.600 ;
        RECT 593.550 507.750 595.350 510.600 ;
        RECT 598.050 507.750 599.850 513.600 ;
        RECT 602.250 507.750 604.050 513.600 ;
        RECT 606.150 507.750 607.950 514.500 ;
        RECT 614.250 513.600 615.450 514.500 ;
        RECT 609.150 507.750 610.950 513.600 ;
        RECT 613.950 507.750 615.750 513.600 ;
        RECT 619.050 507.750 620.850 513.600 ;
        RECT 622.050 507.750 623.850 519.600 ;
        RECT 649.950 517.950 652.050 520.050 ;
        RECT 656.550 513.600 657.750 521.850 ;
        RECT 695.400 513.600 696.600 526.050 ;
        RECT 731.400 513.600 732.600 526.050 ;
        RECT 653.550 507.750 655.350 513.600 ;
        RECT 656.550 507.750 658.350 513.600 ;
        RECT 659.550 507.750 661.350 513.600 ;
        RECT 692.550 507.750 694.350 513.600 ;
        RECT 695.550 507.750 697.350 513.600 ;
        RECT 730.650 507.750 732.450 513.600 ;
        RECT 733.650 507.750 735.450 513.600 ;
        RECT 29.550 497.400 31.350 503.250 ;
        RECT 32.550 497.400 34.350 503.250 ;
        RECT 29.100 486.150 30.900 487.950 ;
        RECT 28.950 484.050 31.050 486.150 ;
        RECT 32.700 480.300 33.900 497.400 ;
        RECT 36.150 491.400 37.950 503.250 ;
        RECT 39.150 491.400 40.950 503.250 ;
        RECT 71.550 491.400 73.350 503.250 ;
        RECT 75.750 491.400 77.550 503.250 ;
        RECT 110.400 497.400 112.200 503.250 ;
        RECT 113.700 491.400 115.500 503.250 ;
        RECT 117.900 491.400 119.700 503.250 ;
        RECT 153.450 491.400 155.250 503.250 ;
        RECT 157.650 491.400 159.450 503.250 ;
        RECT 188.550 497.400 190.350 503.250 ;
        RECT 34.950 485.850 37.050 487.950 ;
        RECT 39.150 486.150 40.350 491.400 ;
        RECT 75.000 490.350 77.550 491.400 ;
        RECT 71.100 486.150 72.900 487.950 ;
        RECT 35.100 484.050 36.900 485.850 ;
        RECT 37.950 484.050 40.350 486.150 ;
        RECT 70.950 484.050 73.050 486.150 ;
        RECT 29.550 479.100 37.050 480.300 ;
        RECT 29.550 471.750 31.350 479.100 ;
        RECT 35.250 478.500 37.050 479.100 ;
        RECT 39.150 477.600 40.350 484.050 ;
        RECT 75.000 483.150 76.050 490.350 ;
        RECT 110.250 489.150 112.050 490.950 ;
        RECT 77.100 486.150 78.900 487.950 ;
        RECT 109.950 487.050 112.050 489.150 ;
        RECT 113.850 486.150 115.050 491.400 ;
        RECT 153.450 490.350 156.000 491.400 ;
        RECT 119.100 486.150 120.900 487.950 ;
        RECT 152.100 486.150 153.900 487.950 ;
        RECT 76.950 484.050 79.050 486.150 ;
        RECT 112.950 484.050 115.050 486.150 ;
        RECT 73.950 481.050 76.050 483.150 ;
        RECT 34.050 471.750 35.850 477.600 ;
        RECT 37.050 476.100 40.350 477.600 ;
        RECT 37.050 471.750 38.850 476.100 ;
        RECT 75.000 474.600 76.050 481.050 ;
        RECT 112.950 480.750 114.150 484.050 ;
        RECT 115.950 482.850 118.050 484.950 ;
        RECT 118.950 484.050 121.050 486.150 ;
        RECT 151.950 484.050 154.050 486.150 ;
        RECT 154.950 483.150 156.000 490.350 ;
        RECT 188.550 490.500 189.750 497.400 ;
        RECT 191.850 491.400 193.650 503.250 ;
        RECT 194.850 491.400 196.650 503.250 ;
        RECT 201.150 491.400 202.950 503.250 ;
        RECT 204.150 497.400 205.950 503.250 ;
        RECT 209.250 497.400 211.050 503.250 ;
        RECT 214.050 497.400 215.850 503.250 ;
        RECT 209.550 496.500 210.750 497.400 ;
        RECT 217.050 496.500 218.850 503.250 ;
        RECT 220.950 497.400 222.750 503.250 ;
        RECT 225.150 497.400 226.950 503.250 ;
        RECT 229.650 500.400 231.450 503.250 ;
        RECT 205.950 494.400 210.750 496.500 ;
        RECT 213.150 494.700 220.050 496.500 ;
        RECT 225.150 495.300 229.050 497.400 ;
        RECT 209.550 493.500 210.750 494.400 ;
        RECT 222.450 493.800 224.250 494.400 ;
        RECT 209.550 492.300 217.050 493.500 ;
        RECT 215.250 491.700 217.050 492.300 ;
        RECT 217.950 492.900 224.250 493.800 ;
        RECT 188.550 489.600 194.250 490.500 ;
        RECT 192.000 488.700 194.250 489.600 ;
        RECT 158.100 486.150 159.900 487.950 ;
        RECT 188.100 486.150 189.900 487.950 ;
        RECT 157.950 484.050 160.050 486.150 ;
        RECT 187.950 484.050 190.050 486.150 ;
        RECT 116.100 481.050 117.900 482.850 ;
        RECT 154.950 481.050 157.050 483.150 ;
        RECT 110.250 479.700 114.000 480.750 ;
        RECT 110.250 477.600 111.450 479.700 ;
        RECT 71.550 471.750 73.350 474.600 ;
        RECT 74.550 471.750 76.350 474.600 ;
        RECT 77.550 471.750 79.350 474.600 ;
        RECT 109.650 471.750 111.450 477.600 ;
        RECT 112.650 476.700 120.450 478.050 ;
        RECT 112.650 471.750 114.450 476.700 ;
        RECT 115.650 471.750 117.450 475.800 ;
        RECT 118.650 471.750 120.450 476.700 ;
        RECT 154.950 474.600 156.000 481.050 ;
        RECT 192.000 480.300 193.050 488.700 ;
        RECT 195.150 486.150 196.350 491.400 ;
        RECT 193.950 484.050 196.350 486.150 ;
        RECT 192.000 479.400 194.250 480.300 ;
        RECT 189.150 478.500 194.250 479.400 ;
        RECT 189.150 474.600 190.350 478.500 ;
        RECT 195.150 477.600 196.350 484.050 ;
        RECT 201.150 490.800 212.250 491.400 ;
        RECT 217.950 490.800 218.850 492.900 ;
        RECT 222.450 492.600 224.250 492.900 ;
        RECT 225.150 492.600 227.850 494.400 ;
        RECT 225.150 491.700 226.050 492.600 ;
        RECT 201.150 490.200 218.850 490.800 ;
        RECT 201.150 477.600 202.050 490.200 ;
        RECT 210.450 489.900 218.850 490.200 ;
        RECT 220.050 490.800 226.050 491.700 ;
        RECT 226.950 490.800 229.050 491.700 ;
        RECT 232.650 491.400 234.450 503.250 ;
        RECT 265.650 491.400 267.450 503.250 ;
        RECT 268.650 492.300 270.450 503.250 ;
        RECT 271.650 493.200 273.450 503.250 ;
        RECT 274.650 492.300 276.450 503.250 ;
        RECT 305.550 497.400 307.350 503.250 ;
        RECT 308.550 497.400 310.350 503.250 ;
        RECT 311.550 497.400 313.350 503.250 ;
        RECT 268.650 491.400 276.450 492.300 ;
        RECT 210.450 489.600 212.250 489.900 ;
        RECT 220.050 486.150 220.950 490.800 ;
        RECT 226.950 489.600 231.150 490.800 ;
        RECT 230.250 487.800 232.050 489.600 ;
        RECT 211.950 485.100 214.050 486.150 ;
        RECT 203.100 483.150 204.900 484.950 ;
        RECT 206.100 484.050 214.050 485.100 ;
        RECT 217.950 484.050 220.950 486.150 ;
        RECT 206.100 483.300 207.900 484.050 ;
        RECT 204.000 482.400 204.900 483.150 ;
        RECT 209.100 482.400 210.900 483.000 ;
        RECT 204.000 481.200 210.900 482.400 ;
        RECT 209.850 480.000 210.900 481.200 ;
        RECT 220.050 480.000 220.950 484.050 ;
        RECT 229.950 483.750 232.050 484.050 ;
        RECT 228.150 481.950 232.050 483.750 ;
        RECT 233.250 481.950 234.450 491.400 ;
        RECT 266.100 486.150 267.300 491.400 ;
        RECT 308.550 489.150 309.750 497.400 ;
        RECT 317.550 491.400 319.350 503.250 ;
        RECT 320.550 500.400 322.350 503.250 ;
        RECT 325.050 497.400 326.850 503.250 ;
        RECT 329.250 497.400 331.050 503.250 ;
        RECT 322.950 495.300 326.850 497.400 ;
        RECT 333.150 496.500 334.950 503.250 ;
        RECT 336.150 497.400 337.950 503.250 ;
        RECT 340.950 497.400 342.750 503.250 ;
        RECT 346.050 497.400 347.850 503.250 ;
        RECT 341.250 496.500 342.450 497.400 ;
        RECT 331.950 494.700 338.850 496.500 ;
        RECT 341.250 494.400 346.050 496.500 ;
        RECT 324.150 492.600 326.850 494.400 ;
        RECT 327.750 493.800 329.550 494.400 ;
        RECT 327.750 492.900 334.050 493.800 ;
        RECT 341.250 493.500 342.450 494.400 ;
        RECT 327.750 492.600 329.550 492.900 ;
        RECT 325.950 491.700 326.850 492.600 ;
        RECT 265.950 484.050 268.050 486.150 ;
        RECT 304.950 485.850 307.050 487.950 ;
        RECT 307.950 487.050 310.050 489.150 ;
        RECT 209.850 479.100 220.950 480.000 ;
        RECT 229.950 479.850 234.450 481.950 ;
        RECT 209.850 478.200 210.900 479.100 ;
        RECT 220.050 478.800 220.950 479.100 ;
        RECT 151.650 471.750 153.450 474.600 ;
        RECT 154.650 471.750 156.450 474.600 ;
        RECT 157.650 471.750 159.450 474.600 ;
        RECT 188.550 471.750 190.350 474.600 ;
        RECT 191.850 471.750 193.650 477.600 ;
        RECT 194.850 471.750 196.650 477.600 ;
        RECT 201.150 471.750 202.950 477.600 ;
        RECT 205.950 475.500 208.050 477.600 ;
        RECT 209.550 476.400 211.350 478.200 ;
        RECT 212.850 477.450 214.650 478.200 ;
        RECT 212.850 476.400 217.800 477.450 ;
        RECT 220.050 477.000 221.850 478.800 ;
        RECT 233.250 477.600 234.450 479.850 ;
        RECT 226.950 476.700 229.050 477.600 ;
        RECT 207.000 474.600 208.050 475.500 ;
        RECT 216.750 474.600 217.800 476.400 ;
        RECT 225.300 475.500 229.050 476.700 ;
        RECT 225.300 474.600 226.350 475.500 ;
        RECT 204.150 471.750 205.950 474.600 ;
        RECT 207.000 473.700 210.750 474.600 ;
        RECT 208.950 471.750 210.750 473.700 ;
        RECT 213.450 471.750 215.250 474.600 ;
        RECT 216.750 471.750 218.550 474.600 ;
        RECT 220.650 471.750 222.450 474.600 ;
        RECT 224.850 471.750 226.650 474.600 ;
        RECT 229.350 471.750 231.150 474.600 ;
        RECT 232.650 471.750 234.450 477.600 ;
        RECT 266.100 477.600 267.300 484.050 ;
        RECT 268.950 482.850 271.050 484.950 ;
        RECT 272.100 483.150 273.900 484.950 ;
        RECT 269.100 481.050 270.900 482.850 ;
        RECT 271.950 481.050 274.050 483.150 ;
        RECT 274.950 482.850 277.050 484.950 ;
        RECT 305.100 484.050 306.900 485.850 ;
        RECT 275.100 481.050 276.900 482.850 ;
        RECT 308.550 479.700 309.750 487.050 ;
        RECT 310.950 485.850 313.050 487.950 ;
        RECT 311.100 484.050 312.900 485.850 ;
        RECT 317.550 481.950 318.750 491.400 ;
        RECT 322.950 490.800 325.050 491.700 ;
        RECT 325.950 490.800 331.950 491.700 ;
        RECT 320.850 489.600 325.050 490.800 ;
        RECT 319.950 487.800 321.750 489.600 ;
        RECT 331.050 486.150 331.950 490.800 ;
        RECT 333.150 490.800 334.050 492.900 ;
        RECT 334.950 492.300 342.450 493.500 ;
        RECT 334.950 491.700 336.750 492.300 ;
        RECT 349.050 491.400 350.850 503.250 ;
        RECT 380.550 491.400 382.350 503.250 ;
        RECT 384.750 491.400 386.550 503.250 ;
        RECT 422.400 497.400 424.200 503.250 ;
        RECT 425.700 491.400 427.500 503.250 ;
        RECT 429.900 491.400 431.700 503.250 ;
        RECT 461.550 497.400 463.350 503.250 ;
        RECT 464.550 497.400 466.350 503.250 ;
        RECT 339.750 490.800 350.850 491.400 ;
        RECT 333.150 490.200 350.850 490.800 ;
        RECT 333.150 489.900 341.550 490.200 ;
        RECT 339.750 489.600 341.550 489.900 ;
        RECT 331.050 484.050 334.050 486.150 ;
        RECT 337.950 485.100 340.050 486.150 ;
        RECT 337.950 484.050 345.900 485.100 ;
        RECT 319.950 483.750 322.050 484.050 ;
        RECT 319.950 481.950 323.850 483.750 ;
        RECT 317.550 479.850 322.050 481.950 ;
        RECT 331.050 480.000 331.950 484.050 ;
        RECT 344.100 483.300 345.900 484.050 ;
        RECT 347.100 483.150 348.900 484.950 ;
        RECT 341.100 482.400 342.900 483.000 ;
        RECT 347.100 482.400 348.000 483.150 ;
        RECT 341.100 481.200 348.000 482.400 ;
        RECT 341.100 480.000 342.150 481.200 ;
        RECT 308.550 478.800 312.150 479.700 ;
        RECT 266.100 475.950 271.800 477.600 ;
        RECT 266.700 471.750 268.500 474.600 ;
        RECT 270.000 471.750 271.800 475.950 ;
        RECT 274.200 471.750 276.000 477.600 ;
        RECT 305.850 471.750 307.650 477.600 ;
        RECT 310.350 471.750 312.150 478.800 ;
        RECT 317.550 477.600 318.750 479.850 ;
        RECT 331.050 479.100 342.150 480.000 ;
        RECT 331.050 478.800 331.950 479.100 ;
        RECT 317.550 471.750 319.350 477.600 ;
        RECT 322.950 476.700 325.050 477.600 ;
        RECT 330.150 477.000 331.950 478.800 ;
        RECT 341.100 478.200 342.150 479.100 ;
        RECT 337.350 477.450 339.150 478.200 ;
        RECT 322.950 475.500 326.700 476.700 ;
        RECT 325.650 474.600 326.700 475.500 ;
        RECT 334.200 476.400 339.150 477.450 ;
        RECT 340.650 476.400 342.450 478.200 ;
        RECT 349.950 477.600 350.850 490.200 ;
        RECT 384.000 490.350 386.550 491.400 ;
        RECT 380.100 486.150 381.900 487.950 ;
        RECT 379.950 484.050 382.050 486.150 ;
        RECT 384.000 483.150 385.050 490.350 ;
        RECT 422.250 489.150 424.050 490.950 ;
        RECT 386.100 486.150 387.900 487.950 ;
        RECT 421.950 487.050 424.050 489.150 ;
        RECT 425.850 486.150 427.050 491.400 ;
        RECT 431.100 486.150 432.900 487.950 ;
        RECT 385.950 484.050 388.050 486.150 ;
        RECT 424.950 484.050 427.050 486.150 ;
        RECT 382.950 481.050 385.050 483.150 ;
        RECT 334.200 474.600 335.250 476.400 ;
        RECT 343.950 475.500 346.050 477.600 ;
        RECT 343.950 474.600 345.000 475.500 ;
        RECT 320.850 471.750 322.650 474.600 ;
        RECT 325.350 471.750 327.150 474.600 ;
        RECT 329.550 471.750 331.350 474.600 ;
        RECT 333.450 471.750 335.250 474.600 ;
        RECT 336.750 471.750 338.550 474.600 ;
        RECT 341.250 473.700 345.000 474.600 ;
        RECT 341.250 471.750 343.050 473.700 ;
        RECT 346.050 471.750 347.850 474.600 ;
        RECT 349.050 471.750 350.850 477.600 ;
        RECT 384.000 474.600 385.050 481.050 ;
        RECT 424.950 480.750 426.150 484.050 ;
        RECT 427.950 482.850 430.050 484.950 ;
        RECT 430.950 484.050 433.050 486.150 ;
        RECT 464.400 484.950 465.600 497.400 ;
        RECT 497.550 492.300 499.350 503.250 ;
        RECT 500.550 493.200 502.350 503.250 ;
        RECT 503.550 492.300 505.350 503.250 ;
        RECT 497.550 491.400 505.350 492.300 ;
        RECT 506.550 491.400 508.350 503.250 ;
        RECT 512.550 491.400 514.350 503.250 ;
        RECT 515.550 500.400 517.350 503.250 ;
        RECT 520.050 497.400 521.850 503.250 ;
        RECT 524.250 497.400 526.050 503.250 ;
        RECT 517.950 495.300 521.850 497.400 ;
        RECT 528.150 496.500 529.950 503.250 ;
        RECT 531.150 497.400 532.950 503.250 ;
        RECT 535.950 497.400 537.750 503.250 ;
        RECT 541.050 497.400 542.850 503.250 ;
        RECT 536.250 496.500 537.450 497.400 ;
        RECT 526.950 494.700 533.850 496.500 ;
        RECT 536.250 494.400 541.050 496.500 ;
        RECT 519.150 492.600 521.850 494.400 ;
        RECT 522.750 493.800 524.550 494.400 ;
        RECT 522.750 492.900 529.050 493.800 ;
        RECT 536.250 493.500 537.450 494.400 ;
        RECT 522.750 492.600 524.550 492.900 ;
        RECT 520.950 491.700 521.850 492.600 ;
        RECT 506.700 486.150 507.900 491.400 ;
        RECT 461.100 483.150 462.900 484.950 ;
        RECT 428.100 481.050 429.900 482.850 ;
        RECT 460.950 481.050 463.050 483.150 ;
        RECT 463.950 482.850 466.050 484.950 ;
        RECT 496.950 482.850 499.050 484.950 ;
        RECT 500.100 483.150 501.900 484.950 ;
        RECT 422.250 479.700 426.000 480.750 ;
        RECT 422.250 477.600 423.450 479.700 ;
        RECT 380.550 471.750 382.350 474.600 ;
        RECT 383.550 471.750 385.350 474.600 ;
        RECT 386.550 471.750 388.350 474.600 ;
        RECT 421.650 471.750 423.450 477.600 ;
        RECT 424.650 476.700 432.450 478.050 ;
        RECT 424.650 471.750 426.450 476.700 ;
        RECT 427.650 471.750 429.450 475.800 ;
        RECT 430.650 471.750 432.450 476.700 ;
        RECT 464.400 474.600 465.600 482.850 ;
        RECT 497.100 481.050 498.900 482.850 ;
        RECT 499.950 481.050 502.050 483.150 ;
        RECT 502.950 482.850 505.050 484.950 ;
        RECT 505.950 484.050 508.050 486.150 ;
        RECT 503.100 481.050 504.900 482.850 ;
        RECT 506.700 477.600 507.900 484.050 ;
        RECT 461.550 471.750 463.350 474.600 ;
        RECT 464.550 471.750 466.350 474.600 ;
        RECT 498.000 471.750 499.800 477.600 ;
        RECT 502.200 475.950 507.900 477.600 ;
        RECT 512.550 481.950 513.750 491.400 ;
        RECT 517.950 490.800 520.050 491.700 ;
        RECT 520.950 490.800 526.950 491.700 ;
        RECT 515.850 489.600 520.050 490.800 ;
        RECT 514.950 487.800 516.750 489.600 ;
        RECT 526.050 486.150 526.950 490.800 ;
        RECT 528.150 490.800 529.050 492.900 ;
        RECT 529.950 492.300 537.450 493.500 ;
        RECT 529.950 491.700 531.750 492.300 ;
        RECT 544.050 491.400 545.850 503.250 ;
        RECT 575.550 492.300 577.350 503.250 ;
        RECT 578.550 493.200 580.350 503.250 ;
        RECT 581.550 492.300 583.350 503.250 ;
        RECT 575.550 491.400 583.350 492.300 ;
        RECT 584.550 491.400 586.350 503.250 ;
        RECT 590.550 491.400 592.350 503.250 ;
        RECT 593.550 500.400 595.350 503.250 ;
        RECT 598.050 497.400 599.850 503.250 ;
        RECT 602.250 497.400 604.050 503.250 ;
        RECT 595.950 495.300 599.850 497.400 ;
        RECT 606.150 496.500 607.950 503.250 ;
        RECT 609.150 497.400 610.950 503.250 ;
        RECT 613.950 497.400 615.750 503.250 ;
        RECT 619.050 497.400 620.850 503.250 ;
        RECT 614.250 496.500 615.450 497.400 ;
        RECT 604.950 494.700 611.850 496.500 ;
        RECT 614.250 494.400 619.050 496.500 ;
        RECT 597.150 492.600 599.850 494.400 ;
        RECT 600.750 493.800 602.550 494.400 ;
        RECT 600.750 492.900 607.050 493.800 ;
        RECT 614.250 493.500 615.450 494.400 ;
        RECT 600.750 492.600 602.550 492.900 ;
        RECT 598.950 491.700 599.850 492.600 ;
        RECT 534.750 490.800 545.850 491.400 ;
        RECT 528.150 490.200 545.850 490.800 ;
        RECT 528.150 489.900 536.550 490.200 ;
        RECT 534.750 489.600 536.550 489.900 ;
        RECT 526.050 484.050 529.050 486.150 ;
        RECT 532.950 485.100 535.050 486.150 ;
        RECT 532.950 484.050 540.900 485.100 ;
        RECT 514.950 483.750 517.050 484.050 ;
        RECT 514.950 481.950 518.850 483.750 ;
        RECT 512.550 479.850 517.050 481.950 ;
        RECT 526.050 480.000 526.950 484.050 ;
        RECT 539.100 483.300 540.900 484.050 ;
        RECT 542.100 483.150 543.900 484.950 ;
        RECT 536.100 482.400 537.900 483.000 ;
        RECT 542.100 482.400 543.000 483.150 ;
        RECT 536.100 481.200 543.000 482.400 ;
        RECT 536.100 480.000 537.150 481.200 ;
        RECT 512.550 477.600 513.750 479.850 ;
        RECT 526.050 479.100 537.150 480.000 ;
        RECT 526.050 478.800 526.950 479.100 ;
        RECT 502.200 471.750 504.000 475.950 ;
        RECT 505.500 471.750 507.300 474.600 ;
        RECT 512.550 471.750 514.350 477.600 ;
        RECT 517.950 476.700 520.050 477.600 ;
        RECT 525.150 477.000 526.950 478.800 ;
        RECT 536.100 478.200 537.150 479.100 ;
        RECT 532.350 477.450 534.150 478.200 ;
        RECT 517.950 475.500 521.700 476.700 ;
        RECT 520.650 474.600 521.700 475.500 ;
        RECT 529.200 476.400 534.150 477.450 ;
        RECT 535.650 476.400 537.450 478.200 ;
        RECT 544.950 477.600 545.850 490.200 ;
        RECT 584.700 486.150 585.900 491.400 ;
        RECT 574.950 482.850 577.050 484.950 ;
        RECT 578.100 483.150 579.900 484.950 ;
        RECT 575.100 481.050 576.900 482.850 ;
        RECT 577.950 481.050 580.050 483.150 ;
        RECT 580.950 482.850 583.050 484.950 ;
        RECT 583.950 484.050 586.050 486.150 ;
        RECT 581.100 481.050 582.900 482.850 ;
        RECT 584.700 477.600 585.900 484.050 ;
        RECT 529.200 474.600 530.250 476.400 ;
        RECT 538.950 475.500 541.050 477.600 ;
        RECT 538.950 474.600 540.000 475.500 ;
        RECT 515.850 471.750 517.650 474.600 ;
        RECT 520.350 471.750 522.150 474.600 ;
        RECT 524.550 471.750 526.350 474.600 ;
        RECT 528.450 471.750 530.250 474.600 ;
        RECT 531.750 471.750 533.550 474.600 ;
        RECT 536.250 473.700 540.000 474.600 ;
        RECT 536.250 471.750 538.050 473.700 ;
        RECT 541.050 471.750 542.850 474.600 ;
        RECT 544.050 471.750 545.850 477.600 ;
        RECT 576.000 471.750 577.800 477.600 ;
        RECT 580.200 475.950 585.900 477.600 ;
        RECT 590.550 481.950 591.750 491.400 ;
        RECT 595.950 490.800 598.050 491.700 ;
        RECT 598.950 490.800 604.950 491.700 ;
        RECT 593.850 489.600 598.050 490.800 ;
        RECT 592.950 487.800 594.750 489.600 ;
        RECT 604.050 486.150 604.950 490.800 ;
        RECT 606.150 490.800 607.050 492.900 ;
        RECT 607.950 492.300 615.450 493.500 ;
        RECT 607.950 491.700 609.750 492.300 ;
        RECT 622.050 491.400 623.850 503.250 ;
        RECT 653.550 492.600 655.350 503.250 ;
        RECT 656.550 493.500 658.350 503.250 ;
        RECT 659.550 502.500 667.350 503.250 ;
        RECT 659.550 492.600 661.350 502.500 ;
        RECT 653.550 491.700 661.350 492.600 ;
        RECT 662.550 491.400 664.350 501.600 ;
        RECT 665.550 491.400 667.350 502.500 ;
        RECT 698.550 492.300 700.350 503.250 ;
        RECT 701.550 493.200 703.350 503.250 ;
        RECT 704.550 492.300 706.350 503.250 ;
        RECT 698.550 491.400 706.350 492.300 ;
        RECT 707.550 491.400 709.350 503.250 ;
        RECT 741.300 491.400 743.100 503.250 ;
        RECT 745.500 491.400 747.300 503.250 ;
        RECT 748.800 497.400 750.600 503.250 ;
        RECT 612.750 490.800 623.850 491.400 ;
        RECT 606.150 490.200 623.850 490.800 ;
        RECT 662.400 490.500 664.200 491.400 ;
        RECT 606.150 489.900 614.550 490.200 ;
        RECT 612.750 489.600 614.550 489.900 ;
        RECT 604.050 484.050 607.050 486.150 ;
        RECT 610.950 485.100 613.050 486.150 ;
        RECT 610.950 484.050 618.900 485.100 ;
        RECT 592.950 483.750 595.050 484.050 ;
        RECT 592.950 481.950 596.850 483.750 ;
        RECT 590.550 479.850 595.050 481.950 ;
        RECT 604.050 480.000 604.950 484.050 ;
        RECT 617.100 483.300 618.900 484.050 ;
        RECT 620.100 483.150 621.900 484.950 ;
        RECT 614.100 482.400 615.900 483.000 ;
        RECT 620.100 482.400 621.000 483.150 ;
        RECT 614.100 481.200 621.000 482.400 ;
        RECT 614.100 480.000 615.150 481.200 ;
        RECT 590.550 477.600 591.750 479.850 ;
        RECT 604.050 479.100 615.150 480.000 ;
        RECT 604.050 478.800 604.950 479.100 ;
        RECT 580.200 471.750 582.000 475.950 ;
        RECT 583.500 471.750 585.300 474.600 ;
        RECT 590.550 471.750 592.350 477.600 ;
        RECT 595.950 476.700 598.050 477.600 ;
        RECT 603.150 477.000 604.950 478.800 ;
        RECT 614.100 478.200 615.150 479.100 ;
        RECT 610.350 477.450 612.150 478.200 ;
        RECT 595.950 475.500 599.700 476.700 ;
        RECT 598.650 474.600 599.700 475.500 ;
        RECT 607.200 476.400 612.150 477.450 ;
        RECT 613.650 476.400 615.450 478.200 ;
        RECT 622.950 477.600 623.850 490.200 ;
        RECT 660.150 489.600 664.200 490.500 ;
        RECT 653.250 486.150 655.050 487.950 ;
        RECT 660.150 486.150 661.050 489.600 ;
        RECT 665.100 486.150 666.900 487.950 ;
        RECT 707.700 486.150 708.900 491.400 ;
        RECT 740.100 486.150 741.900 487.950 ;
        RECT 745.950 486.150 747.150 491.400 ;
        RECT 748.950 489.150 750.750 490.950 ;
        RECT 748.950 487.050 751.050 489.150 ;
        RECT 652.950 484.050 655.050 486.150 ;
        RECT 655.950 482.850 658.050 484.950 ;
        RECT 656.250 481.050 658.050 482.850 ;
        RECT 658.950 484.050 661.050 486.150 ;
        RECT 658.950 477.600 660.000 484.050 ;
        RECT 661.950 482.850 664.050 484.950 ;
        RECT 664.950 484.050 667.050 486.150 ;
        RECT 697.950 482.850 700.050 484.950 ;
        RECT 701.100 483.150 702.900 484.950 ;
        RECT 661.950 481.050 663.750 482.850 ;
        RECT 698.100 481.050 699.900 482.850 ;
        RECT 700.950 481.050 703.050 483.150 ;
        RECT 703.950 482.850 706.050 484.950 ;
        RECT 706.950 484.050 709.050 486.150 ;
        RECT 739.950 484.050 742.050 486.150 ;
        RECT 704.100 481.050 705.900 482.850 ;
        RECT 707.700 477.600 708.900 484.050 ;
        RECT 742.950 482.850 745.050 484.950 ;
        RECT 745.950 484.050 748.050 486.150 ;
        RECT 743.100 481.050 744.900 482.850 ;
        RECT 746.850 480.750 748.050 484.050 ;
        RECT 747.000 479.700 750.750 480.750 ;
        RECT 607.200 474.600 608.250 476.400 ;
        RECT 616.950 475.500 619.050 477.600 ;
        RECT 616.950 474.600 618.000 475.500 ;
        RECT 593.850 471.750 595.650 474.600 ;
        RECT 598.350 471.750 600.150 474.600 ;
        RECT 602.550 471.750 604.350 474.600 ;
        RECT 606.450 471.750 608.250 474.600 ;
        RECT 609.750 471.750 611.550 474.600 ;
        RECT 614.250 473.700 618.000 474.600 ;
        RECT 614.250 471.750 616.050 473.700 ;
        RECT 619.050 471.750 620.850 474.600 ;
        RECT 622.050 471.750 623.850 477.600 ;
        RECT 654.000 471.750 655.800 477.600 ;
        RECT 658.200 471.750 660.000 477.600 ;
        RECT 662.400 471.750 664.200 477.600 ;
        RECT 699.000 471.750 700.800 477.600 ;
        RECT 703.200 475.950 708.900 477.600 ;
        RECT 740.550 476.700 748.350 478.050 ;
        RECT 703.200 471.750 705.000 475.950 ;
        RECT 706.500 471.750 708.300 474.600 ;
        RECT 740.550 471.750 742.350 476.700 ;
        RECT 743.550 471.750 745.350 475.800 ;
        RECT 746.550 471.750 748.350 476.700 ;
        RECT 749.550 477.600 750.750 479.700 ;
        RECT 749.550 471.750 751.350 477.600 ;
        RECT 29.550 464.400 31.350 467.250 ;
        RECT 32.550 464.400 34.350 467.250 ;
        RECT 35.550 464.400 37.350 467.250 ;
        RECT 70.650 464.400 72.450 467.250 ;
        RECT 73.650 464.400 75.450 467.250 ;
        RECT 33.000 457.950 34.050 464.400 ;
        RECT 31.950 455.850 34.050 457.950 ;
        RECT 71.400 456.150 72.600 464.400 ;
        RECT 105.000 461.400 106.800 467.250 ;
        RECT 109.200 463.050 111.000 467.250 ;
        RECT 112.500 464.400 114.300 467.250 ;
        RECT 109.200 461.400 114.900 463.050 ;
        RECT 28.950 452.850 31.050 454.950 ;
        RECT 29.100 451.050 30.900 452.850 ;
        RECT 33.000 448.650 34.050 455.850 ;
        RECT 34.950 452.850 37.050 454.950 ;
        RECT 70.950 454.050 73.050 456.150 ;
        RECT 73.950 455.850 76.050 457.950 ;
        RECT 104.100 456.150 105.900 457.950 ;
        RECT 74.100 454.050 75.900 455.850 ;
        RECT 103.950 454.050 106.050 456.150 ;
        RECT 106.950 455.850 109.050 457.950 ;
        RECT 110.100 456.150 111.900 457.950 ;
        RECT 107.100 454.050 108.900 455.850 ;
        RECT 109.950 454.050 112.050 456.150 ;
        RECT 113.700 454.950 114.900 461.400 ;
        RECT 146.550 462.300 148.350 467.250 ;
        RECT 149.550 463.200 151.350 467.250 ;
        RECT 152.550 462.300 154.350 467.250 ;
        RECT 146.550 460.950 154.350 462.300 ;
        RECT 155.550 461.400 157.350 467.250 ;
        RECT 188.550 461.400 190.350 467.250 ;
        RECT 191.550 461.400 193.350 467.250 ;
        RECT 194.550 461.400 196.350 467.250 ;
        RECT 155.550 459.300 156.750 461.400 ;
        RECT 191.400 460.500 193.200 461.400 ;
        RECT 197.550 460.500 199.350 467.250 ;
        RECT 200.550 461.400 202.350 467.250 ;
        RECT 203.550 461.400 205.350 467.250 ;
        RECT 206.550 461.400 208.350 467.250 ;
        RECT 209.550 461.400 211.350 467.250 ;
        RECT 212.550 461.400 214.350 467.250 ;
        RECT 245.550 464.400 247.350 467.250 ;
        RECT 248.550 464.400 250.350 467.250 ;
        RECT 281.550 464.400 283.350 467.250 ;
        RECT 203.400 460.500 205.200 461.400 ;
        RECT 209.400 460.500 211.200 461.400 ;
        RECT 191.400 459.300 195.450 460.500 ;
        RECT 197.550 459.300 201.300 460.500 ;
        RECT 203.400 459.300 207.300 460.500 ;
        RECT 209.400 460.350 212.100 460.500 ;
        RECT 209.400 459.300 212.250 460.350 ;
        RECT 153.000 458.250 156.750 459.300 ;
        RECT 194.250 458.400 195.450 459.300 ;
        RECT 200.100 458.400 201.300 459.300 ;
        RECT 206.100 458.400 207.300 459.300 ;
        RECT 149.100 456.150 150.900 457.950 ;
        RECT 35.100 451.050 36.900 452.850 ;
        RECT 33.000 447.600 35.550 448.650 ;
        RECT 29.550 435.750 31.350 447.600 ;
        RECT 33.750 435.750 35.550 447.600 ;
        RECT 71.400 441.600 72.600 454.050 ;
        RECT 112.950 452.850 115.050 454.950 ;
        RECT 145.950 452.850 148.050 454.950 ;
        RECT 148.950 454.050 151.050 456.150 ;
        RECT 152.850 454.950 154.050 458.250 ;
        RECT 191.100 456.150 192.900 457.950 ;
        RECT 194.250 456.600 198.300 458.400 ;
        RECT 200.100 456.600 204.300 458.400 ;
        RECT 206.100 456.600 210.300 458.400 ;
        RECT 151.950 452.850 154.050 454.950 ;
        RECT 190.950 454.050 193.050 456.150 ;
        RECT 113.700 447.600 114.900 452.850 ;
        RECT 146.100 451.050 147.900 452.850 ;
        RECT 151.950 447.600 153.150 452.850 ;
        RECT 154.950 449.850 157.050 451.950 ;
        RECT 154.950 448.050 156.750 449.850 ;
        RECT 194.250 449.700 195.450 456.600 ;
        RECT 200.100 449.700 201.300 456.600 ;
        RECT 206.100 449.700 207.300 456.600 ;
        RECT 211.200 456.150 212.250 459.300 ;
        RECT 211.200 454.050 214.050 456.150 ;
        RECT 244.950 455.850 247.050 457.950 ;
        RECT 248.400 456.150 249.600 464.400 ;
        RECT 282.150 460.500 283.350 464.400 ;
        RECT 284.850 461.400 286.650 467.250 ;
        RECT 287.850 461.400 289.650 467.250 ;
        RECT 294.150 461.400 295.950 467.250 ;
        RECT 297.150 464.400 298.950 467.250 ;
        RECT 301.950 465.300 303.750 467.250 ;
        RECT 300.000 464.400 303.750 465.300 ;
        RECT 306.450 464.400 308.250 467.250 ;
        RECT 309.750 464.400 311.550 467.250 ;
        RECT 313.650 464.400 315.450 467.250 ;
        RECT 317.850 464.400 319.650 467.250 ;
        RECT 322.350 464.400 324.150 467.250 ;
        RECT 300.000 463.500 301.050 464.400 ;
        RECT 298.950 461.400 301.050 463.500 ;
        RECT 309.750 462.600 310.800 464.400 ;
        RECT 282.150 459.600 287.250 460.500 ;
        RECT 285.000 458.700 287.250 459.600 ;
        RECT 245.100 454.050 246.900 455.850 ;
        RECT 247.950 454.050 250.050 456.150 ;
        RECT 211.200 449.700 212.250 454.050 ;
        RECT 191.550 448.500 195.450 449.700 ;
        RECT 197.550 448.500 201.300 449.700 ;
        RECT 203.550 448.500 207.300 449.700 ;
        RECT 209.550 448.500 212.250 449.700 ;
        RECT 104.550 446.700 112.350 447.600 ;
        RECT 70.650 435.750 72.450 441.600 ;
        RECT 73.650 435.750 75.450 441.600 ;
        RECT 104.550 435.750 106.350 446.700 ;
        RECT 107.550 435.750 109.350 445.800 ;
        RECT 110.550 435.750 112.350 446.700 ;
        RECT 113.550 435.750 115.350 447.600 ;
        RECT 147.300 435.750 149.100 447.600 ;
        RECT 151.500 435.750 153.300 447.600 ;
        RECT 154.800 435.750 156.600 441.600 ;
        RECT 188.550 435.750 190.350 447.600 ;
        RECT 191.550 435.750 193.350 448.500 ;
        RECT 194.550 435.750 196.350 447.600 ;
        RECT 197.550 435.750 199.350 448.500 ;
        RECT 200.550 435.750 202.350 447.600 ;
        RECT 203.550 435.750 205.350 448.500 ;
        RECT 206.550 435.750 208.350 447.600 ;
        RECT 209.550 435.750 211.350 448.500 ;
        RECT 212.550 435.750 214.350 447.600 ;
        RECT 248.400 441.600 249.600 454.050 ;
        RECT 280.950 452.850 283.050 454.950 ;
        RECT 281.100 451.050 282.900 452.850 ;
        RECT 285.000 450.300 286.050 458.700 ;
        RECT 288.150 454.950 289.350 461.400 ;
        RECT 286.950 452.850 289.350 454.950 ;
        RECT 285.000 449.400 287.250 450.300 ;
        RECT 281.550 448.500 287.250 449.400 ;
        RECT 281.550 441.600 282.750 448.500 ;
        RECT 288.150 447.600 289.350 452.850 ;
        RECT 294.150 448.800 295.050 461.400 ;
        RECT 302.550 460.800 304.350 462.600 ;
        RECT 305.850 461.550 310.800 462.600 ;
        RECT 318.300 463.500 319.350 464.400 ;
        RECT 318.300 462.300 322.050 463.500 ;
        RECT 305.850 460.800 307.650 461.550 ;
        RECT 302.850 459.900 303.900 460.800 ;
        RECT 313.050 460.200 314.850 462.000 ;
        RECT 319.950 461.400 322.050 462.300 ;
        RECT 325.650 461.400 327.450 467.250 ;
        RECT 356.550 464.400 358.350 467.250 ;
        RECT 359.550 464.400 361.350 467.250 ;
        RECT 313.050 459.900 313.950 460.200 ;
        RECT 302.850 459.000 313.950 459.900 ;
        RECT 326.250 459.150 327.450 461.400 ;
        RECT 302.850 457.800 303.900 459.000 ;
        RECT 297.000 456.600 303.900 457.800 ;
        RECT 297.000 455.850 297.900 456.600 ;
        RECT 302.100 456.000 303.900 456.600 ;
        RECT 296.100 454.050 297.900 455.850 ;
        RECT 299.100 454.950 300.900 455.700 ;
        RECT 313.050 454.950 313.950 459.000 ;
        RECT 322.950 457.050 327.450 459.150 ;
        RECT 321.150 455.250 325.050 457.050 ;
        RECT 322.950 454.950 325.050 455.250 ;
        RECT 299.100 453.900 307.050 454.950 ;
        RECT 304.950 452.850 307.050 453.900 ;
        RECT 310.950 452.850 313.950 454.950 ;
        RECT 303.450 449.100 305.250 449.400 ;
        RECT 303.450 448.800 311.850 449.100 ;
        RECT 294.150 448.200 311.850 448.800 ;
        RECT 294.150 447.600 305.250 448.200 ;
        RECT 245.550 435.750 247.350 441.600 ;
        RECT 248.550 435.750 250.350 441.600 ;
        RECT 281.550 435.750 283.350 441.600 ;
        RECT 284.850 435.750 286.650 447.600 ;
        RECT 287.850 435.750 289.650 447.600 ;
        RECT 294.150 435.750 295.950 447.600 ;
        RECT 308.250 446.700 310.050 447.300 ;
        RECT 302.550 445.500 310.050 446.700 ;
        RECT 310.950 446.100 311.850 448.200 ;
        RECT 313.050 448.200 313.950 452.850 ;
        RECT 323.250 449.400 325.050 451.200 ;
        RECT 319.950 448.200 324.150 449.400 ;
        RECT 313.050 447.300 319.050 448.200 ;
        RECT 319.950 447.300 322.050 448.200 ;
        RECT 326.250 447.600 327.450 457.050 ;
        RECT 355.950 455.850 358.050 457.950 ;
        RECT 359.400 456.150 360.600 464.400 ;
        RECT 365.550 461.400 367.350 467.250 ;
        RECT 368.850 464.400 370.650 467.250 ;
        RECT 373.350 464.400 375.150 467.250 ;
        RECT 377.550 464.400 379.350 467.250 ;
        RECT 381.450 464.400 383.250 467.250 ;
        RECT 384.750 464.400 386.550 467.250 ;
        RECT 389.250 465.300 391.050 467.250 ;
        RECT 389.250 464.400 393.000 465.300 ;
        RECT 394.050 464.400 395.850 467.250 ;
        RECT 373.650 463.500 374.700 464.400 ;
        RECT 370.950 462.300 374.700 463.500 ;
        RECT 382.200 462.600 383.250 464.400 ;
        RECT 391.950 463.500 393.000 464.400 ;
        RECT 370.950 461.400 373.050 462.300 ;
        RECT 365.550 459.150 366.750 461.400 ;
        RECT 378.150 460.200 379.950 462.000 ;
        RECT 382.200 461.550 387.150 462.600 ;
        RECT 385.350 460.800 387.150 461.550 ;
        RECT 388.650 460.800 390.450 462.600 ;
        RECT 391.950 461.400 394.050 463.500 ;
        RECT 397.050 461.400 398.850 467.250 ;
        RECT 428.550 464.400 430.350 467.250 ;
        RECT 431.550 464.400 433.350 467.250 ;
        RECT 434.550 464.400 436.350 467.250 ;
        RECT 464.550 464.400 466.350 467.250 ;
        RECT 467.550 464.400 469.350 467.250 ;
        RECT 470.550 464.400 472.350 467.250 ;
        RECT 500.550 464.400 502.350 467.250 ;
        RECT 379.050 459.900 379.950 460.200 ;
        RECT 389.100 459.900 390.150 460.800 ;
        RECT 365.550 457.050 370.050 459.150 ;
        RECT 379.050 459.000 390.150 459.900 ;
        RECT 356.100 454.050 357.900 455.850 ;
        RECT 358.950 454.050 361.050 456.150 ;
        RECT 318.150 446.400 319.050 447.300 ;
        RECT 315.450 446.100 317.250 446.400 ;
        RECT 302.550 444.600 303.750 445.500 ;
        RECT 310.950 445.200 317.250 446.100 ;
        RECT 315.450 444.600 317.250 445.200 ;
        RECT 318.150 444.600 320.850 446.400 ;
        RECT 298.950 442.500 303.750 444.600 ;
        RECT 306.150 442.500 313.050 444.300 ;
        RECT 302.550 441.600 303.750 442.500 ;
        RECT 297.150 435.750 298.950 441.600 ;
        RECT 302.250 435.750 304.050 441.600 ;
        RECT 307.050 435.750 308.850 441.600 ;
        RECT 310.050 435.750 311.850 442.500 ;
        RECT 318.150 441.600 322.050 443.700 ;
        RECT 313.950 435.750 315.750 441.600 ;
        RECT 318.150 435.750 319.950 441.600 ;
        RECT 322.650 435.750 324.450 438.600 ;
        RECT 325.650 435.750 327.450 447.600 ;
        RECT 359.400 441.600 360.600 454.050 ;
        RECT 365.550 447.600 366.750 457.050 ;
        RECT 367.950 455.250 371.850 457.050 ;
        RECT 367.950 454.950 370.050 455.250 ;
        RECT 379.050 454.950 379.950 459.000 ;
        RECT 389.100 457.800 390.150 459.000 ;
        RECT 389.100 456.600 396.000 457.800 ;
        RECT 389.100 456.000 390.900 456.600 ;
        RECT 395.100 455.850 396.000 456.600 ;
        RECT 392.100 454.950 393.900 455.700 ;
        RECT 379.050 452.850 382.050 454.950 ;
        RECT 385.950 453.900 393.900 454.950 ;
        RECT 395.100 454.050 396.900 455.850 ;
        RECT 385.950 452.850 388.050 453.900 ;
        RECT 367.950 449.400 369.750 451.200 ;
        RECT 368.850 448.200 373.050 449.400 ;
        RECT 379.050 448.200 379.950 452.850 ;
        RECT 387.750 449.100 389.550 449.400 ;
        RECT 356.550 435.750 358.350 441.600 ;
        RECT 359.550 435.750 361.350 441.600 ;
        RECT 365.550 435.750 367.350 447.600 ;
        RECT 370.950 447.300 373.050 448.200 ;
        RECT 373.950 447.300 379.950 448.200 ;
        RECT 381.150 448.800 389.550 449.100 ;
        RECT 397.950 448.800 398.850 461.400 ;
        RECT 432.000 457.950 433.050 464.400 ;
        RECT 468.000 457.950 469.050 464.400 ;
        RECT 501.150 460.500 502.350 464.400 ;
        RECT 503.850 461.400 505.650 467.250 ;
        RECT 506.850 461.400 508.650 467.250 ;
        RECT 541.650 461.400 543.450 467.250 ;
        RECT 501.150 459.600 506.250 460.500 ;
        RECT 430.950 455.850 433.050 457.950 ;
        RECT 466.950 455.850 469.050 457.950 ;
        RECT 427.950 452.850 430.050 454.950 ;
        RECT 428.100 451.050 429.900 452.850 ;
        RECT 381.150 448.200 398.850 448.800 ;
        RECT 373.950 446.400 374.850 447.300 ;
        RECT 372.150 444.600 374.850 446.400 ;
        RECT 375.750 446.100 377.550 446.400 ;
        RECT 381.150 446.100 382.050 448.200 ;
        RECT 387.750 447.600 398.850 448.200 ;
        RECT 432.000 448.650 433.050 455.850 ;
        RECT 433.950 452.850 436.050 454.950 ;
        RECT 463.950 452.850 466.050 454.950 ;
        RECT 434.100 451.050 435.900 452.850 ;
        RECT 464.100 451.050 465.900 452.850 ;
        RECT 468.000 448.650 469.050 455.850 ;
        RECT 504.000 458.700 506.250 459.600 ;
        RECT 469.950 452.850 472.050 454.950 ;
        RECT 499.950 452.850 502.050 454.950 ;
        RECT 470.100 451.050 471.900 452.850 ;
        RECT 500.100 451.050 501.900 452.850 ;
        RECT 504.000 450.300 505.050 458.700 ;
        RECT 507.150 454.950 508.350 461.400 ;
        RECT 542.250 459.300 543.450 461.400 ;
        RECT 544.650 462.300 546.450 467.250 ;
        RECT 547.650 463.200 549.450 467.250 ;
        RECT 550.650 462.300 552.450 467.250 ;
        RECT 544.650 460.950 552.450 462.300 ;
        RECT 583.650 461.400 585.450 467.250 ;
        RECT 584.250 459.300 585.450 461.400 ;
        RECT 586.650 462.300 588.450 467.250 ;
        RECT 589.650 463.200 591.450 467.250 ;
        RECT 592.650 462.300 594.450 467.250 ;
        RECT 623.700 464.400 625.500 467.250 ;
        RECT 627.000 463.050 628.800 467.250 ;
        RECT 586.650 460.950 594.450 462.300 ;
        RECT 623.100 461.400 628.800 463.050 ;
        RECT 631.200 461.400 633.000 467.250 ;
        RECT 662.850 461.400 664.650 467.250 ;
        RECT 542.250 458.250 546.000 459.300 ;
        RECT 584.250 458.250 588.000 459.300 ;
        RECT 505.950 452.850 508.350 454.950 ;
        RECT 544.950 454.950 546.150 458.250 ;
        RECT 548.100 456.150 549.900 457.950 ;
        RECT 544.950 452.850 547.050 454.950 ;
        RECT 547.950 454.050 550.050 456.150 ;
        RECT 586.950 454.950 588.150 458.250 ;
        RECT 590.100 456.150 591.900 457.950 ;
        RECT 550.950 452.850 553.050 454.950 ;
        RECT 586.950 452.850 589.050 454.950 ;
        RECT 589.950 454.050 592.050 456.150 ;
        RECT 623.100 454.950 624.300 461.400 ;
        RECT 667.350 460.200 669.150 467.250 ;
        RECT 703.650 464.400 705.450 467.250 ;
        RECT 706.650 464.400 708.450 467.250 ;
        RECT 709.650 464.400 711.450 467.250 ;
        RECT 665.550 459.300 669.150 460.200 ;
        RECT 626.100 456.150 627.900 457.950 ;
        RECT 592.950 452.850 595.050 454.950 ;
        RECT 622.950 452.850 625.050 454.950 ;
        RECT 625.950 454.050 628.050 456.150 ;
        RECT 628.950 455.850 631.050 457.950 ;
        RECT 632.100 456.150 633.900 457.950 ;
        RECT 629.100 454.050 630.900 455.850 ;
        RECT 631.950 454.050 634.050 456.150 ;
        RECT 662.100 453.150 663.900 454.950 ;
        RECT 504.000 449.400 506.250 450.300 ;
        RECT 432.000 447.600 434.550 448.650 ;
        RECT 468.000 447.600 470.550 448.650 ;
        RECT 375.750 445.200 382.050 446.100 ;
        RECT 382.950 446.700 384.750 447.300 ;
        RECT 382.950 445.500 390.450 446.700 ;
        RECT 375.750 444.600 377.550 445.200 ;
        RECT 389.250 444.600 390.450 445.500 ;
        RECT 370.950 441.600 374.850 443.700 ;
        RECT 379.950 442.500 386.850 444.300 ;
        RECT 389.250 442.500 394.050 444.600 ;
        RECT 368.550 435.750 370.350 438.600 ;
        RECT 373.050 435.750 374.850 441.600 ;
        RECT 377.250 435.750 379.050 441.600 ;
        RECT 381.150 435.750 382.950 442.500 ;
        RECT 389.250 441.600 390.450 442.500 ;
        RECT 384.150 435.750 385.950 441.600 ;
        RECT 388.950 435.750 390.750 441.600 ;
        RECT 394.050 435.750 395.850 441.600 ;
        RECT 397.050 435.750 398.850 447.600 ;
        RECT 428.550 435.750 430.350 447.600 ;
        RECT 432.750 435.750 434.550 447.600 ;
        RECT 464.550 435.750 466.350 447.600 ;
        RECT 468.750 435.750 470.550 447.600 ;
        RECT 500.550 448.500 506.250 449.400 ;
        RECT 500.550 441.600 501.750 448.500 ;
        RECT 507.150 447.600 508.350 452.850 ;
        RECT 541.950 449.850 544.050 451.950 ;
        RECT 542.250 448.050 544.050 449.850 ;
        RECT 545.850 447.600 547.050 452.850 ;
        RECT 551.100 451.050 552.900 452.850 ;
        RECT 583.950 449.850 586.050 451.950 ;
        RECT 584.250 448.050 586.050 449.850 ;
        RECT 587.850 447.600 589.050 452.850 ;
        RECT 593.100 451.050 594.900 452.850 ;
        RECT 623.100 447.600 624.300 452.850 ;
        RECT 661.950 451.050 664.050 453.150 ;
        RECT 665.550 451.950 666.750 459.300 ;
        RECT 706.950 457.950 708.000 464.400 ;
        RECT 740.550 462.300 742.350 467.250 ;
        RECT 743.550 463.200 745.350 467.250 ;
        RECT 746.550 462.300 748.350 467.250 ;
        RECT 740.550 460.950 748.350 462.300 ;
        RECT 749.550 461.400 751.350 467.250 ;
        RECT 749.550 459.300 750.750 461.400 ;
        RECT 747.000 458.250 750.750 459.300 ;
        RECT 706.950 455.850 709.050 457.950 ;
        RECT 743.100 456.150 744.900 457.950 ;
        RECT 668.100 453.150 669.900 454.950 ;
        RECT 664.950 449.850 667.050 451.950 ;
        RECT 667.950 451.050 670.050 453.150 ;
        RECT 703.950 452.850 706.050 454.950 ;
        RECT 704.100 451.050 705.900 452.850 ;
        RECT 500.550 435.750 502.350 441.600 ;
        RECT 503.850 435.750 505.650 447.600 ;
        RECT 506.850 435.750 508.650 447.600 ;
        RECT 542.400 435.750 544.200 441.600 ;
        RECT 545.700 435.750 547.500 447.600 ;
        RECT 549.900 435.750 551.700 447.600 ;
        RECT 584.400 435.750 586.200 441.600 ;
        RECT 587.700 435.750 589.500 447.600 ;
        RECT 591.900 435.750 593.700 447.600 ;
        RECT 622.650 435.750 624.450 447.600 ;
        RECT 625.650 446.700 633.450 447.600 ;
        RECT 625.650 435.750 627.450 446.700 ;
        RECT 628.650 435.750 630.450 445.800 ;
        RECT 631.650 435.750 633.450 446.700 ;
        RECT 665.550 441.600 666.750 449.850 ;
        RECT 706.950 448.650 708.000 455.850 ;
        RECT 709.950 452.850 712.050 454.950 ;
        RECT 739.950 452.850 742.050 454.950 ;
        RECT 742.950 454.050 745.050 456.150 ;
        RECT 746.850 454.950 748.050 458.250 ;
        RECT 745.950 452.850 748.050 454.950 ;
        RECT 710.100 451.050 711.900 452.850 ;
        RECT 740.100 451.050 741.900 452.850 ;
        RECT 705.450 447.600 708.000 448.650 ;
        RECT 745.950 447.600 747.150 452.850 ;
        RECT 748.950 449.850 751.050 451.950 ;
        RECT 748.950 448.050 750.750 449.850 ;
        RECT 662.550 435.750 664.350 441.600 ;
        RECT 665.550 435.750 667.350 441.600 ;
        RECT 668.550 435.750 670.350 441.600 ;
        RECT 705.450 435.750 707.250 447.600 ;
        RECT 709.650 435.750 711.450 447.600 ;
        RECT 741.300 435.750 743.100 447.600 ;
        RECT 745.500 435.750 747.300 447.600 ;
        RECT 748.800 435.750 750.600 441.600 ;
        RECT 3.150 419.400 4.950 431.250 ;
        RECT 6.150 425.400 7.950 431.250 ;
        RECT 11.250 425.400 13.050 431.250 ;
        RECT 16.050 425.400 17.850 431.250 ;
        RECT 11.550 424.500 12.750 425.400 ;
        RECT 19.050 424.500 20.850 431.250 ;
        RECT 22.950 425.400 24.750 431.250 ;
        RECT 27.150 425.400 28.950 431.250 ;
        RECT 31.650 428.400 33.450 431.250 ;
        RECT 7.950 422.400 12.750 424.500 ;
        RECT 15.150 422.700 22.050 424.500 ;
        RECT 27.150 423.300 31.050 425.400 ;
        RECT 11.550 421.500 12.750 422.400 ;
        RECT 24.450 421.800 26.250 422.400 ;
        RECT 11.550 420.300 19.050 421.500 ;
        RECT 17.250 419.700 19.050 420.300 ;
        RECT 19.950 420.900 26.250 421.800 ;
        RECT 3.150 418.800 14.250 419.400 ;
        RECT 19.950 418.800 20.850 420.900 ;
        RECT 24.450 420.600 26.250 420.900 ;
        RECT 27.150 420.600 29.850 422.400 ;
        RECT 27.150 419.700 28.050 420.600 ;
        RECT 3.150 418.200 20.850 418.800 ;
        RECT 3.150 405.600 4.050 418.200 ;
        RECT 12.450 417.900 20.850 418.200 ;
        RECT 22.050 418.800 28.050 419.700 ;
        RECT 28.950 418.800 31.050 419.700 ;
        RECT 34.650 419.400 36.450 431.250 ;
        RECT 67.650 419.400 69.450 431.250 ;
        RECT 70.650 420.300 72.450 431.250 ;
        RECT 73.650 421.200 75.450 431.250 ;
        RECT 76.650 420.300 78.450 431.250 ;
        RECT 109.650 425.400 111.450 431.250 ;
        RECT 112.650 425.400 114.450 431.250 ;
        RECT 115.650 425.400 117.450 431.250 ;
        RECT 82.950 423.450 85.050 424.050 ;
        RECT 106.950 423.450 109.050 424.050 ;
        RECT 82.950 422.550 109.050 423.450 ;
        RECT 82.950 421.950 85.050 422.550 ;
        RECT 106.950 421.950 109.050 422.550 ;
        RECT 70.650 419.400 78.450 420.300 ;
        RECT 12.450 417.600 14.250 417.900 ;
        RECT 22.050 414.150 22.950 418.800 ;
        RECT 28.950 417.600 33.150 418.800 ;
        RECT 32.250 415.800 34.050 417.600 ;
        RECT 13.950 413.100 16.050 414.150 ;
        RECT 5.100 411.150 6.900 412.950 ;
        RECT 8.100 412.050 16.050 413.100 ;
        RECT 19.950 412.050 22.950 414.150 ;
        RECT 8.100 411.300 9.900 412.050 ;
        RECT 6.000 410.400 6.900 411.150 ;
        RECT 11.100 410.400 12.900 411.000 ;
        RECT 6.000 409.200 12.900 410.400 ;
        RECT 11.850 408.000 12.900 409.200 ;
        RECT 22.050 408.000 22.950 412.050 ;
        RECT 31.950 411.750 34.050 412.050 ;
        RECT 30.150 409.950 34.050 411.750 ;
        RECT 35.250 409.950 36.450 419.400 ;
        RECT 68.100 414.150 69.300 419.400 ;
        RECT 113.250 417.150 114.450 425.400 ;
        RECT 145.350 419.400 147.150 431.250 ;
        RECT 148.350 419.400 150.150 431.250 ;
        RECT 151.650 425.400 153.450 431.250 ;
        RECT 67.950 412.050 70.050 414.150 ;
        RECT 109.950 413.850 112.050 415.950 ;
        RECT 112.950 415.050 115.050 417.150 ;
        RECT 11.850 407.100 22.950 408.000 ;
        RECT 31.950 407.850 36.450 409.950 ;
        RECT 11.850 406.200 12.900 407.100 ;
        RECT 22.050 406.800 22.950 407.100 ;
        RECT 3.150 399.750 4.950 405.600 ;
        RECT 7.950 403.500 10.050 405.600 ;
        RECT 11.550 404.400 13.350 406.200 ;
        RECT 14.850 405.450 16.650 406.200 ;
        RECT 14.850 404.400 19.800 405.450 ;
        RECT 22.050 405.000 23.850 406.800 ;
        RECT 35.250 405.600 36.450 407.850 ;
        RECT 28.950 404.700 31.050 405.600 ;
        RECT 9.000 402.600 10.050 403.500 ;
        RECT 18.750 402.600 19.800 404.400 ;
        RECT 27.300 403.500 31.050 404.700 ;
        RECT 27.300 402.600 28.350 403.500 ;
        RECT 6.150 399.750 7.950 402.600 ;
        RECT 9.000 401.700 12.750 402.600 ;
        RECT 10.950 399.750 12.750 401.700 ;
        RECT 15.450 399.750 17.250 402.600 ;
        RECT 18.750 399.750 20.550 402.600 ;
        RECT 22.650 399.750 24.450 402.600 ;
        RECT 26.850 399.750 28.650 402.600 ;
        RECT 31.350 399.750 33.150 402.600 ;
        RECT 34.650 399.750 36.450 405.600 ;
        RECT 68.100 405.600 69.300 412.050 ;
        RECT 70.950 410.850 73.050 412.950 ;
        RECT 74.100 411.150 75.900 412.950 ;
        RECT 71.100 409.050 72.900 410.850 ;
        RECT 73.950 409.050 76.050 411.150 ;
        RECT 76.950 410.850 79.050 412.950 ;
        RECT 110.100 412.050 111.900 413.850 ;
        RECT 77.100 409.050 78.900 410.850 ;
        RECT 113.250 407.700 114.450 415.050 ;
        RECT 115.950 413.850 118.050 415.950 ;
        RECT 145.650 414.150 146.850 419.400 ;
        RECT 152.250 418.500 153.450 425.400 ;
        RECT 147.750 417.600 153.450 418.500 ;
        RECT 156.150 419.400 157.950 431.250 ;
        RECT 159.150 425.400 160.950 431.250 ;
        RECT 164.250 425.400 166.050 431.250 ;
        RECT 169.050 425.400 170.850 431.250 ;
        RECT 164.550 424.500 165.750 425.400 ;
        RECT 172.050 424.500 173.850 431.250 ;
        RECT 175.950 425.400 177.750 431.250 ;
        RECT 180.150 425.400 181.950 431.250 ;
        RECT 184.650 428.400 186.450 431.250 ;
        RECT 160.950 422.400 165.750 424.500 ;
        RECT 168.150 422.700 175.050 424.500 ;
        RECT 180.150 423.300 184.050 425.400 ;
        RECT 164.550 421.500 165.750 422.400 ;
        RECT 177.450 421.800 179.250 422.400 ;
        RECT 164.550 420.300 172.050 421.500 ;
        RECT 170.250 419.700 172.050 420.300 ;
        RECT 172.950 420.900 179.250 421.800 ;
        RECT 156.150 418.800 167.250 419.400 ;
        RECT 172.950 418.800 173.850 420.900 ;
        RECT 177.450 420.600 179.250 420.900 ;
        RECT 180.150 420.600 182.850 422.400 ;
        RECT 180.150 419.700 181.050 420.600 ;
        RECT 156.150 418.200 173.850 418.800 ;
        RECT 147.750 416.700 150.000 417.600 ;
        RECT 116.100 412.050 117.900 413.850 ;
        RECT 145.650 412.050 148.050 414.150 ;
        RECT 110.850 406.800 114.450 407.700 ;
        RECT 68.100 403.950 73.800 405.600 ;
        RECT 68.700 399.750 70.500 402.600 ;
        RECT 72.000 399.750 73.800 403.950 ;
        RECT 76.200 399.750 78.000 405.600 ;
        RECT 110.850 399.750 112.650 406.800 ;
        RECT 145.650 405.600 146.850 412.050 ;
        RECT 148.950 408.300 150.000 416.700 ;
        RECT 152.100 414.150 153.900 415.950 ;
        RECT 151.950 412.050 154.050 414.150 ;
        RECT 147.750 407.400 150.000 408.300 ;
        RECT 147.750 406.500 152.850 407.400 ;
        RECT 115.350 399.750 117.150 405.600 ;
        RECT 145.350 399.750 147.150 405.600 ;
        RECT 148.350 399.750 150.150 405.600 ;
        RECT 151.650 402.600 152.850 406.500 ;
        RECT 156.150 405.600 157.050 418.200 ;
        RECT 165.450 417.900 173.850 418.200 ;
        RECT 175.050 418.800 181.050 419.700 ;
        RECT 181.950 418.800 184.050 419.700 ;
        RECT 187.650 419.400 189.450 431.250 ;
        RECT 218.550 425.400 220.350 431.250 ;
        RECT 221.550 425.400 223.350 431.250 ;
        RECT 256.650 425.400 258.450 431.250 ;
        RECT 259.650 425.400 261.450 431.250 ;
        RECT 292.650 425.400 294.450 431.250 ;
        RECT 295.650 425.400 297.450 431.250 ;
        RECT 298.650 425.400 300.450 431.250 ;
        RECT 165.450 417.600 167.250 417.900 ;
        RECT 175.050 414.150 175.950 418.800 ;
        RECT 181.950 417.600 186.150 418.800 ;
        RECT 185.250 415.800 187.050 417.600 ;
        RECT 166.950 413.100 169.050 414.150 ;
        RECT 158.100 411.150 159.900 412.950 ;
        RECT 161.100 412.050 169.050 413.100 ;
        RECT 172.950 412.050 175.950 414.150 ;
        RECT 161.100 411.300 162.900 412.050 ;
        RECT 159.000 410.400 159.900 411.150 ;
        RECT 164.100 410.400 165.900 411.000 ;
        RECT 159.000 409.200 165.900 410.400 ;
        RECT 164.850 408.000 165.900 409.200 ;
        RECT 175.050 408.000 175.950 412.050 ;
        RECT 184.950 411.750 187.050 412.050 ;
        RECT 183.150 409.950 187.050 411.750 ;
        RECT 188.250 409.950 189.450 419.400 ;
        RECT 221.400 412.950 222.600 425.400 ;
        RECT 257.400 412.950 258.600 425.400 ;
        RECT 296.250 417.150 297.450 425.400 ;
        RECT 302.550 419.400 304.350 431.250 ;
        RECT 305.550 428.400 307.350 431.250 ;
        RECT 310.050 425.400 311.850 431.250 ;
        RECT 314.250 425.400 316.050 431.250 ;
        RECT 307.950 423.300 311.850 425.400 ;
        RECT 318.150 424.500 319.950 431.250 ;
        RECT 321.150 425.400 322.950 431.250 ;
        RECT 325.950 425.400 327.750 431.250 ;
        RECT 331.050 425.400 332.850 431.250 ;
        RECT 326.250 424.500 327.450 425.400 ;
        RECT 316.950 422.700 323.850 424.500 ;
        RECT 326.250 422.400 331.050 424.500 ;
        RECT 309.150 420.600 311.850 422.400 ;
        RECT 312.750 421.800 314.550 422.400 ;
        RECT 312.750 420.900 319.050 421.800 ;
        RECT 326.250 421.500 327.450 422.400 ;
        RECT 312.750 420.600 314.550 420.900 ;
        RECT 310.950 419.700 311.850 420.600 ;
        RECT 292.950 413.850 295.050 415.950 ;
        RECT 295.950 415.050 298.050 417.150 ;
        RECT 218.100 411.150 219.900 412.950 ;
        RECT 164.850 407.100 175.950 408.000 ;
        RECT 184.950 407.850 189.450 409.950 ;
        RECT 217.950 409.050 220.050 411.150 ;
        RECT 220.950 410.850 223.050 412.950 ;
        RECT 256.950 410.850 259.050 412.950 ;
        RECT 260.100 411.150 261.900 412.950 ;
        RECT 293.100 412.050 294.900 413.850 ;
        RECT 164.850 406.200 165.900 407.100 ;
        RECT 175.050 406.800 175.950 407.100 ;
        RECT 151.650 399.750 153.450 402.600 ;
        RECT 156.150 399.750 157.950 405.600 ;
        RECT 160.950 403.500 163.050 405.600 ;
        RECT 164.550 404.400 166.350 406.200 ;
        RECT 167.850 405.450 169.650 406.200 ;
        RECT 167.850 404.400 172.800 405.450 ;
        RECT 175.050 405.000 176.850 406.800 ;
        RECT 188.250 405.600 189.450 407.850 ;
        RECT 181.950 404.700 184.050 405.600 ;
        RECT 162.000 402.600 163.050 403.500 ;
        RECT 171.750 402.600 172.800 404.400 ;
        RECT 180.300 403.500 184.050 404.700 ;
        RECT 180.300 402.600 181.350 403.500 ;
        RECT 159.150 399.750 160.950 402.600 ;
        RECT 162.000 401.700 165.750 402.600 ;
        RECT 163.950 399.750 165.750 401.700 ;
        RECT 168.450 399.750 170.250 402.600 ;
        RECT 171.750 399.750 173.550 402.600 ;
        RECT 175.650 399.750 177.450 402.600 ;
        RECT 179.850 399.750 181.650 402.600 ;
        RECT 184.350 399.750 186.150 402.600 ;
        RECT 187.650 399.750 189.450 405.600 ;
        RECT 221.400 402.600 222.600 410.850 ;
        RECT 257.400 402.600 258.600 410.850 ;
        RECT 259.950 409.050 262.050 411.150 ;
        RECT 296.250 407.700 297.450 415.050 ;
        RECT 298.950 413.850 301.050 415.950 ;
        RECT 299.100 412.050 300.900 413.850 ;
        RECT 293.850 406.800 297.450 407.700 ;
        RECT 302.550 409.950 303.750 419.400 ;
        RECT 307.950 418.800 310.050 419.700 ;
        RECT 310.950 418.800 316.950 419.700 ;
        RECT 305.850 417.600 310.050 418.800 ;
        RECT 304.950 415.800 306.750 417.600 ;
        RECT 316.050 414.150 316.950 418.800 ;
        RECT 318.150 418.800 319.050 420.900 ;
        RECT 319.950 420.300 327.450 421.500 ;
        RECT 319.950 419.700 321.750 420.300 ;
        RECT 334.050 419.400 335.850 431.250 ;
        RECT 324.750 418.800 335.850 419.400 ;
        RECT 318.150 418.200 335.850 418.800 ;
        RECT 318.150 417.900 326.550 418.200 ;
        RECT 324.750 417.600 326.550 417.900 ;
        RECT 316.050 412.050 319.050 414.150 ;
        RECT 322.950 413.100 325.050 414.150 ;
        RECT 322.950 412.050 330.900 413.100 ;
        RECT 304.950 411.750 307.050 412.050 ;
        RECT 304.950 409.950 308.850 411.750 ;
        RECT 302.550 407.850 307.050 409.950 ;
        RECT 316.050 408.000 316.950 412.050 ;
        RECT 329.100 411.300 330.900 412.050 ;
        RECT 332.100 411.150 333.900 412.950 ;
        RECT 326.100 410.400 327.900 411.000 ;
        RECT 332.100 410.400 333.000 411.150 ;
        RECT 326.100 409.200 333.000 410.400 ;
        RECT 326.100 408.000 327.150 409.200 ;
        RECT 218.550 399.750 220.350 402.600 ;
        RECT 221.550 399.750 223.350 402.600 ;
        RECT 256.650 399.750 258.450 402.600 ;
        RECT 259.650 399.750 261.450 402.600 ;
        RECT 293.850 399.750 295.650 406.800 ;
        RECT 302.550 405.600 303.750 407.850 ;
        RECT 316.050 407.100 327.150 408.000 ;
        RECT 316.050 406.800 316.950 407.100 ;
        RECT 298.350 399.750 300.150 405.600 ;
        RECT 302.550 399.750 304.350 405.600 ;
        RECT 307.950 404.700 310.050 405.600 ;
        RECT 315.150 405.000 316.950 406.800 ;
        RECT 326.100 406.200 327.150 407.100 ;
        RECT 322.350 405.450 324.150 406.200 ;
        RECT 307.950 403.500 311.700 404.700 ;
        RECT 310.650 402.600 311.700 403.500 ;
        RECT 319.200 404.400 324.150 405.450 ;
        RECT 325.650 404.400 327.450 406.200 ;
        RECT 334.950 405.600 335.850 418.200 ;
        RECT 319.200 402.600 320.250 404.400 ;
        RECT 328.950 403.500 331.050 405.600 ;
        RECT 328.950 402.600 330.000 403.500 ;
        RECT 305.850 399.750 307.650 402.600 ;
        RECT 310.350 399.750 312.150 402.600 ;
        RECT 314.550 399.750 316.350 402.600 ;
        RECT 318.450 399.750 320.250 402.600 ;
        RECT 321.750 399.750 323.550 402.600 ;
        RECT 326.250 401.700 330.000 402.600 ;
        RECT 326.250 399.750 328.050 401.700 ;
        RECT 331.050 399.750 332.850 402.600 ;
        RECT 334.050 399.750 335.850 405.600 ;
        RECT 339.150 419.400 340.950 431.250 ;
        RECT 342.150 425.400 343.950 431.250 ;
        RECT 347.250 425.400 349.050 431.250 ;
        RECT 352.050 425.400 353.850 431.250 ;
        RECT 347.550 424.500 348.750 425.400 ;
        RECT 355.050 424.500 356.850 431.250 ;
        RECT 358.950 425.400 360.750 431.250 ;
        RECT 363.150 425.400 364.950 431.250 ;
        RECT 367.650 428.400 369.450 431.250 ;
        RECT 343.950 422.400 348.750 424.500 ;
        RECT 351.150 422.700 358.050 424.500 ;
        RECT 363.150 423.300 367.050 425.400 ;
        RECT 347.550 421.500 348.750 422.400 ;
        RECT 360.450 421.800 362.250 422.400 ;
        RECT 347.550 420.300 355.050 421.500 ;
        RECT 353.250 419.700 355.050 420.300 ;
        RECT 355.950 420.900 362.250 421.800 ;
        RECT 339.150 418.800 350.250 419.400 ;
        RECT 355.950 418.800 356.850 420.900 ;
        RECT 360.450 420.600 362.250 420.900 ;
        RECT 363.150 420.600 365.850 422.400 ;
        RECT 363.150 419.700 364.050 420.600 ;
        RECT 339.150 418.200 356.850 418.800 ;
        RECT 339.150 405.600 340.050 418.200 ;
        RECT 348.450 417.900 356.850 418.200 ;
        RECT 358.050 418.800 364.050 419.700 ;
        RECT 364.950 418.800 367.050 419.700 ;
        RECT 370.650 419.400 372.450 431.250 ;
        RECT 401.550 425.400 403.350 431.250 ;
        RECT 404.550 425.400 406.350 431.250 ;
        RECT 348.450 417.600 350.250 417.900 ;
        RECT 358.050 414.150 358.950 418.800 ;
        RECT 364.950 417.600 369.150 418.800 ;
        RECT 368.250 415.800 370.050 417.600 ;
        RECT 349.950 413.100 352.050 414.150 ;
        RECT 341.100 411.150 342.900 412.950 ;
        RECT 344.100 412.050 352.050 413.100 ;
        RECT 355.950 412.050 358.950 414.150 ;
        RECT 344.100 411.300 345.900 412.050 ;
        RECT 342.000 410.400 342.900 411.150 ;
        RECT 347.100 410.400 348.900 411.000 ;
        RECT 342.000 409.200 348.900 410.400 ;
        RECT 347.850 408.000 348.900 409.200 ;
        RECT 358.050 408.000 358.950 412.050 ;
        RECT 367.950 411.750 370.050 412.050 ;
        RECT 366.150 409.950 370.050 411.750 ;
        RECT 371.250 409.950 372.450 419.400 ;
        RECT 404.400 412.950 405.600 425.400 ;
        RECT 437.550 420.300 439.350 431.250 ;
        RECT 440.550 421.200 442.350 431.250 ;
        RECT 443.550 420.300 445.350 431.250 ;
        RECT 437.550 419.400 445.350 420.300 ;
        RECT 446.550 419.400 448.350 431.250 ;
        RECT 479.400 425.400 481.200 431.250 ;
        RECT 482.700 419.400 484.500 431.250 ;
        RECT 486.900 419.400 488.700 431.250 ;
        RECT 522.450 419.400 524.250 431.250 ;
        RECT 526.650 419.400 528.450 431.250 ;
        RECT 554.550 419.400 556.350 431.250 ;
        RECT 559.050 419.550 560.850 431.250 ;
        RECT 562.050 420.900 563.850 431.250 ;
        RECT 599.400 425.400 601.200 431.250 ;
        RECT 562.050 419.550 564.450 420.900 ;
        RECT 406.950 414.450 409.050 415.050 ;
        RECT 433.950 414.450 436.050 415.050 ;
        RECT 406.950 413.550 436.050 414.450 ;
        RECT 446.700 414.150 447.900 419.400 ;
        RECT 479.250 417.150 481.050 418.950 ;
        RECT 478.950 415.050 481.050 417.150 ;
        RECT 482.850 414.150 484.050 419.400 ;
        RECT 522.450 418.350 525.000 419.400 ;
        RECT 488.100 414.150 489.900 415.950 ;
        RECT 521.100 414.150 522.900 415.950 ;
        RECT 406.950 412.950 409.050 413.550 ;
        RECT 433.950 412.950 436.050 413.550 ;
        RECT 401.100 411.150 402.900 412.950 ;
        RECT 347.850 407.100 358.950 408.000 ;
        RECT 367.950 407.850 372.450 409.950 ;
        RECT 400.950 409.050 403.050 411.150 ;
        RECT 403.950 410.850 406.050 412.950 ;
        RECT 436.950 410.850 439.050 412.950 ;
        RECT 440.100 411.150 441.900 412.950 ;
        RECT 347.850 406.200 348.900 407.100 ;
        RECT 358.050 406.800 358.950 407.100 ;
        RECT 339.150 399.750 340.950 405.600 ;
        RECT 343.950 403.500 346.050 405.600 ;
        RECT 347.550 404.400 349.350 406.200 ;
        RECT 350.850 405.450 352.650 406.200 ;
        RECT 350.850 404.400 355.800 405.450 ;
        RECT 358.050 405.000 359.850 406.800 ;
        RECT 371.250 405.600 372.450 407.850 ;
        RECT 364.950 404.700 367.050 405.600 ;
        RECT 345.000 402.600 346.050 403.500 ;
        RECT 354.750 402.600 355.800 404.400 ;
        RECT 363.300 403.500 367.050 404.700 ;
        RECT 363.300 402.600 364.350 403.500 ;
        RECT 342.150 399.750 343.950 402.600 ;
        RECT 345.000 401.700 348.750 402.600 ;
        RECT 346.950 399.750 348.750 401.700 ;
        RECT 351.450 399.750 353.250 402.600 ;
        RECT 354.750 399.750 356.550 402.600 ;
        RECT 358.650 399.750 360.450 402.600 ;
        RECT 362.850 399.750 364.650 402.600 ;
        RECT 367.350 399.750 369.150 402.600 ;
        RECT 370.650 399.750 372.450 405.600 ;
        RECT 404.400 402.600 405.600 410.850 ;
        RECT 437.100 409.050 438.900 410.850 ;
        RECT 439.950 409.050 442.050 411.150 ;
        RECT 442.950 410.850 445.050 412.950 ;
        RECT 445.950 412.050 448.050 414.150 ;
        RECT 481.950 412.050 484.050 414.150 ;
        RECT 443.100 409.050 444.900 410.850 ;
        RECT 446.700 405.600 447.900 412.050 ;
        RECT 481.950 408.750 483.150 412.050 ;
        RECT 484.950 410.850 487.050 412.950 ;
        RECT 487.950 412.050 490.050 414.150 ;
        RECT 520.950 412.050 523.050 414.150 ;
        RECT 523.950 411.150 525.000 418.350 ;
        RECT 554.550 418.200 555.750 419.400 ;
        RECT 559.950 418.200 561.750 418.650 ;
        RECT 554.550 417.000 561.750 418.200 ;
        RECT 559.950 416.850 561.750 417.000 ;
        RECT 527.100 414.150 528.900 415.950 ;
        RECT 557.100 414.150 558.900 415.950 ;
        RECT 526.950 412.050 529.050 414.150 ;
        RECT 554.100 411.150 555.900 412.950 ;
        RECT 556.950 412.050 559.050 414.150 ;
        RECT 485.100 409.050 486.900 410.850 ;
        RECT 523.950 409.050 526.050 411.150 ;
        RECT 553.950 409.050 556.050 411.150 ;
        RECT 479.250 407.700 483.000 408.750 ;
        RECT 479.250 405.600 480.450 407.700 ;
        RECT 401.550 399.750 403.350 402.600 ;
        RECT 404.550 399.750 406.350 402.600 ;
        RECT 438.000 399.750 439.800 405.600 ;
        RECT 442.200 403.950 447.900 405.600 ;
        RECT 442.200 399.750 444.000 403.950 ;
        RECT 445.500 399.750 447.300 402.600 ;
        RECT 478.650 399.750 480.450 405.600 ;
        RECT 481.650 404.700 489.450 406.050 ;
        RECT 481.650 399.750 483.450 404.700 ;
        RECT 484.650 399.750 486.450 403.800 ;
        RECT 487.650 399.750 489.450 404.700 ;
        RECT 523.950 402.600 525.000 409.050 ;
        RECT 560.700 408.600 561.600 416.850 ;
        RECT 563.100 412.950 564.450 419.550 ;
        RECT 602.700 419.400 604.500 431.250 ;
        RECT 606.900 419.400 608.700 431.250 ;
        RECT 638.550 425.400 640.350 431.250 ;
        RECT 641.550 425.400 643.350 431.250 ;
        RECT 644.550 425.400 646.350 431.250 ;
        RECT 599.250 417.150 601.050 418.950 ;
        RECT 598.950 415.050 601.050 417.150 ;
        RECT 602.850 414.150 604.050 419.400 ;
        RECT 641.550 417.150 642.750 425.400 ;
        RECT 674.550 420.300 676.350 431.250 ;
        RECT 677.550 421.200 679.350 431.250 ;
        RECT 680.550 420.300 682.350 431.250 ;
        RECT 674.550 419.400 682.350 420.300 ;
        RECT 683.550 419.400 685.350 431.250 ;
        RECT 716.550 420.300 718.350 431.250 ;
        RECT 719.550 421.200 721.350 431.250 ;
        RECT 722.550 420.300 724.350 431.250 ;
        RECT 716.550 419.400 724.350 420.300 ;
        RECT 725.550 419.400 727.350 431.250 ;
        RECT 608.100 414.150 609.900 415.950 ;
        RECT 562.950 410.850 565.050 412.950 ;
        RECT 559.950 407.700 561.750 408.600 ;
        RECT 558.450 406.800 561.750 407.700 ;
        RECT 558.450 402.600 559.350 406.800 ;
        RECT 564.000 405.600 565.050 410.850 ;
        RECT 601.950 412.050 604.050 414.150 ;
        RECT 601.950 408.750 603.150 412.050 ;
        RECT 604.950 410.850 607.050 412.950 ;
        RECT 607.950 412.050 610.050 414.150 ;
        RECT 637.950 413.850 640.050 415.950 ;
        RECT 640.950 415.050 643.050 417.150 ;
        RECT 638.100 412.050 639.900 413.850 ;
        RECT 605.100 409.050 606.900 410.850 ;
        RECT 599.250 407.700 603.000 408.750 ;
        RECT 641.550 407.700 642.750 415.050 ;
        RECT 643.950 413.850 646.050 415.950 ;
        RECT 683.700 414.150 684.900 419.400 ;
        RECT 725.700 414.150 726.900 419.400 ;
        RECT 644.100 412.050 645.900 413.850 ;
        RECT 673.950 410.850 676.050 412.950 ;
        RECT 677.100 411.150 678.900 412.950 ;
        RECT 674.100 409.050 675.900 410.850 ;
        RECT 676.950 409.050 679.050 411.150 ;
        RECT 679.950 410.850 682.050 412.950 ;
        RECT 682.950 412.050 685.050 414.150 ;
        RECT 680.100 409.050 681.900 410.850 ;
        RECT 599.250 405.600 600.450 407.700 ;
        RECT 641.550 406.800 645.150 407.700 ;
        RECT 520.650 399.750 522.450 402.600 ;
        RECT 523.650 399.750 525.450 402.600 ;
        RECT 526.650 399.750 528.450 402.600 ;
        RECT 554.550 399.750 556.350 402.600 ;
        RECT 557.550 399.750 559.350 402.600 ;
        RECT 560.550 399.750 562.350 402.600 ;
        RECT 563.550 399.750 565.350 405.600 ;
        RECT 598.650 399.750 600.450 405.600 ;
        RECT 601.650 404.700 609.450 406.050 ;
        RECT 601.650 399.750 603.450 404.700 ;
        RECT 604.650 399.750 606.450 403.800 ;
        RECT 607.650 399.750 609.450 404.700 ;
        RECT 638.850 399.750 640.650 405.600 ;
        RECT 643.350 399.750 645.150 406.800 ;
        RECT 683.700 405.600 684.900 412.050 ;
        RECT 715.950 410.850 718.050 412.950 ;
        RECT 719.100 411.150 720.900 412.950 ;
        RECT 716.100 409.050 717.900 410.850 ;
        RECT 718.950 409.050 721.050 411.150 ;
        RECT 721.950 410.850 724.050 412.950 ;
        RECT 724.950 412.050 727.050 414.150 ;
        RECT 722.100 409.050 723.900 410.850 ;
        RECT 725.700 405.600 726.900 412.050 ;
        RECT 675.000 399.750 676.800 405.600 ;
        RECT 679.200 403.950 684.900 405.600 ;
        RECT 679.200 399.750 681.000 403.950 ;
        RECT 682.500 399.750 684.300 402.600 ;
        RECT 717.000 399.750 718.800 405.600 ;
        RECT 721.200 403.950 726.900 405.600 ;
        RECT 721.200 399.750 723.000 403.950 ;
        RECT 724.500 399.750 726.300 402.600 ;
        RECT 28.650 389.400 30.450 395.250 ;
        RECT 29.250 387.300 30.450 389.400 ;
        RECT 31.650 390.300 33.450 395.250 ;
        RECT 34.650 391.200 36.450 395.250 ;
        RECT 37.650 390.300 39.450 395.250 ;
        RECT 31.650 388.950 39.450 390.300 ;
        RECT 71.850 388.200 73.650 395.250 ;
        RECT 76.350 389.400 78.150 395.250 ;
        RECT 71.850 387.300 75.450 388.200 ;
        RECT 29.250 386.250 33.000 387.300 ;
        RECT 31.950 382.950 33.150 386.250 ;
        RECT 35.100 384.150 36.900 385.950 ;
        RECT 31.950 380.850 34.050 382.950 ;
        RECT 34.950 382.050 37.050 384.150 ;
        RECT 37.950 380.850 40.050 382.950 ;
        RECT 71.100 381.150 72.900 382.950 ;
        RECT 28.950 377.850 31.050 379.950 ;
        RECT 29.250 376.050 31.050 377.850 ;
        RECT 32.850 375.600 34.050 380.850 ;
        RECT 38.100 379.050 39.900 380.850 ;
        RECT 70.950 379.050 73.050 381.150 ;
        RECT 74.250 379.950 75.450 387.300 ;
        RECT 107.550 387.900 109.350 395.250 ;
        RECT 112.050 389.400 113.850 395.250 ;
        RECT 115.050 390.900 116.850 395.250 ;
        RECT 115.050 389.400 118.350 390.900 ;
        RECT 151.650 389.400 153.450 395.250 ;
        RECT 154.650 389.400 156.450 395.250 ;
        RECT 187.650 392.400 189.450 395.250 ;
        RECT 190.650 392.400 192.450 395.250 ;
        RECT 193.650 392.400 195.450 395.250 ;
        RECT 113.250 387.900 115.050 388.500 ;
        RECT 107.550 386.700 115.050 387.900 ;
        RECT 77.100 381.150 78.900 382.950 ;
        RECT 73.950 377.850 76.050 379.950 ;
        RECT 76.950 379.050 79.050 381.150 ;
        RECT 106.950 380.850 109.050 382.950 ;
        RECT 107.100 379.050 108.900 380.850 ;
        RECT 29.400 363.750 31.200 369.600 ;
        RECT 32.700 363.750 34.500 375.600 ;
        RECT 36.900 363.750 38.700 375.600 ;
        RECT 74.250 369.600 75.450 377.850 ;
        RECT 110.700 369.600 111.900 386.700 ;
        RECT 117.150 382.950 118.350 389.400 ;
        RECT 152.400 382.950 153.600 389.400 ;
        RECT 190.950 385.950 192.000 392.400 ;
        RECT 227.850 388.200 229.650 395.250 ;
        RECT 232.350 389.400 234.150 395.250 ;
        RECT 260.550 390.300 262.350 395.250 ;
        RECT 263.550 391.200 265.350 395.250 ;
        RECT 266.550 390.300 268.350 395.250 ;
        RECT 260.550 388.950 268.350 390.300 ;
        RECT 269.550 389.400 271.350 395.250 ;
        RECT 303.000 389.400 304.800 395.250 ;
        RECT 307.200 391.050 309.000 395.250 ;
        RECT 310.500 392.400 312.300 395.250 ;
        RECT 341.550 392.400 343.350 395.250 ;
        RECT 344.550 392.400 346.350 395.250 ;
        RECT 347.550 392.400 349.350 395.250 ;
        RECT 377.550 392.400 379.350 395.250 ;
        RECT 307.200 389.400 312.900 391.050 ;
        RECT 227.850 387.300 231.450 388.200 ;
        RECT 269.550 387.300 270.750 389.400 ;
        RECT 155.100 384.150 156.900 385.950 ;
        RECT 113.100 381.150 114.900 382.950 ;
        RECT 112.950 379.050 115.050 381.150 ;
        RECT 115.950 380.850 118.350 382.950 ;
        RECT 151.950 380.850 154.050 382.950 ;
        RECT 154.950 382.050 157.050 384.150 ;
        RECT 190.950 383.850 193.050 385.950 ;
        RECT 187.950 380.850 190.050 382.950 ;
        RECT 117.150 375.600 118.350 380.850 ;
        RECT 152.400 375.600 153.600 380.850 ;
        RECT 188.100 379.050 189.900 380.850 ;
        RECT 190.950 376.650 192.000 383.850 ;
        RECT 193.950 380.850 196.050 382.950 ;
        RECT 227.100 381.150 228.900 382.950 ;
        RECT 194.100 379.050 195.900 380.850 ;
        RECT 226.950 379.050 229.050 381.150 ;
        RECT 230.250 379.950 231.450 387.300 ;
        RECT 267.000 386.250 270.750 387.300 ;
        RECT 263.100 384.150 264.900 385.950 ;
        RECT 233.100 381.150 234.900 382.950 ;
        RECT 229.950 377.850 232.050 379.950 ;
        RECT 232.950 379.050 235.050 381.150 ;
        RECT 259.950 380.850 262.050 382.950 ;
        RECT 262.950 382.050 265.050 384.150 ;
        RECT 266.850 382.950 268.050 386.250 ;
        RECT 302.100 384.150 303.900 385.950 ;
        RECT 265.950 380.850 268.050 382.950 ;
        RECT 301.950 382.050 304.050 384.150 ;
        RECT 304.950 383.850 307.050 385.950 ;
        RECT 308.100 384.150 309.900 385.950 ;
        RECT 305.100 382.050 306.900 383.850 ;
        RECT 307.950 382.050 310.050 384.150 ;
        RECT 311.700 382.950 312.900 389.400 ;
        RECT 345.000 385.950 346.050 392.400 ;
        RECT 378.150 388.500 379.350 392.400 ;
        RECT 380.850 389.400 382.650 395.250 ;
        RECT 383.850 389.400 385.650 395.250 ;
        RECT 378.150 387.600 383.250 388.500 ;
        RECT 343.950 383.850 346.050 385.950 ;
        RECT 310.950 380.850 313.050 382.950 ;
        RECT 340.950 380.850 343.050 382.950 ;
        RECT 260.100 379.050 261.900 380.850 ;
        RECT 189.450 375.600 192.000 376.650 ;
        RECT 70.650 363.750 72.450 369.600 ;
        RECT 73.650 363.750 75.450 369.600 ;
        RECT 76.650 363.750 78.450 369.600 ;
        RECT 107.550 363.750 109.350 369.600 ;
        RECT 110.550 363.750 112.350 369.600 ;
        RECT 114.150 363.750 115.950 375.600 ;
        RECT 117.150 363.750 118.950 375.600 ;
        RECT 151.650 363.750 153.450 375.600 ;
        RECT 154.650 363.750 156.450 375.600 ;
        RECT 189.450 363.750 191.250 375.600 ;
        RECT 193.650 363.750 195.450 375.600 ;
        RECT 230.250 369.600 231.450 377.850 ;
        RECT 265.950 375.600 267.150 380.850 ;
        RECT 268.950 377.850 271.050 379.950 ;
        RECT 268.950 376.050 270.750 377.850 ;
        RECT 311.700 375.600 312.900 380.850 ;
        RECT 341.100 379.050 342.900 380.850 ;
        RECT 345.000 376.650 346.050 383.850 ;
        RECT 381.000 386.700 383.250 387.600 ;
        RECT 346.950 380.850 349.050 382.950 ;
        RECT 376.950 380.850 379.050 382.950 ;
        RECT 347.100 379.050 348.900 380.850 ;
        RECT 377.100 379.050 378.900 380.850 ;
        RECT 381.000 378.300 382.050 386.700 ;
        RECT 384.150 382.950 385.350 389.400 ;
        RECT 419.850 388.200 421.650 395.250 ;
        RECT 424.350 389.400 426.150 395.250 ;
        RECT 457.650 389.400 459.450 395.250 ;
        RECT 419.850 387.300 423.450 388.200 ;
        RECT 382.950 380.850 385.350 382.950 ;
        RECT 419.100 381.150 420.900 382.950 ;
        RECT 381.000 377.400 383.250 378.300 ;
        RECT 345.000 375.600 347.550 376.650 ;
        RECT 226.650 363.750 228.450 369.600 ;
        RECT 229.650 363.750 231.450 369.600 ;
        RECT 232.650 363.750 234.450 369.600 ;
        RECT 261.300 363.750 263.100 375.600 ;
        RECT 265.500 363.750 267.300 375.600 ;
        RECT 302.550 374.700 310.350 375.600 ;
        RECT 268.800 363.750 270.600 369.600 ;
        RECT 302.550 363.750 304.350 374.700 ;
        RECT 305.550 363.750 307.350 373.800 ;
        RECT 308.550 363.750 310.350 374.700 ;
        RECT 311.550 363.750 313.350 375.600 ;
        RECT 341.550 363.750 343.350 375.600 ;
        RECT 345.750 363.750 347.550 375.600 ;
        RECT 377.550 376.500 383.250 377.400 ;
        RECT 377.550 369.600 378.750 376.500 ;
        RECT 384.150 375.600 385.350 380.850 ;
        RECT 418.950 379.050 421.050 381.150 ;
        RECT 422.250 379.950 423.450 387.300 ;
        RECT 458.250 387.300 459.450 389.400 ;
        RECT 460.650 390.300 462.450 395.250 ;
        RECT 463.650 391.200 465.450 395.250 ;
        RECT 466.650 390.300 468.450 395.250 ;
        RECT 460.650 388.950 468.450 390.300 ;
        RECT 498.000 389.400 499.800 395.250 ;
        RECT 502.200 391.050 504.000 395.250 ;
        RECT 505.500 392.400 507.300 395.250 ;
        RECT 502.200 389.400 507.900 391.050 ;
        RECT 541.650 389.400 543.450 395.250 ;
        RECT 458.250 386.250 462.000 387.300 ;
        RECT 460.950 382.950 462.150 386.250 ;
        RECT 464.100 384.150 465.900 385.950 ;
        RECT 497.100 384.150 498.900 385.950 ;
        RECT 425.100 381.150 426.900 382.950 ;
        RECT 421.950 377.850 424.050 379.950 ;
        RECT 424.950 379.050 427.050 381.150 ;
        RECT 460.950 380.850 463.050 382.950 ;
        RECT 463.950 382.050 466.050 384.150 ;
        RECT 466.950 380.850 469.050 382.950 ;
        RECT 496.950 382.050 499.050 384.150 ;
        RECT 499.950 383.850 502.050 385.950 ;
        RECT 503.100 384.150 504.900 385.950 ;
        RECT 500.100 382.050 501.900 383.850 ;
        RECT 502.950 382.050 505.050 384.150 ;
        RECT 506.700 382.950 507.900 389.400 ;
        RECT 542.250 387.300 543.450 389.400 ;
        RECT 544.650 390.300 546.450 395.250 ;
        RECT 547.650 391.200 549.450 395.250 ;
        RECT 550.650 390.300 552.450 395.250 ;
        RECT 583.650 392.400 585.450 395.250 ;
        RECT 586.650 392.400 588.450 395.250 ;
        RECT 589.650 392.400 591.450 395.250 ;
        RECT 620.550 392.400 622.350 395.250 ;
        RECT 623.550 392.400 625.350 395.250 ;
        RECT 544.650 388.950 552.450 390.300 ;
        RECT 571.950 387.450 574.050 388.050 ;
        RECT 583.950 387.450 586.050 388.050 ;
        RECT 542.250 386.250 546.000 387.300 ;
        RECT 571.950 386.550 586.050 387.450 ;
        RECT 544.950 382.950 546.150 386.250 ;
        RECT 571.950 385.950 574.050 386.550 ;
        RECT 583.950 385.950 586.050 386.550 ;
        RECT 586.950 385.950 588.000 392.400 ;
        RECT 548.100 384.150 549.900 385.950 ;
        RECT 505.950 380.850 508.050 382.950 ;
        RECT 544.950 380.850 547.050 382.950 ;
        RECT 547.950 382.050 550.050 384.150 ;
        RECT 586.950 383.850 589.050 385.950 ;
        RECT 619.950 383.850 622.050 385.950 ;
        RECT 623.400 384.150 624.600 392.400 ;
        RECT 658.650 389.400 660.450 395.250 ;
        RECT 659.250 387.300 660.450 389.400 ;
        RECT 661.650 390.300 663.450 395.250 ;
        RECT 664.650 391.200 666.450 395.250 ;
        RECT 667.650 390.300 669.450 395.250 ;
        RECT 698.550 392.400 700.350 395.250 ;
        RECT 701.550 392.400 703.350 395.250 ;
        RECT 731.550 392.400 733.350 395.250 ;
        RECT 734.550 392.400 736.350 395.250 ;
        RECT 661.650 388.950 669.450 390.300 ;
        RECT 659.250 386.250 663.000 387.300 ;
        RECT 550.950 380.850 553.050 382.950 ;
        RECT 583.950 380.850 586.050 382.950 ;
        RECT 457.950 377.850 460.050 379.950 ;
        RECT 377.550 363.750 379.350 369.600 ;
        RECT 380.850 363.750 382.650 375.600 ;
        RECT 383.850 363.750 385.650 375.600 ;
        RECT 422.250 369.600 423.450 377.850 ;
        RECT 458.250 376.050 460.050 377.850 ;
        RECT 461.850 375.600 463.050 380.850 ;
        RECT 467.100 379.050 468.900 380.850 ;
        RECT 506.700 375.600 507.900 380.850 ;
        RECT 541.950 377.850 544.050 379.950 ;
        RECT 542.250 376.050 544.050 377.850 ;
        RECT 545.850 375.600 547.050 380.850 ;
        RECT 551.100 379.050 552.900 380.850 ;
        RECT 584.100 379.050 585.900 380.850 ;
        RECT 586.950 376.650 588.000 383.850 ;
        RECT 589.950 380.850 592.050 382.950 ;
        RECT 620.100 382.050 621.900 383.850 ;
        RECT 622.950 382.050 625.050 384.150 ;
        RECT 661.950 382.950 663.150 386.250 ;
        RECT 665.100 384.150 666.900 385.950 ;
        RECT 590.100 379.050 591.900 380.850 ;
        RECT 585.450 375.600 588.000 376.650 ;
        RECT 418.650 363.750 420.450 369.600 ;
        RECT 421.650 363.750 423.450 369.600 ;
        RECT 424.650 363.750 426.450 369.600 ;
        RECT 458.400 363.750 460.200 369.600 ;
        RECT 461.700 363.750 463.500 375.600 ;
        RECT 465.900 363.750 467.700 375.600 ;
        RECT 497.550 374.700 505.350 375.600 ;
        RECT 497.550 363.750 499.350 374.700 ;
        RECT 500.550 363.750 502.350 373.800 ;
        RECT 503.550 363.750 505.350 374.700 ;
        RECT 506.550 363.750 508.350 375.600 ;
        RECT 542.400 363.750 544.200 369.600 ;
        RECT 545.700 363.750 547.500 375.600 ;
        RECT 549.900 363.750 551.700 375.600 ;
        RECT 585.450 363.750 587.250 375.600 ;
        RECT 589.650 363.750 591.450 375.600 ;
        RECT 623.400 369.600 624.600 382.050 ;
        RECT 661.950 380.850 664.050 382.950 ;
        RECT 664.950 382.050 667.050 384.150 ;
        RECT 697.950 383.850 700.050 385.950 ;
        RECT 701.400 384.150 702.600 392.400 ;
        RECT 667.950 380.850 670.050 382.950 ;
        RECT 698.100 382.050 699.900 383.850 ;
        RECT 700.950 382.050 703.050 384.150 ;
        RECT 730.950 383.850 733.050 385.950 ;
        RECT 734.400 384.150 735.600 392.400 ;
        RECT 731.100 382.050 732.900 383.850 ;
        RECT 733.950 382.050 736.050 384.150 ;
        RECT 658.950 377.850 661.050 379.950 ;
        RECT 659.250 376.050 661.050 377.850 ;
        RECT 662.850 375.600 664.050 380.850 ;
        RECT 668.100 379.050 669.900 380.850 ;
        RECT 620.550 363.750 622.350 369.600 ;
        RECT 623.550 363.750 625.350 369.600 ;
        RECT 659.400 363.750 661.200 369.600 ;
        RECT 662.700 363.750 664.500 375.600 ;
        RECT 666.900 363.750 668.700 375.600 ;
        RECT 701.400 369.600 702.600 382.050 ;
        RECT 734.400 369.600 735.600 382.050 ;
        RECT 698.550 363.750 700.350 369.600 ;
        RECT 701.550 363.750 703.350 369.600 ;
        RECT 731.550 363.750 733.350 369.600 ;
        RECT 734.550 363.750 736.350 369.600 ;
        RECT 26.550 347.400 28.350 359.250 ;
        RECT 29.550 346.500 31.350 359.250 ;
        RECT 32.550 347.400 34.350 359.250 ;
        RECT 35.550 346.500 37.350 359.250 ;
        RECT 38.550 347.400 40.350 359.250 ;
        RECT 41.550 346.500 43.350 359.250 ;
        RECT 44.550 347.400 46.350 359.250 ;
        RECT 47.550 346.500 49.350 359.250 ;
        RECT 50.550 347.400 52.350 359.250 ;
        RECT 84.300 347.400 86.100 359.250 ;
        RECT 88.500 347.400 90.300 359.250 ;
        RECT 91.800 353.400 93.600 359.250 ;
        RECT 99.150 347.400 100.950 359.250 ;
        RECT 102.150 353.400 103.950 359.250 ;
        RECT 107.250 353.400 109.050 359.250 ;
        RECT 112.050 353.400 113.850 359.250 ;
        RECT 107.550 352.500 108.750 353.400 ;
        RECT 115.050 352.500 116.850 359.250 ;
        RECT 118.950 353.400 120.750 359.250 ;
        RECT 123.150 353.400 124.950 359.250 ;
        RECT 127.650 356.400 129.450 359.250 ;
        RECT 103.950 350.400 108.750 352.500 ;
        RECT 111.150 350.700 118.050 352.500 ;
        RECT 123.150 351.300 127.050 353.400 ;
        RECT 107.550 349.500 108.750 350.400 ;
        RECT 120.450 349.800 122.250 350.400 ;
        RECT 107.550 348.300 115.050 349.500 ;
        RECT 113.250 347.700 115.050 348.300 ;
        RECT 115.950 348.900 122.250 349.800 ;
        RECT 29.550 345.300 33.450 346.500 ;
        RECT 35.550 345.300 39.300 346.500 ;
        RECT 41.550 345.300 45.300 346.500 ;
        RECT 47.550 345.300 50.250 346.500 ;
        RECT 28.950 338.850 31.050 340.950 ;
        RECT 29.100 337.050 30.900 338.850 ;
        RECT 32.250 338.400 33.450 345.300 ;
        RECT 38.100 338.400 39.300 345.300 ;
        RECT 44.100 338.400 45.300 345.300 ;
        RECT 49.200 340.950 50.250 345.300 ;
        RECT 83.100 342.150 84.900 343.950 ;
        RECT 88.950 342.150 90.150 347.400 ;
        RECT 91.950 345.150 93.750 346.950 ;
        RECT 99.150 346.800 110.250 347.400 ;
        RECT 115.950 346.800 116.850 348.900 ;
        RECT 120.450 348.600 122.250 348.900 ;
        RECT 123.150 348.600 125.850 350.400 ;
        RECT 123.150 347.700 124.050 348.600 ;
        RECT 99.150 346.200 116.850 346.800 ;
        RECT 91.950 343.050 94.050 345.150 ;
        RECT 49.200 338.850 52.050 340.950 ;
        RECT 82.950 340.050 85.050 342.150 ;
        RECT 85.950 338.850 88.050 340.950 ;
        RECT 88.950 340.050 91.050 342.150 ;
        RECT 32.250 336.600 36.300 338.400 ;
        RECT 38.100 336.600 42.300 338.400 ;
        RECT 44.100 336.600 48.300 338.400 ;
        RECT 32.250 335.700 33.450 336.600 ;
        RECT 38.100 335.700 39.300 336.600 ;
        RECT 44.100 335.700 45.300 336.600 ;
        RECT 49.200 335.700 50.250 338.850 ;
        RECT 86.100 337.050 87.900 338.850 ;
        RECT 89.850 336.750 91.050 340.050 ;
        RECT 90.000 335.700 93.750 336.750 ;
        RECT 29.400 334.500 33.450 335.700 ;
        RECT 35.550 334.500 39.300 335.700 ;
        RECT 41.400 334.500 45.300 335.700 ;
        RECT 47.400 334.650 50.250 335.700 ;
        RECT 47.400 334.500 50.100 334.650 ;
        RECT 29.400 333.600 31.200 334.500 ;
        RECT 26.550 327.750 28.350 333.600 ;
        RECT 29.550 327.750 31.350 333.600 ;
        RECT 32.550 327.750 34.350 333.600 ;
        RECT 35.550 327.750 37.350 334.500 ;
        RECT 41.400 333.600 43.200 334.500 ;
        RECT 47.400 333.600 49.200 334.500 ;
        RECT 38.550 327.750 40.350 333.600 ;
        RECT 41.550 327.750 43.350 333.600 ;
        RECT 44.550 327.750 46.350 333.600 ;
        RECT 47.550 327.750 49.350 333.600 ;
        RECT 50.550 327.750 52.350 333.600 ;
        RECT 83.550 332.700 91.350 334.050 ;
        RECT 83.550 327.750 85.350 332.700 ;
        RECT 86.550 327.750 88.350 331.800 ;
        RECT 89.550 327.750 91.350 332.700 ;
        RECT 92.550 333.600 93.750 335.700 ;
        RECT 99.150 333.600 100.050 346.200 ;
        RECT 108.450 345.900 116.850 346.200 ;
        RECT 118.050 346.800 124.050 347.700 ;
        RECT 124.950 346.800 127.050 347.700 ;
        RECT 130.650 347.400 132.450 359.250 ;
        RECT 158.550 353.400 160.350 359.250 ;
        RECT 161.550 353.400 163.350 359.250 ;
        RECT 108.450 345.600 110.250 345.900 ;
        RECT 118.050 342.150 118.950 346.800 ;
        RECT 124.950 345.600 129.150 346.800 ;
        RECT 128.250 343.800 130.050 345.600 ;
        RECT 109.950 341.100 112.050 342.150 ;
        RECT 101.100 339.150 102.900 340.950 ;
        RECT 104.100 340.050 112.050 341.100 ;
        RECT 115.950 340.050 118.950 342.150 ;
        RECT 104.100 339.300 105.900 340.050 ;
        RECT 102.000 338.400 102.900 339.150 ;
        RECT 107.100 338.400 108.900 339.000 ;
        RECT 102.000 337.200 108.900 338.400 ;
        RECT 107.850 336.000 108.900 337.200 ;
        RECT 118.050 336.000 118.950 340.050 ;
        RECT 127.950 339.750 130.050 340.050 ;
        RECT 126.150 337.950 130.050 339.750 ;
        RECT 131.250 337.950 132.450 347.400 ;
        RECT 161.400 340.950 162.600 353.400 ;
        RECT 195.300 347.400 197.100 359.250 ;
        RECT 199.500 347.400 201.300 359.250 ;
        RECT 202.800 353.400 204.600 359.250 ;
        RECT 239.400 353.400 241.200 359.250 ;
        RECT 242.700 347.400 244.500 359.250 ;
        RECT 246.900 347.400 248.700 359.250 ;
        RECT 279.300 347.400 281.100 359.250 ;
        RECT 283.500 347.400 285.300 359.250 ;
        RECT 286.800 353.400 288.600 359.250 ;
        RECT 320.400 353.400 322.200 359.250 ;
        RECT 323.700 347.400 325.500 359.250 ;
        RECT 327.900 347.400 329.700 359.250 ;
        RECT 332.550 347.400 334.350 359.250 ;
        RECT 335.550 356.400 337.350 359.250 ;
        RECT 340.050 353.400 341.850 359.250 ;
        RECT 344.250 353.400 346.050 359.250 ;
        RECT 337.950 351.300 341.850 353.400 ;
        RECT 348.150 352.500 349.950 359.250 ;
        RECT 351.150 353.400 352.950 359.250 ;
        RECT 355.950 353.400 357.750 359.250 ;
        RECT 361.050 353.400 362.850 359.250 ;
        RECT 356.250 352.500 357.450 353.400 ;
        RECT 346.950 350.700 353.850 352.500 ;
        RECT 356.250 350.400 361.050 352.500 ;
        RECT 339.150 348.600 341.850 350.400 ;
        RECT 342.750 349.800 344.550 350.400 ;
        RECT 342.750 348.900 349.050 349.800 ;
        RECT 356.250 349.500 357.450 350.400 ;
        RECT 342.750 348.600 344.550 348.900 ;
        RECT 340.950 347.700 341.850 348.600 ;
        RECT 194.100 342.150 195.900 343.950 ;
        RECT 199.950 342.150 201.150 347.400 ;
        RECT 202.950 345.150 204.750 346.950 ;
        RECT 239.250 345.150 241.050 346.950 ;
        RECT 202.950 343.050 205.050 345.150 ;
        RECT 238.950 343.050 241.050 345.150 ;
        RECT 242.850 342.150 244.050 347.400 ;
        RECT 248.100 342.150 249.900 343.950 ;
        RECT 278.100 342.150 279.900 343.950 ;
        RECT 283.950 342.150 285.150 347.400 ;
        RECT 286.950 345.150 288.750 346.950 ;
        RECT 320.250 345.150 322.050 346.950 ;
        RECT 286.950 343.050 289.050 345.150 ;
        RECT 319.950 343.050 322.050 345.150 ;
        RECT 323.850 342.150 325.050 347.400 ;
        RECT 329.100 342.150 330.900 343.950 ;
        RECT 158.100 339.150 159.900 340.950 ;
        RECT 107.850 335.100 118.950 336.000 ;
        RECT 127.950 335.850 132.450 337.950 ;
        RECT 157.950 337.050 160.050 339.150 ;
        RECT 160.950 338.850 163.050 340.950 ;
        RECT 193.950 340.050 196.050 342.150 ;
        RECT 196.950 338.850 199.050 340.950 ;
        RECT 199.950 340.050 202.050 342.150 ;
        RECT 107.850 334.200 108.900 335.100 ;
        RECT 118.050 334.800 118.950 335.100 ;
        RECT 92.550 327.750 94.350 333.600 ;
        RECT 99.150 327.750 100.950 333.600 ;
        RECT 103.950 331.500 106.050 333.600 ;
        RECT 107.550 332.400 109.350 334.200 ;
        RECT 110.850 333.450 112.650 334.200 ;
        RECT 110.850 332.400 115.800 333.450 ;
        RECT 118.050 333.000 119.850 334.800 ;
        RECT 131.250 333.600 132.450 335.850 ;
        RECT 124.950 332.700 127.050 333.600 ;
        RECT 105.000 330.600 106.050 331.500 ;
        RECT 114.750 330.600 115.800 332.400 ;
        RECT 123.300 331.500 127.050 332.700 ;
        RECT 123.300 330.600 124.350 331.500 ;
        RECT 102.150 327.750 103.950 330.600 ;
        RECT 105.000 329.700 108.750 330.600 ;
        RECT 106.950 327.750 108.750 329.700 ;
        RECT 111.450 327.750 113.250 330.600 ;
        RECT 114.750 327.750 116.550 330.600 ;
        RECT 118.650 327.750 120.450 330.600 ;
        RECT 122.850 327.750 124.650 330.600 ;
        RECT 127.350 327.750 129.150 330.600 ;
        RECT 130.650 327.750 132.450 333.600 ;
        RECT 161.400 330.600 162.600 338.850 ;
        RECT 197.100 337.050 198.900 338.850 ;
        RECT 200.850 336.750 202.050 340.050 ;
        RECT 241.950 340.050 244.050 342.150 ;
        RECT 241.950 336.750 243.150 340.050 ;
        RECT 244.950 338.850 247.050 340.950 ;
        RECT 247.950 340.050 250.050 342.150 ;
        RECT 277.950 340.050 280.050 342.150 ;
        RECT 280.950 338.850 283.050 340.950 ;
        RECT 283.950 340.050 286.050 342.150 ;
        RECT 245.100 337.050 246.900 338.850 ;
        RECT 281.100 337.050 282.900 338.850 ;
        RECT 284.850 336.750 286.050 340.050 ;
        RECT 322.950 340.050 325.050 342.150 ;
        RECT 322.950 336.750 324.150 340.050 ;
        RECT 325.950 338.850 328.050 340.950 ;
        RECT 328.950 340.050 331.050 342.150 ;
        RECT 326.100 337.050 327.900 338.850 ;
        RECT 332.550 337.950 333.750 347.400 ;
        RECT 337.950 346.800 340.050 347.700 ;
        RECT 340.950 346.800 346.950 347.700 ;
        RECT 335.850 345.600 340.050 346.800 ;
        RECT 334.950 343.800 336.750 345.600 ;
        RECT 346.050 342.150 346.950 346.800 ;
        RECT 348.150 346.800 349.050 348.900 ;
        RECT 349.950 348.300 357.450 349.500 ;
        RECT 349.950 347.700 351.750 348.300 ;
        RECT 364.050 347.400 365.850 359.250 ;
        RECT 397.050 347.400 398.850 359.250 ;
        RECT 400.050 347.400 401.850 359.250 ;
        RECT 403.650 353.400 405.450 359.250 ;
        RECT 406.650 353.400 408.450 359.250 ;
        RECT 440.400 353.400 442.200 359.250 ;
        RECT 354.750 346.800 365.850 347.400 ;
        RECT 348.150 346.200 365.850 346.800 ;
        RECT 348.150 345.900 356.550 346.200 ;
        RECT 354.750 345.600 356.550 345.900 ;
        RECT 346.050 340.050 349.050 342.150 ;
        RECT 352.950 341.100 355.050 342.150 ;
        RECT 352.950 340.050 360.900 341.100 ;
        RECT 334.950 339.750 337.050 340.050 ;
        RECT 334.950 337.950 338.850 339.750 ;
        RECT 201.000 335.700 204.750 336.750 ;
        RECT 194.550 332.700 202.350 334.050 ;
        RECT 158.550 327.750 160.350 330.600 ;
        RECT 161.550 327.750 163.350 330.600 ;
        RECT 194.550 327.750 196.350 332.700 ;
        RECT 197.550 327.750 199.350 331.800 ;
        RECT 200.550 327.750 202.350 332.700 ;
        RECT 203.550 333.600 204.750 335.700 ;
        RECT 239.250 335.700 243.000 336.750 ;
        RECT 285.000 335.700 288.750 336.750 ;
        RECT 239.250 333.600 240.450 335.700 ;
        RECT 203.550 327.750 205.350 333.600 ;
        RECT 238.650 327.750 240.450 333.600 ;
        RECT 241.650 332.700 249.450 334.050 ;
        RECT 241.650 327.750 243.450 332.700 ;
        RECT 244.650 327.750 246.450 331.800 ;
        RECT 247.650 327.750 249.450 332.700 ;
        RECT 278.550 332.700 286.350 334.050 ;
        RECT 278.550 327.750 280.350 332.700 ;
        RECT 281.550 327.750 283.350 331.800 ;
        RECT 284.550 327.750 286.350 332.700 ;
        RECT 287.550 333.600 288.750 335.700 ;
        RECT 320.250 335.700 324.000 336.750 ;
        RECT 332.550 335.850 337.050 337.950 ;
        RECT 346.050 336.000 346.950 340.050 ;
        RECT 359.100 339.300 360.900 340.050 ;
        RECT 362.100 339.150 363.900 340.950 ;
        RECT 356.100 338.400 357.900 339.000 ;
        RECT 362.100 338.400 363.000 339.150 ;
        RECT 356.100 337.200 363.000 338.400 ;
        RECT 356.100 336.000 357.150 337.200 ;
        RECT 320.250 333.600 321.450 335.700 ;
        RECT 287.550 327.750 289.350 333.600 ;
        RECT 319.650 327.750 321.450 333.600 ;
        RECT 322.650 332.700 330.450 334.050 ;
        RECT 322.650 327.750 324.450 332.700 ;
        RECT 325.650 327.750 327.450 331.800 ;
        RECT 328.650 327.750 330.450 332.700 ;
        RECT 332.550 333.600 333.750 335.850 ;
        RECT 346.050 335.100 357.150 336.000 ;
        RECT 346.050 334.800 346.950 335.100 ;
        RECT 332.550 327.750 334.350 333.600 ;
        RECT 337.950 332.700 340.050 333.600 ;
        RECT 345.150 333.000 346.950 334.800 ;
        RECT 356.100 334.200 357.150 335.100 ;
        RECT 352.350 333.450 354.150 334.200 ;
        RECT 337.950 331.500 341.700 332.700 ;
        RECT 340.650 330.600 341.700 331.500 ;
        RECT 349.200 332.400 354.150 333.450 ;
        RECT 355.650 332.400 357.450 334.200 ;
        RECT 364.950 333.600 365.850 346.200 ;
        RECT 349.200 330.600 350.250 332.400 ;
        RECT 358.950 331.500 361.050 333.600 ;
        RECT 358.950 330.600 360.000 331.500 ;
        RECT 335.850 327.750 337.650 330.600 ;
        RECT 340.350 327.750 342.150 330.600 ;
        RECT 344.550 327.750 346.350 330.600 ;
        RECT 348.450 327.750 350.250 330.600 ;
        RECT 351.750 327.750 353.550 330.600 ;
        RECT 356.250 329.700 360.000 330.600 ;
        RECT 356.250 327.750 358.050 329.700 ;
        RECT 361.050 327.750 362.850 330.600 ;
        RECT 364.050 327.750 365.850 333.600 ;
        RECT 397.650 342.150 398.850 347.400 ;
        RECT 397.650 340.050 400.050 342.150 ;
        RECT 400.950 341.850 403.050 343.950 ;
        RECT 401.100 340.050 402.900 341.850 ;
        RECT 397.650 333.600 398.850 340.050 ;
        RECT 404.100 336.300 405.300 353.400 ;
        RECT 443.700 347.400 445.500 359.250 ;
        RECT 447.900 347.400 449.700 359.250 ;
        RECT 480.300 347.400 482.100 359.250 ;
        RECT 484.500 347.400 486.300 359.250 ;
        RECT 487.800 353.400 489.600 359.250 ;
        RECT 521.550 353.400 523.350 359.250 ;
        RECT 440.250 345.150 442.050 346.950 ;
        RECT 407.100 342.150 408.900 343.950 ;
        RECT 439.950 343.050 442.050 345.150 ;
        RECT 443.850 342.150 445.050 347.400 ;
        RECT 449.100 342.150 450.900 343.950 ;
        RECT 479.100 342.150 480.900 343.950 ;
        RECT 484.950 342.150 486.150 347.400 ;
        RECT 487.950 345.150 489.750 346.950 ;
        RECT 521.550 346.500 522.750 353.400 ;
        RECT 524.850 347.400 526.650 359.250 ;
        RECT 527.850 347.400 529.650 359.250 ;
        RECT 533.550 347.400 535.350 359.250 ;
        RECT 536.550 356.400 538.350 359.250 ;
        RECT 541.050 353.400 542.850 359.250 ;
        RECT 545.250 353.400 547.050 359.250 ;
        RECT 538.950 351.300 542.850 353.400 ;
        RECT 549.150 352.500 550.950 359.250 ;
        RECT 552.150 353.400 553.950 359.250 ;
        RECT 556.950 353.400 558.750 359.250 ;
        RECT 562.050 353.400 563.850 359.250 ;
        RECT 557.250 352.500 558.450 353.400 ;
        RECT 547.950 350.700 554.850 352.500 ;
        RECT 557.250 350.400 562.050 352.500 ;
        RECT 540.150 348.600 542.850 350.400 ;
        RECT 543.750 349.800 545.550 350.400 ;
        RECT 543.750 348.900 550.050 349.800 ;
        RECT 557.250 349.500 558.450 350.400 ;
        RECT 543.750 348.600 545.550 348.900 ;
        RECT 541.950 347.700 542.850 348.600 ;
        RECT 521.550 345.600 527.250 346.500 ;
        RECT 487.950 343.050 490.050 345.150 ;
        RECT 525.000 344.700 527.250 345.600 ;
        RECT 521.100 342.150 522.900 343.950 ;
        RECT 406.950 340.050 409.050 342.150 ;
        RECT 442.950 340.050 445.050 342.150 ;
        RECT 442.950 336.750 444.150 340.050 ;
        RECT 445.950 338.850 448.050 340.950 ;
        RECT 448.950 340.050 451.050 342.150 ;
        RECT 478.950 340.050 481.050 342.150 ;
        RECT 481.950 338.850 484.050 340.950 ;
        RECT 484.950 340.050 487.050 342.150 ;
        RECT 520.950 340.050 523.050 342.150 ;
        RECT 446.100 337.050 447.900 338.850 ;
        RECT 482.100 337.050 483.900 338.850 ;
        RECT 485.850 336.750 487.050 340.050 ;
        RECT 400.950 335.100 408.450 336.300 ;
        RECT 400.950 334.500 402.750 335.100 ;
        RECT 397.650 332.100 400.950 333.600 ;
        RECT 399.150 327.750 400.950 332.100 ;
        RECT 402.150 327.750 403.950 333.600 ;
        RECT 406.650 327.750 408.450 335.100 ;
        RECT 440.250 335.700 444.000 336.750 ;
        RECT 486.000 335.700 489.750 336.750 ;
        RECT 440.250 333.600 441.450 335.700 ;
        RECT 439.650 327.750 441.450 333.600 ;
        RECT 442.650 332.700 450.450 334.050 ;
        RECT 442.650 327.750 444.450 332.700 ;
        RECT 445.650 327.750 447.450 331.800 ;
        RECT 448.650 327.750 450.450 332.700 ;
        RECT 479.550 332.700 487.350 334.050 ;
        RECT 479.550 327.750 481.350 332.700 ;
        RECT 482.550 327.750 484.350 331.800 ;
        RECT 485.550 327.750 487.350 332.700 ;
        RECT 488.550 333.600 489.750 335.700 ;
        RECT 525.000 336.300 526.050 344.700 ;
        RECT 528.150 342.150 529.350 347.400 ;
        RECT 526.950 340.050 529.350 342.150 ;
        RECT 525.000 335.400 527.250 336.300 ;
        RECT 522.150 334.500 527.250 335.400 ;
        RECT 488.550 327.750 490.350 333.600 ;
        RECT 522.150 330.600 523.350 334.500 ;
        RECT 528.150 333.600 529.350 340.050 ;
        RECT 533.550 337.950 534.750 347.400 ;
        RECT 538.950 346.800 541.050 347.700 ;
        RECT 541.950 346.800 547.950 347.700 ;
        RECT 536.850 345.600 541.050 346.800 ;
        RECT 535.950 343.800 537.750 345.600 ;
        RECT 547.050 342.150 547.950 346.800 ;
        RECT 549.150 346.800 550.050 348.900 ;
        RECT 550.950 348.300 558.450 349.500 ;
        RECT 550.950 347.700 552.750 348.300 ;
        RECT 565.050 347.400 566.850 359.250 ;
        RECT 599.400 353.400 601.200 359.250 ;
        RECT 602.700 347.400 604.500 359.250 ;
        RECT 606.900 347.400 608.700 359.250 ;
        RECT 642.450 347.400 644.250 359.250 ;
        RECT 646.650 347.400 648.450 359.250 ;
        RECT 676.650 353.400 678.450 359.250 ;
        RECT 679.650 353.400 681.450 359.250 ;
        RECT 682.650 353.400 684.450 359.250 ;
        RECT 555.750 346.800 566.850 347.400 ;
        RECT 549.150 346.200 566.850 346.800 ;
        RECT 549.150 345.900 557.550 346.200 ;
        RECT 555.750 345.600 557.550 345.900 ;
        RECT 547.050 340.050 550.050 342.150 ;
        RECT 553.950 341.100 556.050 342.150 ;
        RECT 553.950 340.050 561.900 341.100 ;
        RECT 535.950 339.750 538.050 340.050 ;
        RECT 535.950 337.950 539.850 339.750 ;
        RECT 533.550 335.850 538.050 337.950 ;
        RECT 547.050 336.000 547.950 340.050 ;
        RECT 560.100 339.300 561.900 340.050 ;
        RECT 563.100 339.150 564.900 340.950 ;
        RECT 557.100 338.400 558.900 339.000 ;
        RECT 563.100 338.400 564.000 339.150 ;
        RECT 557.100 337.200 564.000 338.400 ;
        RECT 557.100 336.000 558.150 337.200 ;
        RECT 533.550 333.600 534.750 335.850 ;
        RECT 547.050 335.100 558.150 336.000 ;
        RECT 547.050 334.800 547.950 335.100 ;
        RECT 521.550 327.750 523.350 330.600 ;
        RECT 524.850 327.750 526.650 333.600 ;
        RECT 527.850 327.750 529.650 333.600 ;
        RECT 533.550 327.750 535.350 333.600 ;
        RECT 538.950 332.700 541.050 333.600 ;
        RECT 546.150 333.000 547.950 334.800 ;
        RECT 557.100 334.200 558.150 335.100 ;
        RECT 553.350 333.450 555.150 334.200 ;
        RECT 538.950 331.500 542.700 332.700 ;
        RECT 541.650 330.600 542.700 331.500 ;
        RECT 550.200 332.400 555.150 333.450 ;
        RECT 556.650 332.400 558.450 334.200 ;
        RECT 565.950 333.600 566.850 346.200 ;
        RECT 599.250 345.150 601.050 346.950 ;
        RECT 598.950 343.050 601.050 345.150 ;
        RECT 602.850 342.150 604.050 347.400 ;
        RECT 642.450 346.350 645.000 347.400 ;
        RECT 608.100 342.150 609.900 343.950 ;
        RECT 641.100 342.150 642.900 343.950 ;
        RECT 601.950 340.050 604.050 342.150 ;
        RECT 601.950 336.750 603.150 340.050 ;
        RECT 604.950 338.850 607.050 340.950 ;
        RECT 607.950 340.050 610.050 342.150 ;
        RECT 640.950 340.050 643.050 342.150 ;
        RECT 643.950 339.150 645.000 346.350 ;
        RECT 680.250 345.150 681.450 353.400 ;
        RECT 713.550 348.300 715.350 359.250 ;
        RECT 716.550 349.200 718.350 359.250 ;
        RECT 719.550 348.300 721.350 359.250 ;
        RECT 713.550 347.400 721.350 348.300 ;
        RECT 722.550 347.400 724.350 359.250 ;
        RECT 757.650 353.400 759.450 359.250 ;
        RECT 760.650 353.400 762.450 359.250 ;
        RECT 647.100 342.150 648.900 343.950 ;
        RECT 646.950 340.050 649.050 342.150 ;
        RECT 676.950 341.850 679.050 343.950 ;
        RECT 679.950 343.050 682.050 345.150 ;
        RECT 677.100 340.050 678.900 341.850 ;
        RECT 605.100 337.050 606.900 338.850 ;
        RECT 643.950 337.050 646.050 339.150 ;
        RECT 599.250 335.700 603.000 336.750 ;
        RECT 599.250 333.600 600.450 335.700 ;
        RECT 550.200 330.600 551.250 332.400 ;
        RECT 559.950 331.500 562.050 333.600 ;
        RECT 559.950 330.600 561.000 331.500 ;
        RECT 536.850 327.750 538.650 330.600 ;
        RECT 541.350 327.750 543.150 330.600 ;
        RECT 545.550 327.750 547.350 330.600 ;
        RECT 549.450 327.750 551.250 330.600 ;
        RECT 552.750 327.750 554.550 330.600 ;
        RECT 557.250 329.700 561.000 330.600 ;
        RECT 557.250 327.750 559.050 329.700 ;
        RECT 562.050 327.750 563.850 330.600 ;
        RECT 565.050 327.750 566.850 333.600 ;
        RECT 598.650 327.750 600.450 333.600 ;
        RECT 601.650 332.700 609.450 334.050 ;
        RECT 601.650 327.750 603.450 332.700 ;
        RECT 604.650 327.750 606.450 331.800 ;
        RECT 607.650 327.750 609.450 332.700 ;
        RECT 643.950 330.600 645.000 337.050 ;
        RECT 680.250 335.700 681.450 343.050 ;
        RECT 682.950 341.850 685.050 343.950 ;
        RECT 722.700 342.150 723.900 347.400 ;
        RECT 683.100 340.050 684.900 341.850 ;
        RECT 712.950 338.850 715.050 340.950 ;
        RECT 716.100 339.150 717.900 340.950 ;
        RECT 713.100 337.050 714.900 338.850 ;
        RECT 715.950 337.050 718.050 339.150 ;
        RECT 718.950 338.850 721.050 340.950 ;
        RECT 721.950 340.050 724.050 342.150 ;
        RECT 758.400 340.950 759.600 353.400 ;
        RECT 719.100 337.050 720.900 338.850 ;
        RECT 677.850 334.800 681.450 335.700 ;
        RECT 640.650 327.750 642.450 330.600 ;
        RECT 643.650 327.750 645.450 330.600 ;
        RECT 646.650 327.750 648.450 330.600 ;
        RECT 677.850 327.750 679.650 334.800 ;
        RECT 722.700 333.600 723.900 340.050 ;
        RECT 757.950 338.850 760.050 340.950 ;
        RECT 761.100 339.150 762.900 340.950 ;
        RECT 682.350 327.750 684.150 333.600 ;
        RECT 714.000 327.750 715.800 333.600 ;
        RECT 718.200 331.950 723.900 333.600 ;
        RECT 718.200 327.750 720.000 331.950 ;
        RECT 758.400 330.600 759.600 338.850 ;
        RECT 760.950 337.050 763.050 339.150 ;
        RECT 721.500 327.750 723.300 330.600 ;
        RECT 757.650 327.750 759.450 330.600 ;
        RECT 760.650 327.750 762.450 330.600 ;
        RECT 3.150 317.400 4.950 323.250 ;
        RECT 6.150 320.400 7.950 323.250 ;
        RECT 10.950 321.300 12.750 323.250 ;
        RECT 9.000 320.400 12.750 321.300 ;
        RECT 15.450 320.400 17.250 323.250 ;
        RECT 18.750 320.400 20.550 323.250 ;
        RECT 22.650 320.400 24.450 323.250 ;
        RECT 26.850 320.400 28.650 323.250 ;
        RECT 31.350 320.400 33.150 323.250 ;
        RECT 9.000 319.500 10.050 320.400 ;
        RECT 7.950 317.400 10.050 319.500 ;
        RECT 18.750 318.600 19.800 320.400 ;
        RECT 3.150 304.800 4.050 317.400 ;
        RECT 11.550 316.800 13.350 318.600 ;
        RECT 14.850 317.550 19.800 318.600 ;
        RECT 27.300 319.500 28.350 320.400 ;
        RECT 27.300 318.300 31.050 319.500 ;
        RECT 14.850 316.800 16.650 317.550 ;
        RECT 11.850 315.900 12.900 316.800 ;
        RECT 22.050 316.200 23.850 318.000 ;
        RECT 28.950 317.400 31.050 318.300 ;
        RECT 34.650 317.400 36.450 323.250 ;
        RECT 22.050 315.900 22.950 316.200 ;
        RECT 11.850 315.000 22.950 315.900 ;
        RECT 35.250 315.150 36.450 317.400 ;
        RECT 11.850 313.800 12.900 315.000 ;
        RECT 6.000 312.600 12.900 313.800 ;
        RECT 6.000 311.850 6.900 312.600 ;
        RECT 11.100 312.000 12.900 312.600 ;
        RECT 5.100 310.050 6.900 311.850 ;
        RECT 8.100 310.950 9.900 311.700 ;
        RECT 22.050 310.950 22.950 315.000 ;
        RECT 31.950 313.050 36.450 315.150 ;
        RECT 30.150 311.250 34.050 313.050 ;
        RECT 31.950 310.950 34.050 311.250 ;
        RECT 8.100 309.900 16.050 310.950 ;
        RECT 13.950 308.850 16.050 309.900 ;
        RECT 19.950 308.850 22.950 310.950 ;
        RECT 12.450 305.100 14.250 305.400 ;
        RECT 12.450 304.800 20.850 305.100 ;
        RECT 3.150 304.200 20.850 304.800 ;
        RECT 3.150 303.600 14.250 304.200 ;
        RECT 3.150 291.750 4.950 303.600 ;
        RECT 17.250 302.700 19.050 303.300 ;
        RECT 11.550 301.500 19.050 302.700 ;
        RECT 19.950 302.100 20.850 304.200 ;
        RECT 22.050 304.200 22.950 308.850 ;
        RECT 32.250 305.400 34.050 307.200 ;
        RECT 28.950 304.200 33.150 305.400 ;
        RECT 22.050 303.300 28.050 304.200 ;
        RECT 28.950 303.300 31.050 304.200 ;
        RECT 35.250 303.600 36.450 313.050 ;
        RECT 27.150 302.400 28.050 303.300 ;
        RECT 24.450 302.100 26.250 302.400 ;
        RECT 11.550 300.600 12.750 301.500 ;
        RECT 19.950 301.200 26.250 302.100 ;
        RECT 24.450 300.600 26.250 301.200 ;
        RECT 27.150 300.600 29.850 302.400 ;
        RECT 7.950 298.500 12.750 300.600 ;
        RECT 15.150 298.500 22.050 300.300 ;
        RECT 11.550 297.600 12.750 298.500 ;
        RECT 6.150 291.750 7.950 297.600 ;
        RECT 11.250 291.750 13.050 297.600 ;
        RECT 16.050 291.750 17.850 297.600 ;
        RECT 19.050 291.750 20.850 298.500 ;
        RECT 27.150 297.600 31.050 299.700 ;
        RECT 22.950 291.750 24.750 297.600 ;
        RECT 27.150 291.750 28.950 297.600 ;
        RECT 31.650 291.750 33.450 294.600 ;
        RECT 34.650 291.750 36.450 303.600 ;
        RECT 38.550 317.400 40.350 323.250 ;
        RECT 41.850 320.400 43.650 323.250 ;
        RECT 46.350 320.400 48.150 323.250 ;
        RECT 50.550 320.400 52.350 323.250 ;
        RECT 54.450 320.400 56.250 323.250 ;
        RECT 57.750 320.400 59.550 323.250 ;
        RECT 62.250 321.300 64.050 323.250 ;
        RECT 62.250 320.400 66.000 321.300 ;
        RECT 67.050 320.400 68.850 323.250 ;
        RECT 46.650 319.500 47.700 320.400 ;
        RECT 43.950 318.300 47.700 319.500 ;
        RECT 55.200 318.600 56.250 320.400 ;
        RECT 64.950 319.500 66.000 320.400 ;
        RECT 43.950 317.400 46.050 318.300 ;
        RECT 38.550 315.150 39.750 317.400 ;
        RECT 51.150 316.200 52.950 318.000 ;
        RECT 55.200 317.550 60.150 318.600 ;
        RECT 58.350 316.800 60.150 317.550 ;
        RECT 61.650 316.800 63.450 318.600 ;
        RECT 64.950 317.400 67.050 319.500 ;
        RECT 70.050 317.400 71.850 323.250 ;
        RECT 104.700 320.400 106.500 323.250 ;
        RECT 108.000 319.050 109.800 323.250 ;
        RECT 52.050 315.900 52.950 316.200 ;
        RECT 62.100 315.900 63.150 316.800 ;
        RECT 38.550 313.050 43.050 315.150 ;
        RECT 52.050 315.000 63.150 315.900 ;
        RECT 38.550 303.600 39.750 313.050 ;
        RECT 40.950 311.250 44.850 313.050 ;
        RECT 40.950 310.950 43.050 311.250 ;
        RECT 52.050 310.950 52.950 315.000 ;
        RECT 62.100 313.800 63.150 315.000 ;
        RECT 62.100 312.600 69.000 313.800 ;
        RECT 62.100 312.000 63.900 312.600 ;
        RECT 68.100 311.850 69.000 312.600 ;
        RECT 65.100 310.950 66.900 311.700 ;
        RECT 52.050 308.850 55.050 310.950 ;
        RECT 58.950 309.900 66.900 310.950 ;
        RECT 68.100 310.050 69.900 311.850 ;
        RECT 58.950 308.850 61.050 309.900 ;
        RECT 40.950 305.400 42.750 307.200 ;
        RECT 41.850 304.200 46.050 305.400 ;
        RECT 52.050 304.200 52.950 308.850 ;
        RECT 60.750 305.100 62.550 305.400 ;
        RECT 38.550 291.750 40.350 303.600 ;
        RECT 43.950 303.300 46.050 304.200 ;
        RECT 46.950 303.300 52.950 304.200 ;
        RECT 54.150 304.800 62.550 305.100 ;
        RECT 70.950 304.800 71.850 317.400 ;
        RECT 104.100 317.400 109.800 319.050 ;
        RECT 112.200 317.400 114.000 323.250 ;
        RECT 145.350 317.400 147.150 323.250 ;
        RECT 148.350 317.400 150.150 323.250 ;
        RECT 151.650 320.400 153.450 323.250 ;
        RECT 185.700 320.400 187.500 323.250 ;
        RECT 104.100 310.950 105.300 317.400 ;
        RECT 107.100 312.150 108.900 313.950 ;
        RECT 103.950 308.850 106.050 310.950 ;
        RECT 106.950 310.050 109.050 312.150 ;
        RECT 109.950 311.850 112.050 313.950 ;
        RECT 113.100 312.150 114.900 313.950 ;
        RECT 110.100 310.050 111.900 311.850 ;
        RECT 112.950 310.050 115.050 312.150 ;
        RECT 145.650 310.950 146.850 317.400 ;
        RECT 151.650 316.500 152.850 320.400 ;
        RECT 189.000 319.050 190.800 323.250 ;
        RECT 147.750 315.600 152.850 316.500 ;
        RECT 185.100 317.400 190.800 319.050 ;
        RECT 193.200 317.400 195.000 323.250 ;
        RECT 226.650 317.400 228.450 323.250 ;
        RECT 147.750 314.700 150.000 315.600 ;
        RECT 145.650 308.850 148.050 310.950 ;
        RECT 54.150 304.200 71.850 304.800 ;
        RECT 46.950 302.400 47.850 303.300 ;
        RECT 45.150 300.600 47.850 302.400 ;
        RECT 48.750 302.100 50.550 302.400 ;
        RECT 54.150 302.100 55.050 304.200 ;
        RECT 60.750 303.600 71.850 304.200 ;
        RECT 104.100 303.600 105.300 308.850 ;
        RECT 145.650 303.600 146.850 308.850 ;
        RECT 148.950 306.300 150.000 314.700 ;
        RECT 185.100 310.950 186.300 317.400 ;
        RECT 227.250 315.300 228.450 317.400 ;
        RECT 229.650 318.300 231.450 323.250 ;
        RECT 232.650 319.200 234.450 323.250 ;
        RECT 235.650 318.300 237.450 323.250 ;
        RECT 263.550 320.400 265.350 323.250 ;
        RECT 266.550 320.400 268.350 323.250 ;
        RECT 299.550 320.400 301.350 323.250 ;
        RECT 229.650 316.950 237.450 318.300 ;
        RECT 227.250 314.250 231.000 315.300 ;
        RECT 188.100 312.150 189.900 313.950 ;
        RECT 151.950 308.850 154.050 310.950 ;
        RECT 184.950 308.850 187.050 310.950 ;
        RECT 187.950 310.050 190.050 312.150 ;
        RECT 190.950 311.850 193.050 313.950 ;
        RECT 194.100 312.150 195.900 313.950 ;
        RECT 191.100 310.050 192.900 311.850 ;
        RECT 193.950 310.050 196.050 312.150 ;
        RECT 229.950 310.950 231.150 314.250 ;
        RECT 233.100 312.150 234.900 313.950 ;
        RECT 229.950 308.850 232.050 310.950 ;
        RECT 232.950 310.050 235.050 312.150 ;
        RECT 262.950 311.850 265.050 313.950 ;
        RECT 266.400 312.150 267.600 320.400 ;
        RECT 300.150 316.500 301.350 320.400 ;
        RECT 302.850 317.400 304.650 323.250 ;
        RECT 305.850 317.400 307.650 323.250 ;
        RECT 338.550 320.400 340.350 323.250 ;
        RECT 341.550 320.400 343.350 323.250 ;
        RECT 300.150 315.600 305.250 316.500 ;
        RECT 303.000 314.700 305.250 315.600 ;
        RECT 235.950 308.850 238.050 310.950 ;
        RECT 263.100 310.050 264.900 311.850 ;
        RECT 265.950 310.050 268.050 312.150 ;
        RECT 152.100 307.050 153.900 308.850 ;
        RECT 147.750 305.400 150.000 306.300 ;
        RECT 147.750 304.500 153.450 305.400 ;
        RECT 48.750 301.200 55.050 302.100 ;
        RECT 55.950 302.700 57.750 303.300 ;
        RECT 55.950 301.500 63.450 302.700 ;
        RECT 48.750 300.600 50.550 301.200 ;
        RECT 62.250 300.600 63.450 301.500 ;
        RECT 43.950 297.600 47.850 299.700 ;
        RECT 52.950 298.500 59.850 300.300 ;
        RECT 62.250 298.500 67.050 300.600 ;
        RECT 41.550 291.750 43.350 294.600 ;
        RECT 46.050 291.750 47.850 297.600 ;
        RECT 50.250 291.750 52.050 297.600 ;
        RECT 54.150 291.750 55.950 298.500 ;
        RECT 62.250 297.600 63.450 298.500 ;
        RECT 57.150 291.750 58.950 297.600 ;
        RECT 61.950 291.750 63.750 297.600 ;
        RECT 67.050 291.750 68.850 297.600 ;
        RECT 70.050 291.750 71.850 303.600 ;
        RECT 103.650 291.750 105.450 303.600 ;
        RECT 106.650 302.700 114.450 303.600 ;
        RECT 106.650 291.750 108.450 302.700 ;
        RECT 109.650 291.750 111.450 301.800 ;
        RECT 112.650 291.750 114.450 302.700 ;
        RECT 145.350 291.750 147.150 303.600 ;
        RECT 148.350 291.750 150.150 303.600 ;
        RECT 152.250 297.600 153.450 304.500 ;
        RECT 185.100 303.600 186.300 308.850 ;
        RECT 226.950 305.850 229.050 307.950 ;
        RECT 227.250 304.050 229.050 305.850 ;
        RECT 230.850 303.600 232.050 308.850 ;
        RECT 236.100 307.050 237.900 308.850 ;
        RECT 151.650 291.750 153.450 297.600 ;
        RECT 184.650 291.750 186.450 303.600 ;
        RECT 187.650 302.700 195.450 303.600 ;
        RECT 187.650 291.750 189.450 302.700 ;
        RECT 190.650 291.750 192.450 301.800 ;
        RECT 193.650 291.750 195.450 302.700 ;
        RECT 227.400 291.750 229.200 297.600 ;
        RECT 230.700 291.750 232.500 303.600 ;
        RECT 234.900 291.750 236.700 303.600 ;
        RECT 266.400 297.600 267.600 310.050 ;
        RECT 298.950 308.850 301.050 310.950 ;
        RECT 299.100 307.050 300.900 308.850 ;
        RECT 303.000 306.300 304.050 314.700 ;
        RECT 306.150 310.950 307.350 317.400 ;
        RECT 337.950 311.850 340.050 313.950 ;
        RECT 341.400 312.150 342.600 320.400 ;
        RECT 374.550 318.300 376.350 323.250 ;
        RECT 377.550 319.200 379.350 323.250 ;
        RECT 380.550 318.300 382.350 323.250 ;
        RECT 374.550 316.950 382.350 318.300 ;
        RECT 383.550 317.400 385.350 323.250 ;
        RECT 415.650 317.400 417.450 323.250 ;
        RECT 383.550 315.300 384.750 317.400 ;
        RECT 381.000 314.250 384.750 315.300 ;
        RECT 416.250 315.300 417.450 317.400 ;
        RECT 418.650 318.300 420.450 323.250 ;
        RECT 421.650 319.200 423.450 323.250 ;
        RECT 424.650 318.300 426.450 323.250 ;
        RECT 418.650 316.950 426.450 318.300 ;
        RECT 452.850 317.400 454.650 323.250 ;
        RECT 457.350 316.200 459.150 323.250 ;
        RECT 491.550 320.400 493.350 323.250 ;
        RECT 455.550 315.300 459.150 316.200 ;
        RECT 492.150 316.500 493.350 320.400 ;
        RECT 494.850 317.400 496.650 323.250 ;
        RECT 497.850 317.400 499.650 323.250 ;
        RECT 534.150 318.900 535.950 323.250 ;
        RECT 532.650 317.400 535.950 318.900 ;
        RECT 537.150 317.400 538.950 323.250 ;
        RECT 492.150 315.600 497.250 316.500 ;
        RECT 416.250 314.250 420.000 315.300 ;
        RECT 377.100 312.150 378.900 313.950 ;
        RECT 304.950 308.850 307.350 310.950 ;
        RECT 338.100 310.050 339.900 311.850 ;
        RECT 340.950 310.050 343.050 312.150 ;
        RECT 303.000 305.400 305.250 306.300 ;
        RECT 299.550 304.500 305.250 305.400 ;
        RECT 299.550 297.600 300.750 304.500 ;
        RECT 306.150 303.600 307.350 308.850 ;
        RECT 263.550 291.750 265.350 297.600 ;
        RECT 266.550 291.750 268.350 297.600 ;
        RECT 299.550 291.750 301.350 297.600 ;
        RECT 302.850 291.750 304.650 303.600 ;
        RECT 305.850 291.750 307.650 303.600 ;
        RECT 341.400 297.600 342.600 310.050 ;
        RECT 373.950 308.850 376.050 310.950 ;
        RECT 376.950 310.050 379.050 312.150 ;
        RECT 380.850 310.950 382.050 314.250 ;
        RECT 379.950 308.850 382.050 310.950 ;
        RECT 418.950 310.950 420.150 314.250 ;
        RECT 422.100 312.150 423.900 313.950 ;
        RECT 418.950 308.850 421.050 310.950 ;
        RECT 421.950 310.050 424.050 312.150 ;
        RECT 424.950 308.850 427.050 310.950 ;
        RECT 452.100 309.150 453.900 310.950 ;
        RECT 374.100 307.050 375.900 308.850 ;
        RECT 379.950 303.600 381.150 308.850 ;
        RECT 382.950 305.850 385.050 307.950 ;
        RECT 415.950 305.850 418.050 307.950 ;
        RECT 382.950 304.050 384.750 305.850 ;
        RECT 416.250 304.050 418.050 305.850 ;
        RECT 419.850 303.600 421.050 308.850 ;
        RECT 425.100 307.050 426.900 308.850 ;
        RECT 451.950 307.050 454.050 309.150 ;
        RECT 455.550 307.950 456.750 315.300 ;
        RECT 495.000 314.700 497.250 315.600 ;
        RECT 458.100 309.150 459.900 310.950 ;
        RECT 454.950 305.850 457.050 307.950 ;
        RECT 457.950 307.050 460.050 309.150 ;
        RECT 490.950 308.850 493.050 310.950 ;
        RECT 491.100 307.050 492.900 308.850 ;
        RECT 495.000 306.300 496.050 314.700 ;
        RECT 498.150 310.950 499.350 317.400 ;
        RECT 496.950 308.850 499.350 310.950 ;
        RECT 338.550 291.750 340.350 297.600 ;
        RECT 341.550 291.750 343.350 297.600 ;
        RECT 375.300 291.750 377.100 303.600 ;
        RECT 379.500 291.750 381.300 303.600 ;
        RECT 382.800 291.750 384.600 297.600 ;
        RECT 416.400 291.750 418.200 297.600 ;
        RECT 419.700 291.750 421.500 303.600 ;
        RECT 423.900 291.750 425.700 303.600 ;
        RECT 455.550 297.600 456.750 305.850 ;
        RECT 495.000 305.400 497.250 306.300 ;
        RECT 491.550 304.500 497.250 305.400 ;
        RECT 491.550 297.600 492.750 304.500 ;
        RECT 498.150 303.600 499.350 308.850 ;
        RECT 532.650 310.950 533.850 317.400 ;
        RECT 535.950 315.900 537.750 316.500 ;
        RECT 541.650 315.900 543.450 323.250 ;
        RECT 535.950 314.700 543.450 315.900 ;
        RECT 575.850 316.200 577.650 323.250 ;
        RECT 580.350 317.400 582.150 323.250 ;
        RECT 614.850 316.200 616.650 323.250 ;
        RECT 619.350 317.400 621.150 323.250 ;
        RECT 651.000 317.400 652.800 323.250 ;
        RECT 655.200 319.050 657.000 323.250 ;
        RECT 658.500 320.400 660.300 323.250 ;
        RECT 692.550 320.400 694.350 323.250 ;
        RECT 695.550 320.400 697.350 323.250 ;
        RECT 698.550 320.400 700.350 323.250 ;
        RECT 655.200 317.400 660.900 319.050 ;
        RECT 575.850 315.300 579.450 316.200 ;
        RECT 614.850 315.300 618.450 316.200 ;
        RECT 532.650 308.850 535.050 310.950 ;
        RECT 536.100 309.150 537.900 310.950 ;
        RECT 532.650 303.600 533.850 308.850 ;
        RECT 535.950 307.050 538.050 309.150 ;
        RECT 452.550 291.750 454.350 297.600 ;
        RECT 455.550 291.750 457.350 297.600 ;
        RECT 458.550 291.750 460.350 297.600 ;
        RECT 491.550 291.750 493.350 297.600 ;
        RECT 494.850 291.750 496.650 303.600 ;
        RECT 497.850 291.750 499.650 303.600 ;
        RECT 532.050 291.750 533.850 303.600 ;
        RECT 535.050 291.750 536.850 303.600 ;
        RECT 539.100 297.600 540.300 314.700 ;
        RECT 541.950 308.850 544.050 310.950 ;
        RECT 575.100 309.150 576.900 310.950 ;
        RECT 542.100 307.050 543.900 308.850 ;
        RECT 574.950 307.050 577.050 309.150 ;
        RECT 578.250 307.950 579.450 315.300 ;
        RECT 581.100 309.150 582.900 310.950 ;
        RECT 614.100 309.150 615.900 310.950 ;
        RECT 577.950 305.850 580.050 307.950 ;
        RECT 580.950 307.050 583.050 309.150 ;
        RECT 613.950 307.050 616.050 309.150 ;
        RECT 617.250 307.950 618.450 315.300 ;
        RECT 619.950 315.450 622.050 316.050 ;
        RECT 619.950 314.550 624.450 315.450 ;
        RECT 619.950 313.950 622.050 314.550 ;
        RECT 620.100 309.150 621.900 310.950 ;
        RECT 616.950 305.850 619.050 307.950 ;
        RECT 619.950 307.050 622.050 309.150 ;
        RECT 578.250 297.600 579.450 305.850 ;
        RECT 617.250 297.600 618.450 305.850 ;
        RECT 619.950 303.450 622.050 304.050 ;
        RECT 623.550 303.450 624.450 314.550 ;
        RECT 650.100 312.150 651.900 313.950 ;
        RECT 649.950 310.050 652.050 312.150 ;
        RECT 652.950 311.850 655.050 313.950 ;
        RECT 656.100 312.150 657.900 313.950 ;
        RECT 653.100 310.050 654.900 311.850 ;
        RECT 655.950 310.050 658.050 312.150 ;
        RECT 659.700 310.950 660.900 317.400 ;
        RECT 696.000 313.950 697.050 320.400 ;
        RECT 728.550 315.900 730.350 323.250 ;
        RECT 733.050 317.400 734.850 323.250 ;
        RECT 736.050 318.900 737.850 323.250 ;
        RECT 736.050 317.400 739.350 318.900 ;
        RECT 734.250 315.900 736.050 316.500 ;
        RECT 728.550 314.700 736.050 315.900 ;
        RECT 694.950 311.850 697.050 313.950 ;
        RECT 658.950 308.850 661.050 310.950 ;
        RECT 691.950 308.850 694.050 310.950 ;
        RECT 659.700 303.600 660.900 308.850 ;
        RECT 692.100 307.050 693.900 308.850 ;
        RECT 696.000 304.650 697.050 311.850 ;
        RECT 697.950 308.850 700.050 310.950 ;
        RECT 727.950 308.850 730.050 310.950 ;
        RECT 698.100 307.050 699.900 308.850 ;
        RECT 728.100 307.050 729.900 308.850 ;
        RECT 696.000 303.600 698.550 304.650 ;
        RECT 619.950 302.550 624.450 303.450 ;
        RECT 650.550 302.700 658.350 303.600 ;
        RECT 619.950 301.950 622.050 302.550 ;
        RECT 538.650 291.750 540.450 297.600 ;
        RECT 541.650 291.750 543.450 297.600 ;
        RECT 574.650 291.750 576.450 297.600 ;
        RECT 577.650 291.750 579.450 297.600 ;
        RECT 580.650 291.750 582.450 297.600 ;
        RECT 613.650 291.750 615.450 297.600 ;
        RECT 616.650 291.750 618.450 297.600 ;
        RECT 619.650 291.750 621.450 297.600 ;
        RECT 650.550 291.750 652.350 302.700 ;
        RECT 653.550 291.750 655.350 301.800 ;
        RECT 656.550 291.750 658.350 302.700 ;
        RECT 659.550 291.750 661.350 303.600 ;
        RECT 692.550 291.750 694.350 303.600 ;
        RECT 696.750 291.750 698.550 303.600 ;
        RECT 731.700 297.600 732.900 314.700 ;
        RECT 738.150 310.950 739.350 317.400 ;
        RECT 734.100 309.150 735.900 310.950 ;
        RECT 733.950 307.050 736.050 309.150 ;
        RECT 736.950 308.850 739.350 310.950 ;
        RECT 738.150 303.600 739.350 308.850 ;
        RECT 728.550 291.750 730.350 297.600 ;
        RECT 731.550 291.750 733.350 297.600 ;
        RECT 735.150 291.750 736.950 303.600 ;
        RECT 738.150 291.750 739.950 303.600 ;
        RECT 31.650 275.400 33.450 287.250 ;
        RECT 34.650 276.300 36.450 287.250 ;
        RECT 37.650 277.200 39.450 287.250 ;
        RECT 40.650 276.300 42.450 287.250 ;
        RECT 34.650 275.400 42.450 276.300 ;
        RECT 72.300 275.400 74.100 287.250 ;
        RECT 76.500 275.400 78.300 287.250 ;
        RECT 79.800 281.400 81.600 287.250 ;
        RECT 114.450 275.400 116.250 287.250 ;
        RECT 118.650 275.400 120.450 287.250 ;
        RECT 123.150 275.400 124.950 287.250 ;
        RECT 126.150 281.400 127.950 287.250 ;
        RECT 131.250 281.400 133.050 287.250 ;
        RECT 136.050 281.400 137.850 287.250 ;
        RECT 131.550 280.500 132.750 281.400 ;
        RECT 139.050 280.500 140.850 287.250 ;
        RECT 142.950 281.400 144.750 287.250 ;
        RECT 147.150 281.400 148.950 287.250 ;
        RECT 151.650 284.400 153.450 287.250 ;
        RECT 127.950 278.400 132.750 280.500 ;
        RECT 135.150 278.700 142.050 280.500 ;
        RECT 147.150 279.300 151.050 281.400 ;
        RECT 131.550 277.500 132.750 278.400 ;
        RECT 144.450 277.800 146.250 278.400 ;
        RECT 131.550 276.300 139.050 277.500 ;
        RECT 137.250 275.700 139.050 276.300 ;
        RECT 139.950 276.900 146.250 277.800 ;
        RECT 32.100 270.150 33.300 275.400 ;
        RECT 71.100 270.150 72.900 271.950 ;
        RECT 76.950 270.150 78.150 275.400 ;
        RECT 79.950 273.150 81.750 274.950 ;
        RECT 114.450 274.350 117.000 275.400 ;
        RECT 79.950 271.050 82.050 273.150 ;
        RECT 113.100 270.150 114.900 271.950 ;
        RECT 31.950 268.050 34.050 270.150 ;
        RECT 32.100 261.600 33.300 268.050 ;
        RECT 34.950 266.850 37.050 268.950 ;
        RECT 38.100 267.150 39.900 268.950 ;
        RECT 35.100 265.050 36.900 266.850 ;
        RECT 37.950 265.050 40.050 267.150 ;
        RECT 40.950 266.850 43.050 268.950 ;
        RECT 70.950 268.050 73.050 270.150 ;
        RECT 73.950 266.850 76.050 268.950 ;
        RECT 76.950 268.050 79.050 270.150 ;
        RECT 112.950 268.050 115.050 270.150 ;
        RECT 41.100 265.050 42.900 266.850 ;
        RECT 74.100 265.050 75.900 266.850 ;
        RECT 77.850 264.750 79.050 268.050 ;
        RECT 115.950 267.150 117.000 274.350 ;
        RECT 123.150 274.800 134.250 275.400 ;
        RECT 139.950 274.800 140.850 276.900 ;
        RECT 144.450 276.600 146.250 276.900 ;
        RECT 147.150 276.600 149.850 278.400 ;
        RECT 147.150 275.700 148.050 276.600 ;
        RECT 123.150 274.200 140.850 274.800 ;
        RECT 119.100 270.150 120.900 271.950 ;
        RECT 118.950 268.050 121.050 270.150 ;
        RECT 115.950 265.050 118.050 267.150 ;
        RECT 78.000 263.700 81.750 264.750 ;
        RECT 32.100 259.950 37.800 261.600 ;
        RECT 32.700 255.750 34.500 258.600 ;
        RECT 36.000 255.750 37.800 259.950 ;
        RECT 40.200 255.750 42.000 261.600 ;
        RECT 71.550 260.700 79.350 262.050 ;
        RECT 71.550 255.750 73.350 260.700 ;
        RECT 74.550 255.750 76.350 259.800 ;
        RECT 77.550 255.750 79.350 260.700 ;
        RECT 80.550 261.600 81.750 263.700 ;
        RECT 80.550 255.750 82.350 261.600 ;
        RECT 115.950 258.600 117.000 265.050 ;
        RECT 123.150 261.600 124.050 274.200 ;
        RECT 132.450 273.900 140.850 274.200 ;
        RECT 142.050 274.800 148.050 275.700 ;
        RECT 148.950 274.800 151.050 275.700 ;
        RECT 154.650 275.400 156.450 287.250 ;
        RECT 186.300 275.400 188.100 287.250 ;
        RECT 190.500 275.400 192.300 287.250 ;
        RECT 193.800 281.400 195.600 287.250 ;
        RECT 201.150 275.400 202.950 287.250 ;
        RECT 204.150 281.400 205.950 287.250 ;
        RECT 209.250 281.400 211.050 287.250 ;
        RECT 214.050 281.400 215.850 287.250 ;
        RECT 209.550 280.500 210.750 281.400 ;
        RECT 217.050 280.500 218.850 287.250 ;
        RECT 220.950 281.400 222.750 287.250 ;
        RECT 225.150 281.400 226.950 287.250 ;
        RECT 229.650 284.400 231.450 287.250 ;
        RECT 205.950 278.400 210.750 280.500 ;
        RECT 213.150 278.700 220.050 280.500 ;
        RECT 225.150 279.300 229.050 281.400 ;
        RECT 209.550 277.500 210.750 278.400 ;
        RECT 222.450 277.800 224.250 278.400 ;
        RECT 209.550 276.300 217.050 277.500 ;
        RECT 215.250 275.700 217.050 276.300 ;
        RECT 217.950 276.900 224.250 277.800 ;
        RECT 132.450 273.600 134.250 273.900 ;
        RECT 142.050 270.150 142.950 274.800 ;
        RECT 148.950 273.600 153.150 274.800 ;
        RECT 152.250 271.800 154.050 273.600 ;
        RECT 133.950 269.100 136.050 270.150 ;
        RECT 125.100 267.150 126.900 268.950 ;
        RECT 128.100 268.050 136.050 269.100 ;
        RECT 139.950 268.050 142.950 270.150 ;
        RECT 128.100 267.300 129.900 268.050 ;
        RECT 126.000 266.400 126.900 267.150 ;
        RECT 131.100 266.400 132.900 267.000 ;
        RECT 126.000 265.200 132.900 266.400 ;
        RECT 131.850 264.000 132.900 265.200 ;
        RECT 142.050 264.000 142.950 268.050 ;
        RECT 151.950 267.750 154.050 268.050 ;
        RECT 150.150 265.950 154.050 267.750 ;
        RECT 155.250 265.950 156.450 275.400 ;
        RECT 185.100 270.150 186.900 271.950 ;
        RECT 190.950 270.150 192.150 275.400 ;
        RECT 193.950 273.150 195.750 274.950 ;
        RECT 201.150 274.800 212.250 275.400 ;
        RECT 217.950 274.800 218.850 276.900 ;
        RECT 222.450 276.600 224.250 276.900 ;
        RECT 225.150 276.600 227.850 278.400 ;
        RECT 225.150 275.700 226.050 276.600 ;
        RECT 201.150 274.200 218.850 274.800 ;
        RECT 193.950 271.050 196.050 273.150 ;
        RECT 184.950 268.050 187.050 270.150 ;
        RECT 187.950 266.850 190.050 268.950 ;
        RECT 190.950 268.050 193.050 270.150 ;
        RECT 131.850 263.100 142.950 264.000 ;
        RECT 151.950 263.850 156.450 265.950 ;
        RECT 188.100 265.050 189.900 266.850 ;
        RECT 191.850 264.750 193.050 268.050 ;
        RECT 131.850 262.200 132.900 263.100 ;
        RECT 142.050 262.800 142.950 263.100 ;
        RECT 112.650 255.750 114.450 258.600 ;
        RECT 115.650 255.750 117.450 258.600 ;
        RECT 118.650 255.750 120.450 258.600 ;
        RECT 123.150 255.750 124.950 261.600 ;
        RECT 127.950 259.500 130.050 261.600 ;
        RECT 131.550 260.400 133.350 262.200 ;
        RECT 134.850 261.450 136.650 262.200 ;
        RECT 134.850 260.400 139.800 261.450 ;
        RECT 142.050 261.000 143.850 262.800 ;
        RECT 155.250 261.600 156.450 263.850 ;
        RECT 192.000 263.700 195.750 264.750 ;
        RECT 148.950 260.700 151.050 261.600 ;
        RECT 129.000 258.600 130.050 259.500 ;
        RECT 138.750 258.600 139.800 260.400 ;
        RECT 147.300 259.500 151.050 260.700 ;
        RECT 147.300 258.600 148.350 259.500 ;
        RECT 126.150 255.750 127.950 258.600 ;
        RECT 129.000 257.700 132.750 258.600 ;
        RECT 130.950 255.750 132.750 257.700 ;
        RECT 135.450 255.750 137.250 258.600 ;
        RECT 138.750 255.750 140.550 258.600 ;
        RECT 142.650 255.750 144.450 258.600 ;
        RECT 146.850 255.750 148.650 258.600 ;
        RECT 151.350 255.750 153.150 258.600 ;
        RECT 154.650 255.750 156.450 261.600 ;
        RECT 185.550 260.700 193.350 262.050 ;
        RECT 185.550 255.750 187.350 260.700 ;
        RECT 188.550 255.750 190.350 259.800 ;
        RECT 191.550 255.750 193.350 260.700 ;
        RECT 194.550 261.600 195.750 263.700 ;
        RECT 201.150 261.600 202.050 274.200 ;
        RECT 210.450 273.900 218.850 274.200 ;
        RECT 220.050 274.800 226.050 275.700 ;
        RECT 226.950 274.800 229.050 275.700 ;
        RECT 232.650 275.400 234.450 287.250 ;
        RECT 263.550 276.300 265.350 287.250 ;
        RECT 266.550 277.200 268.350 287.250 ;
        RECT 269.550 276.300 271.350 287.250 ;
        RECT 263.550 275.400 271.350 276.300 ;
        RECT 272.550 275.400 274.350 287.250 ;
        RECT 305.400 281.400 307.200 287.250 ;
        RECT 308.700 275.400 310.500 287.250 ;
        RECT 312.900 275.400 314.700 287.250 ;
        RECT 346.650 275.400 348.450 287.250 ;
        RECT 349.650 276.300 351.450 287.250 ;
        RECT 352.650 277.200 354.450 287.250 ;
        RECT 355.650 276.300 357.450 287.250 ;
        RECT 386.550 281.400 388.350 287.250 ;
        RECT 389.550 281.400 391.350 287.250 ;
        RECT 392.550 281.400 394.350 287.250 ;
        RECT 427.650 281.400 429.450 287.250 ;
        RECT 430.650 281.400 432.450 287.250 ;
        RECT 349.650 275.400 357.450 276.300 ;
        RECT 210.450 273.600 212.250 273.900 ;
        RECT 220.050 270.150 220.950 274.800 ;
        RECT 226.950 273.600 231.150 274.800 ;
        RECT 230.250 271.800 232.050 273.600 ;
        RECT 211.950 269.100 214.050 270.150 ;
        RECT 203.100 267.150 204.900 268.950 ;
        RECT 206.100 268.050 214.050 269.100 ;
        RECT 217.950 268.050 220.950 270.150 ;
        RECT 206.100 267.300 207.900 268.050 ;
        RECT 204.000 266.400 204.900 267.150 ;
        RECT 209.100 266.400 210.900 267.000 ;
        RECT 204.000 265.200 210.900 266.400 ;
        RECT 209.850 264.000 210.900 265.200 ;
        RECT 220.050 264.000 220.950 268.050 ;
        RECT 229.950 267.750 232.050 268.050 ;
        RECT 228.150 265.950 232.050 267.750 ;
        RECT 233.250 265.950 234.450 275.400 ;
        RECT 272.700 270.150 273.900 275.400 ;
        RECT 305.250 273.150 307.050 274.950 ;
        RECT 304.950 271.050 307.050 273.150 ;
        RECT 308.850 270.150 310.050 275.400 ;
        RECT 314.100 270.150 315.900 271.950 ;
        RECT 347.100 270.150 348.300 275.400 ;
        RECT 389.550 273.150 390.750 281.400 ;
        RECT 262.950 266.850 265.050 268.950 ;
        RECT 266.100 267.150 267.900 268.950 ;
        RECT 209.850 263.100 220.950 264.000 ;
        RECT 229.950 263.850 234.450 265.950 ;
        RECT 263.100 265.050 264.900 266.850 ;
        RECT 265.950 265.050 268.050 267.150 ;
        RECT 268.950 266.850 271.050 268.950 ;
        RECT 271.950 268.050 274.050 270.150 ;
        RECT 307.950 268.050 310.050 270.150 ;
        RECT 269.100 265.050 270.900 266.850 ;
        RECT 209.850 262.200 210.900 263.100 ;
        RECT 220.050 262.800 220.950 263.100 ;
        RECT 194.550 255.750 196.350 261.600 ;
        RECT 201.150 255.750 202.950 261.600 ;
        RECT 205.950 259.500 208.050 261.600 ;
        RECT 209.550 260.400 211.350 262.200 ;
        RECT 212.850 261.450 214.650 262.200 ;
        RECT 212.850 260.400 217.800 261.450 ;
        RECT 220.050 261.000 221.850 262.800 ;
        RECT 233.250 261.600 234.450 263.850 ;
        RECT 272.700 261.600 273.900 268.050 ;
        RECT 307.950 264.750 309.150 268.050 ;
        RECT 310.950 266.850 313.050 268.950 ;
        RECT 313.950 268.050 316.050 270.150 ;
        RECT 346.950 268.050 349.050 270.150 ;
        RECT 385.950 269.850 388.050 271.950 ;
        RECT 388.950 271.050 391.050 273.150 ;
        RECT 311.100 265.050 312.900 266.850 ;
        RECT 305.250 263.700 309.000 264.750 ;
        RECT 305.250 261.600 306.450 263.700 ;
        RECT 226.950 260.700 229.050 261.600 ;
        RECT 207.000 258.600 208.050 259.500 ;
        RECT 216.750 258.600 217.800 260.400 ;
        RECT 225.300 259.500 229.050 260.700 ;
        RECT 225.300 258.600 226.350 259.500 ;
        RECT 204.150 255.750 205.950 258.600 ;
        RECT 207.000 257.700 210.750 258.600 ;
        RECT 208.950 255.750 210.750 257.700 ;
        RECT 213.450 255.750 215.250 258.600 ;
        RECT 216.750 255.750 218.550 258.600 ;
        RECT 220.650 255.750 222.450 258.600 ;
        RECT 224.850 255.750 226.650 258.600 ;
        RECT 229.350 255.750 231.150 258.600 ;
        RECT 232.650 255.750 234.450 261.600 ;
        RECT 264.000 255.750 265.800 261.600 ;
        RECT 268.200 259.950 273.900 261.600 ;
        RECT 268.200 255.750 270.000 259.950 ;
        RECT 271.500 255.750 273.300 258.600 ;
        RECT 304.650 255.750 306.450 261.600 ;
        RECT 307.650 260.700 315.450 262.050 ;
        RECT 307.650 255.750 309.450 260.700 ;
        RECT 310.650 255.750 312.450 259.800 ;
        RECT 313.650 255.750 315.450 260.700 ;
        RECT 347.100 261.600 348.300 268.050 ;
        RECT 349.950 266.850 352.050 268.950 ;
        RECT 353.100 267.150 354.900 268.950 ;
        RECT 350.100 265.050 351.900 266.850 ;
        RECT 352.950 265.050 355.050 267.150 ;
        RECT 355.950 266.850 358.050 268.950 ;
        RECT 386.100 268.050 387.900 269.850 ;
        RECT 356.100 265.050 357.900 266.850 ;
        RECT 389.550 263.700 390.750 271.050 ;
        RECT 391.950 269.850 394.050 271.950 ;
        RECT 392.100 268.050 393.900 269.850 ;
        RECT 428.400 268.950 429.600 281.400 ;
        RECT 434.550 275.400 436.350 287.250 ;
        RECT 437.550 284.400 439.350 287.250 ;
        RECT 442.050 281.400 443.850 287.250 ;
        RECT 446.250 281.400 448.050 287.250 ;
        RECT 439.950 279.300 443.850 281.400 ;
        RECT 450.150 280.500 451.950 287.250 ;
        RECT 453.150 281.400 454.950 287.250 ;
        RECT 457.950 281.400 459.750 287.250 ;
        RECT 463.050 281.400 464.850 287.250 ;
        RECT 458.250 280.500 459.450 281.400 ;
        RECT 448.950 278.700 455.850 280.500 ;
        RECT 458.250 278.400 463.050 280.500 ;
        RECT 441.150 276.600 443.850 278.400 ;
        RECT 444.750 277.800 446.550 278.400 ;
        RECT 444.750 276.900 451.050 277.800 ;
        RECT 458.250 277.500 459.450 278.400 ;
        RECT 444.750 276.600 446.550 276.900 ;
        RECT 442.950 275.700 443.850 276.600 ;
        RECT 427.950 266.850 430.050 268.950 ;
        RECT 431.100 267.150 432.900 268.950 ;
        RECT 389.550 262.800 393.150 263.700 ;
        RECT 347.100 259.950 352.800 261.600 ;
        RECT 347.700 255.750 349.500 258.600 ;
        RECT 351.000 255.750 352.800 259.950 ;
        RECT 355.200 255.750 357.000 261.600 ;
        RECT 386.850 255.750 388.650 261.600 ;
        RECT 391.350 255.750 393.150 262.800 ;
        RECT 428.400 258.600 429.600 266.850 ;
        RECT 430.950 265.050 433.050 267.150 ;
        RECT 434.550 265.950 435.750 275.400 ;
        RECT 439.950 274.800 442.050 275.700 ;
        RECT 442.950 274.800 448.950 275.700 ;
        RECT 437.850 273.600 442.050 274.800 ;
        RECT 436.950 271.800 438.750 273.600 ;
        RECT 448.050 270.150 448.950 274.800 ;
        RECT 450.150 274.800 451.050 276.900 ;
        RECT 451.950 276.300 459.450 277.500 ;
        RECT 451.950 275.700 453.750 276.300 ;
        RECT 466.050 275.400 467.850 287.250 ;
        RECT 499.050 275.400 500.850 287.250 ;
        RECT 502.050 275.400 503.850 287.250 ;
        RECT 505.650 281.400 507.450 287.250 ;
        RECT 508.650 281.400 510.450 287.250 ;
        RECT 456.750 274.800 467.850 275.400 ;
        RECT 450.150 274.200 467.850 274.800 ;
        RECT 450.150 273.900 458.550 274.200 ;
        RECT 456.750 273.600 458.550 273.900 ;
        RECT 448.050 268.050 451.050 270.150 ;
        RECT 454.950 269.100 457.050 270.150 ;
        RECT 454.950 268.050 462.900 269.100 ;
        RECT 436.950 267.750 439.050 268.050 ;
        RECT 436.950 265.950 440.850 267.750 ;
        RECT 434.550 263.850 439.050 265.950 ;
        RECT 448.050 264.000 448.950 268.050 ;
        RECT 461.100 267.300 462.900 268.050 ;
        RECT 464.100 267.150 465.900 268.950 ;
        RECT 458.100 266.400 459.900 267.000 ;
        RECT 464.100 266.400 465.000 267.150 ;
        RECT 458.100 265.200 465.000 266.400 ;
        RECT 458.100 264.000 459.150 265.200 ;
        RECT 434.550 261.600 435.750 263.850 ;
        RECT 448.050 263.100 459.150 264.000 ;
        RECT 448.050 262.800 448.950 263.100 ;
        RECT 427.650 255.750 429.450 258.600 ;
        RECT 430.650 255.750 432.450 258.600 ;
        RECT 434.550 255.750 436.350 261.600 ;
        RECT 439.950 260.700 442.050 261.600 ;
        RECT 447.150 261.000 448.950 262.800 ;
        RECT 458.100 262.200 459.150 263.100 ;
        RECT 454.350 261.450 456.150 262.200 ;
        RECT 439.950 259.500 443.700 260.700 ;
        RECT 442.650 258.600 443.700 259.500 ;
        RECT 451.200 260.400 456.150 261.450 ;
        RECT 457.650 260.400 459.450 262.200 ;
        RECT 466.950 261.600 467.850 274.200 ;
        RECT 451.200 258.600 452.250 260.400 ;
        RECT 460.950 259.500 463.050 261.600 ;
        RECT 460.950 258.600 462.000 259.500 ;
        RECT 437.850 255.750 439.650 258.600 ;
        RECT 442.350 255.750 444.150 258.600 ;
        RECT 446.550 255.750 448.350 258.600 ;
        RECT 450.450 255.750 452.250 258.600 ;
        RECT 453.750 255.750 455.550 258.600 ;
        RECT 458.250 257.700 462.000 258.600 ;
        RECT 458.250 255.750 460.050 257.700 ;
        RECT 463.050 255.750 464.850 258.600 ;
        RECT 466.050 255.750 467.850 261.600 ;
        RECT 499.650 270.150 500.850 275.400 ;
        RECT 499.650 268.050 502.050 270.150 ;
        RECT 502.950 269.850 505.050 271.950 ;
        RECT 503.100 268.050 504.900 269.850 ;
        RECT 499.650 261.600 500.850 268.050 ;
        RECT 506.100 264.300 507.300 281.400 ;
        RECT 512.550 275.400 514.350 287.250 ;
        RECT 515.550 284.400 517.350 287.250 ;
        RECT 520.050 281.400 521.850 287.250 ;
        RECT 524.250 281.400 526.050 287.250 ;
        RECT 517.950 279.300 521.850 281.400 ;
        RECT 528.150 280.500 529.950 287.250 ;
        RECT 531.150 281.400 532.950 287.250 ;
        RECT 535.950 281.400 537.750 287.250 ;
        RECT 541.050 281.400 542.850 287.250 ;
        RECT 536.250 280.500 537.450 281.400 ;
        RECT 526.950 278.700 533.850 280.500 ;
        RECT 536.250 278.400 541.050 280.500 ;
        RECT 519.150 276.600 521.850 278.400 ;
        RECT 522.750 277.800 524.550 278.400 ;
        RECT 522.750 276.900 529.050 277.800 ;
        RECT 536.250 277.500 537.450 278.400 ;
        RECT 522.750 276.600 524.550 276.900 ;
        RECT 520.950 275.700 521.850 276.600 ;
        RECT 509.100 270.150 510.900 271.950 ;
        RECT 508.950 268.050 511.050 270.150 ;
        RECT 512.550 265.950 513.750 275.400 ;
        RECT 517.950 274.800 520.050 275.700 ;
        RECT 520.950 274.800 526.950 275.700 ;
        RECT 515.850 273.600 520.050 274.800 ;
        RECT 514.950 271.800 516.750 273.600 ;
        RECT 526.050 270.150 526.950 274.800 ;
        RECT 528.150 274.800 529.050 276.900 ;
        RECT 529.950 276.300 537.450 277.500 ;
        RECT 529.950 275.700 531.750 276.300 ;
        RECT 544.050 275.400 545.850 287.250 ;
        RECT 534.750 274.800 545.850 275.400 ;
        RECT 528.150 274.200 545.850 274.800 ;
        RECT 528.150 273.900 536.550 274.200 ;
        RECT 534.750 273.600 536.550 273.900 ;
        RECT 526.050 268.050 529.050 270.150 ;
        RECT 532.950 269.100 535.050 270.150 ;
        RECT 532.950 268.050 540.900 269.100 ;
        RECT 514.950 267.750 517.050 268.050 ;
        RECT 514.950 265.950 518.850 267.750 ;
        RECT 502.950 263.100 510.450 264.300 ;
        RECT 502.950 262.500 504.750 263.100 ;
        RECT 499.650 260.100 502.950 261.600 ;
        RECT 501.150 255.750 502.950 260.100 ;
        RECT 504.150 255.750 505.950 261.600 ;
        RECT 508.650 255.750 510.450 263.100 ;
        RECT 512.550 263.850 517.050 265.950 ;
        RECT 526.050 264.000 526.950 268.050 ;
        RECT 539.100 267.300 540.900 268.050 ;
        RECT 542.100 267.150 543.900 268.950 ;
        RECT 536.100 266.400 537.900 267.000 ;
        RECT 542.100 266.400 543.000 267.150 ;
        RECT 536.100 265.200 543.000 266.400 ;
        RECT 536.100 264.000 537.150 265.200 ;
        RECT 512.550 261.600 513.750 263.850 ;
        RECT 526.050 263.100 537.150 264.000 ;
        RECT 526.050 262.800 526.950 263.100 ;
        RECT 512.550 255.750 514.350 261.600 ;
        RECT 517.950 260.700 520.050 261.600 ;
        RECT 525.150 261.000 526.950 262.800 ;
        RECT 536.100 262.200 537.150 263.100 ;
        RECT 532.350 261.450 534.150 262.200 ;
        RECT 517.950 259.500 521.700 260.700 ;
        RECT 520.650 258.600 521.700 259.500 ;
        RECT 529.200 260.400 534.150 261.450 ;
        RECT 535.650 260.400 537.450 262.200 ;
        RECT 544.950 261.600 545.850 274.200 ;
        RECT 529.200 258.600 530.250 260.400 ;
        RECT 538.950 259.500 541.050 261.600 ;
        RECT 538.950 258.600 540.000 259.500 ;
        RECT 515.850 255.750 517.650 258.600 ;
        RECT 520.350 255.750 522.150 258.600 ;
        RECT 524.550 255.750 526.350 258.600 ;
        RECT 528.450 255.750 530.250 258.600 ;
        RECT 531.750 255.750 533.550 258.600 ;
        RECT 536.250 257.700 540.000 258.600 ;
        RECT 536.250 255.750 538.050 257.700 ;
        RECT 541.050 255.750 542.850 258.600 ;
        RECT 544.050 255.750 545.850 261.600 ;
        RECT 548.550 275.400 550.350 287.250 ;
        RECT 551.550 284.400 553.350 287.250 ;
        RECT 556.050 281.400 557.850 287.250 ;
        RECT 560.250 281.400 562.050 287.250 ;
        RECT 553.950 279.300 557.850 281.400 ;
        RECT 564.150 280.500 565.950 287.250 ;
        RECT 567.150 281.400 568.950 287.250 ;
        RECT 571.950 281.400 573.750 287.250 ;
        RECT 577.050 281.400 578.850 287.250 ;
        RECT 572.250 280.500 573.450 281.400 ;
        RECT 562.950 278.700 569.850 280.500 ;
        RECT 572.250 278.400 577.050 280.500 ;
        RECT 555.150 276.600 557.850 278.400 ;
        RECT 558.750 277.800 560.550 278.400 ;
        RECT 558.750 276.900 565.050 277.800 ;
        RECT 572.250 277.500 573.450 278.400 ;
        RECT 558.750 276.600 560.550 276.900 ;
        RECT 556.950 275.700 557.850 276.600 ;
        RECT 548.550 265.950 549.750 275.400 ;
        RECT 553.950 274.800 556.050 275.700 ;
        RECT 556.950 274.800 562.950 275.700 ;
        RECT 551.850 273.600 556.050 274.800 ;
        RECT 550.950 271.800 552.750 273.600 ;
        RECT 562.050 270.150 562.950 274.800 ;
        RECT 564.150 274.800 565.050 276.900 ;
        RECT 565.950 276.300 573.450 277.500 ;
        RECT 565.950 275.700 567.750 276.300 ;
        RECT 580.050 275.400 581.850 287.250 ;
        RECT 611.550 281.400 613.350 287.250 ;
        RECT 614.550 281.400 616.350 287.250 ;
        RECT 617.550 281.400 619.350 287.250 ;
        RECT 570.750 274.800 581.850 275.400 ;
        RECT 564.150 274.200 581.850 274.800 ;
        RECT 564.150 273.900 572.550 274.200 ;
        RECT 570.750 273.600 572.550 273.900 ;
        RECT 562.050 268.050 565.050 270.150 ;
        RECT 568.950 269.100 571.050 270.150 ;
        RECT 568.950 268.050 576.900 269.100 ;
        RECT 550.950 267.750 553.050 268.050 ;
        RECT 550.950 265.950 554.850 267.750 ;
        RECT 548.550 263.850 553.050 265.950 ;
        RECT 562.050 264.000 562.950 268.050 ;
        RECT 575.100 267.300 576.900 268.050 ;
        RECT 578.100 267.150 579.900 268.950 ;
        RECT 572.100 266.400 573.900 267.000 ;
        RECT 578.100 266.400 579.000 267.150 ;
        RECT 572.100 265.200 579.000 266.400 ;
        RECT 572.100 264.000 573.150 265.200 ;
        RECT 548.550 261.600 549.750 263.850 ;
        RECT 562.050 263.100 573.150 264.000 ;
        RECT 562.050 262.800 562.950 263.100 ;
        RECT 548.550 255.750 550.350 261.600 ;
        RECT 553.950 260.700 556.050 261.600 ;
        RECT 561.150 261.000 562.950 262.800 ;
        RECT 572.100 262.200 573.150 263.100 ;
        RECT 568.350 261.450 570.150 262.200 ;
        RECT 553.950 259.500 557.700 260.700 ;
        RECT 556.650 258.600 557.700 259.500 ;
        RECT 565.200 260.400 570.150 261.450 ;
        RECT 571.650 260.400 573.450 262.200 ;
        RECT 580.950 261.600 581.850 274.200 ;
        RECT 614.550 273.150 615.750 281.400 ;
        RECT 652.650 275.400 654.450 287.250 ;
        RECT 655.650 276.300 657.450 287.250 ;
        RECT 658.650 277.200 660.450 287.250 ;
        RECT 661.650 276.300 663.450 287.250 ;
        RECT 655.650 275.400 663.450 276.300 ;
        RECT 692.550 275.400 694.350 287.250 ;
        RECT 696.750 275.400 698.550 287.250 ;
        RECT 610.950 269.850 613.050 271.950 ;
        RECT 613.950 271.050 616.050 273.150 ;
        RECT 611.100 268.050 612.900 269.850 ;
        RECT 614.550 263.700 615.750 271.050 ;
        RECT 616.950 269.850 619.050 271.950 ;
        RECT 653.100 270.150 654.300 275.400 ;
        RECT 696.000 274.350 698.550 275.400 ;
        RECT 732.450 275.400 734.250 287.250 ;
        RECT 736.650 275.400 738.450 287.250 ;
        RECT 732.450 274.350 735.000 275.400 ;
        RECT 692.100 270.150 693.900 271.950 ;
        RECT 617.100 268.050 618.900 269.850 ;
        RECT 652.950 268.050 655.050 270.150 ;
        RECT 614.550 262.800 618.150 263.700 ;
        RECT 565.200 258.600 566.250 260.400 ;
        RECT 574.950 259.500 577.050 261.600 ;
        RECT 574.950 258.600 576.000 259.500 ;
        RECT 551.850 255.750 553.650 258.600 ;
        RECT 556.350 255.750 558.150 258.600 ;
        RECT 560.550 255.750 562.350 258.600 ;
        RECT 564.450 255.750 566.250 258.600 ;
        RECT 567.750 255.750 569.550 258.600 ;
        RECT 572.250 257.700 576.000 258.600 ;
        RECT 572.250 255.750 574.050 257.700 ;
        RECT 577.050 255.750 578.850 258.600 ;
        RECT 580.050 255.750 581.850 261.600 ;
        RECT 611.850 255.750 613.650 261.600 ;
        RECT 616.350 255.750 618.150 262.800 ;
        RECT 653.100 261.600 654.300 268.050 ;
        RECT 655.950 266.850 658.050 268.950 ;
        RECT 659.100 267.150 660.900 268.950 ;
        RECT 656.100 265.050 657.900 266.850 ;
        RECT 658.950 265.050 661.050 267.150 ;
        RECT 661.950 266.850 664.050 268.950 ;
        RECT 691.950 268.050 694.050 270.150 ;
        RECT 696.000 267.150 697.050 274.350 ;
        RECT 698.100 270.150 699.900 271.950 ;
        RECT 731.100 270.150 732.900 271.950 ;
        RECT 697.950 268.050 700.050 270.150 ;
        RECT 730.950 268.050 733.050 270.150 ;
        RECT 662.100 265.050 663.900 266.850 ;
        RECT 694.950 265.050 697.050 267.150 ;
        RECT 653.100 259.950 658.800 261.600 ;
        RECT 653.700 255.750 655.500 258.600 ;
        RECT 657.000 255.750 658.800 259.950 ;
        RECT 661.200 255.750 663.000 261.600 ;
        RECT 696.000 258.600 697.050 265.050 ;
        RECT 733.950 267.150 735.000 274.350 ;
        RECT 737.100 270.150 738.900 271.950 ;
        RECT 736.950 268.050 739.050 270.150 ;
        RECT 733.950 265.050 736.050 267.150 ;
        RECT 733.950 258.600 735.000 265.050 ;
        RECT 692.550 255.750 694.350 258.600 ;
        RECT 695.550 255.750 697.350 258.600 ;
        RECT 698.550 255.750 700.350 258.600 ;
        RECT 730.650 255.750 732.450 258.600 ;
        RECT 733.650 255.750 735.450 258.600 ;
        RECT 736.650 255.750 738.450 258.600 ;
        RECT 32.850 244.200 34.650 251.250 ;
        RECT 37.350 245.400 39.150 251.250 ;
        RECT 70.650 248.400 72.450 251.250 ;
        RECT 73.650 248.400 75.450 251.250 ;
        RECT 76.650 248.400 78.450 251.250 ;
        RECT 32.850 243.300 36.450 244.200 ;
        RECT 32.100 237.150 33.900 238.950 ;
        RECT 31.950 235.050 34.050 237.150 ;
        RECT 35.250 235.950 36.450 243.300 ;
        RECT 73.950 241.950 75.000 248.400 ;
        RECT 107.850 244.200 109.650 251.250 ;
        RECT 112.350 245.400 114.150 251.250 ;
        RECT 143.850 245.400 145.650 251.250 ;
        RECT 148.350 244.200 150.150 251.250 ;
        RECT 185.700 248.400 187.500 251.250 ;
        RECT 189.000 247.050 190.800 251.250 ;
        RECT 107.850 243.300 111.450 244.200 ;
        RECT 73.950 239.850 76.050 241.950 ;
        RECT 38.100 237.150 39.900 238.950 ;
        RECT 34.950 233.850 37.050 235.950 ;
        RECT 37.950 235.050 40.050 237.150 ;
        RECT 70.950 236.850 73.050 238.950 ;
        RECT 71.100 235.050 72.900 236.850 ;
        RECT 35.250 225.600 36.450 233.850 ;
        RECT 73.950 232.650 75.000 239.850 ;
        RECT 76.950 236.850 79.050 238.950 ;
        RECT 107.100 237.150 108.900 238.950 ;
        RECT 77.100 235.050 78.900 236.850 ;
        RECT 106.950 235.050 109.050 237.150 ;
        RECT 110.250 235.950 111.450 243.300 ;
        RECT 146.550 243.300 150.150 244.200 ;
        RECT 185.100 245.400 190.800 247.050 ;
        RECT 193.200 245.400 195.000 251.250 ;
        RECT 224.550 246.300 226.350 251.250 ;
        RECT 227.550 247.200 229.350 251.250 ;
        RECT 230.550 246.300 232.350 251.250 ;
        RECT 113.100 237.150 114.900 238.950 ;
        RECT 143.100 237.150 144.900 238.950 ;
        RECT 109.950 233.850 112.050 235.950 ;
        RECT 112.950 235.050 115.050 237.150 ;
        RECT 142.950 235.050 145.050 237.150 ;
        RECT 146.550 235.950 147.750 243.300 ;
        RECT 185.100 238.950 186.300 245.400 ;
        RECT 224.550 244.950 232.350 246.300 ;
        RECT 233.550 245.400 235.350 251.250 ;
        RECT 268.650 245.400 270.450 251.250 ;
        RECT 271.650 245.400 273.450 251.250 ;
        RECT 274.650 245.400 276.450 251.250 ;
        RECT 277.650 245.400 279.450 251.250 ;
        RECT 280.650 245.400 282.450 251.250 ;
        RECT 233.550 243.300 234.750 245.400 ;
        RECT 271.800 244.500 273.600 245.400 ;
        RECT 277.800 244.500 279.600 245.400 ;
        RECT 283.650 244.500 285.450 251.250 ;
        RECT 286.650 245.400 288.450 251.250 ;
        RECT 289.650 245.400 291.450 251.250 ;
        RECT 292.650 245.400 294.450 251.250 ;
        RECT 323.550 245.400 325.350 251.250 ;
        RECT 326.550 245.400 328.350 251.250 ;
        RECT 329.550 245.400 331.350 251.250 ;
        RECT 289.800 244.500 291.600 245.400 ;
        RECT 270.900 244.350 273.600 244.500 ;
        RECT 231.000 242.250 234.750 243.300 ;
        RECT 270.750 243.300 273.600 244.350 ;
        RECT 275.700 243.300 279.600 244.500 ;
        RECT 281.700 243.300 285.450 244.500 ;
        RECT 287.550 243.300 291.600 244.500 ;
        RECT 326.400 244.500 328.200 245.400 ;
        RECT 332.550 244.500 334.350 251.250 ;
        RECT 335.550 245.400 337.350 251.250 ;
        RECT 338.550 245.400 340.350 251.250 ;
        RECT 341.550 245.400 343.350 251.250 ;
        RECT 344.550 245.400 346.350 251.250 ;
        RECT 347.550 245.400 349.350 251.250 ;
        RECT 354.150 245.400 355.950 251.250 ;
        RECT 357.150 248.400 358.950 251.250 ;
        RECT 361.950 249.300 363.750 251.250 ;
        RECT 360.000 248.400 363.750 249.300 ;
        RECT 366.450 248.400 368.250 251.250 ;
        RECT 369.750 248.400 371.550 251.250 ;
        RECT 373.650 248.400 375.450 251.250 ;
        RECT 377.850 248.400 379.650 251.250 ;
        RECT 382.350 248.400 384.150 251.250 ;
        RECT 360.000 247.500 361.050 248.400 ;
        RECT 358.950 245.400 361.050 247.500 ;
        RECT 369.750 246.600 370.800 248.400 ;
        RECT 338.400 244.500 340.200 245.400 ;
        RECT 344.400 244.500 346.200 245.400 ;
        RECT 326.400 243.300 330.450 244.500 ;
        RECT 332.550 243.300 336.300 244.500 ;
        RECT 338.400 243.300 342.300 244.500 ;
        RECT 344.400 244.350 347.100 244.500 ;
        RECT 344.400 243.300 347.250 244.350 ;
        RECT 188.100 240.150 189.900 241.950 ;
        RECT 149.100 237.150 150.900 238.950 ;
        RECT 145.950 233.850 148.050 235.950 ;
        RECT 148.950 235.050 151.050 237.150 ;
        RECT 184.950 236.850 187.050 238.950 ;
        RECT 187.950 238.050 190.050 240.150 ;
        RECT 190.950 239.850 193.050 241.950 ;
        RECT 194.100 240.150 195.900 241.950 ;
        RECT 227.100 240.150 228.900 241.950 ;
        RECT 191.100 238.050 192.900 239.850 ;
        RECT 193.950 238.050 196.050 240.150 ;
        RECT 223.950 236.850 226.050 238.950 ;
        RECT 226.950 238.050 229.050 240.150 ;
        RECT 230.850 238.950 232.050 242.250 ;
        RECT 270.750 240.150 271.800 243.300 ;
        RECT 275.700 242.400 276.900 243.300 ;
        RECT 281.700 242.400 282.900 243.300 ;
        RECT 287.550 242.400 288.750 243.300 ;
        RECT 272.700 240.600 276.900 242.400 ;
        RECT 278.700 240.600 282.900 242.400 ;
        RECT 284.700 240.600 288.750 242.400 ;
        RECT 329.250 242.400 330.450 243.300 ;
        RECT 335.100 242.400 336.300 243.300 ;
        RECT 341.100 242.400 342.300 243.300 ;
        RECT 229.950 236.850 232.050 238.950 ;
        RECT 268.950 238.050 271.800 240.150 ;
        RECT 72.450 231.600 75.000 232.650 ;
        RECT 31.650 219.750 33.450 225.600 ;
        RECT 34.650 219.750 36.450 225.600 ;
        RECT 37.650 219.750 39.450 225.600 ;
        RECT 72.450 219.750 74.250 231.600 ;
        RECT 76.650 219.750 78.450 231.600 ;
        RECT 110.250 225.600 111.450 233.850 ;
        RECT 146.550 225.600 147.750 233.850 ;
        RECT 185.100 231.600 186.300 236.850 ;
        RECT 224.100 235.050 225.900 236.850 ;
        RECT 229.950 231.600 231.150 236.850 ;
        RECT 232.950 233.850 235.050 235.950 ;
        RECT 232.950 232.050 234.750 233.850 ;
        RECT 270.750 233.700 271.800 238.050 ;
        RECT 275.700 233.700 276.900 240.600 ;
        RECT 281.700 233.700 282.900 240.600 ;
        RECT 287.550 233.700 288.750 240.600 ;
        RECT 290.100 240.150 291.900 241.950 ;
        RECT 326.100 240.150 327.900 241.950 ;
        RECT 329.250 240.600 333.300 242.400 ;
        RECT 335.100 240.600 339.300 242.400 ;
        RECT 341.100 240.600 345.300 242.400 ;
        RECT 289.950 238.050 292.050 240.150 ;
        RECT 325.950 238.050 328.050 240.150 ;
        RECT 329.250 233.700 330.450 240.600 ;
        RECT 335.100 233.700 336.300 240.600 ;
        RECT 341.100 233.700 342.300 240.600 ;
        RECT 346.200 240.150 347.250 243.300 ;
        RECT 346.200 238.050 349.050 240.150 ;
        RECT 346.200 233.700 347.250 238.050 ;
        RECT 270.750 232.500 273.450 233.700 ;
        RECT 275.700 232.500 279.450 233.700 ;
        RECT 281.700 232.500 285.450 233.700 ;
        RECT 287.550 232.500 291.450 233.700 ;
        RECT 106.650 219.750 108.450 225.600 ;
        RECT 109.650 219.750 111.450 225.600 ;
        RECT 112.650 219.750 114.450 225.600 ;
        RECT 143.550 219.750 145.350 225.600 ;
        RECT 146.550 219.750 148.350 225.600 ;
        RECT 149.550 219.750 151.350 225.600 ;
        RECT 184.650 219.750 186.450 231.600 ;
        RECT 187.650 230.700 195.450 231.600 ;
        RECT 187.650 219.750 189.450 230.700 ;
        RECT 190.650 219.750 192.450 229.800 ;
        RECT 193.650 219.750 195.450 230.700 ;
        RECT 225.300 219.750 227.100 231.600 ;
        RECT 229.500 219.750 231.300 231.600 ;
        RECT 232.800 219.750 234.600 225.600 ;
        RECT 268.650 219.750 270.450 231.600 ;
        RECT 271.650 219.750 273.450 232.500 ;
        RECT 274.650 219.750 276.450 231.600 ;
        RECT 277.650 219.750 279.450 232.500 ;
        RECT 280.650 219.750 282.450 231.600 ;
        RECT 283.650 219.750 285.450 232.500 ;
        RECT 286.650 219.750 288.450 231.600 ;
        RECT 289.650 219.750 291.450 232.500 ;
        RECT 326.550 232.500 330.450 233.700 ;
        RECT 332.550 232.500 336.300 233.700 ;
        RECT 338.550 232.500 342.300 233.700 ;
        RECT 344.550 232.500 347.250 233.700 ;
        RECT 354.150 232.800 355.050 245.400 ;
        RECT 362.550 244.800 364.350 246.600 ;
        RECT 365.850 245.550 370.800 246.600 ;
        RECT 378.300 247.500 379.350 248.400 ;
        RECT 378.300 246.300 382.050 247.500 ;
        RECT 365.850 244.800 367.650 245.550 ;
        RECT 362.850 243.900 363.900 244.800 ;
        RECT 373.050 244.200 374.850 246.000 ;
        RECT 379.950 245.400 382.050 246.300 ;
        RECT 385.650 245.400 387.450 251.250 ;
        RECT 416.850 245.400 418.650 251.250 ;
        RECT 373.050 243.900 373.950 244.200 ;
        RECT 362.850 243.000 373.950 243.900 ;
        RECT 386.250 243.150 387.450 245.400 ;
        RECT 421.350 244.200 423.150 251.250 ;
        RECT 362.850 241.800 363.900 243.000 ;
        RECT 357.000 240.600 363.900 241.800 ;
        RECT 357.000 239.850 357.900 240.600 ;
        RECT 362.100 240.000 363.900 240.600 ;
        RECT 356.100 238.050 357.900 239.850 ;
        RECT 359.100 238.950 360.900 239.700 ;
        RECT 373.050 238.950 373.950 243.000 ;
        RECT 382.950 241.050 387.450 243.150 ;
        RECT 381.150 239.250 385.050 241.050 ;
        RECT 382.950 238.950 385.050 239.250 ;
        RECT 359.100 237.900 367.050 238.950 ;
        RECT 364.950 236.850 367.050 237.900 ;
        RECT 370.950 236.850 373.950 238.950 ;
        RECT 363.450 233.100 365.250 233.400 ;
        RECT 363.450 232.800 371.850 233.100 ;
        RECT 292.650 219.750 294.450 231.600 ;
        RECT 323.550 219.750 325.350 231.600 ;
        RECT 326.550 219.750 328.350 232.500 ;
        RECT 329.550 219.750 331.350 231.600 ;
        RECT 332.550 219.750 334.350 232.500 ;
        RECT 335.550 219.750 337.350 231.600 ;
        RECT 338.550 219.750 340.350 232.500 ;
        RECT 341.550 219.750 343.350 231.600 ;
        RECT 344.550 219.750 346.350 232.500 ;
        RECT 354.150 232.200 371.850 232.800 ;
        RECT 354.150 231.600 365.250 232.200 ;
        RECT 347.550 219.750 349.350 231.600 ;
        RECT 354.150 219.750 355.950 231.600 ;
        RECT 368.250 230.700 370.050 231.300 ;
        RECT 362.550 229.500 370.050 230.700 ;
        RECT 370.950 230.100 371.850 232.200 ;
        RECT 373.050 232.200 373.950 236.850 ;
        RECT 383.250 233.400 385.050 235.200 ;
        RECT 379.950 232.200 384.150 233.400 ;
        RECT 373.050 231.300 379.050 232.200 ;
        RECT 379.950 231.300 382.050 232.200 ;
        RECT 386.250 231.600 387.450 241.050 ;
        RECT 419.550 243.300 423.150 244.200 ;
        RECT 429.150 245.400 430.950 251.250 ;
        RECT 432.150 248.400 433.950 251.250 ;
        RECT 436.950 249.300 438.750 251.250 ;
        RECT 435.000 248.400 438.750 249.300 ;
        RECT 441.450 248.400 443.250 251.250 ;
        RECT 444.750 248.400 446.550 251.250 ;
        RECT 448.650 248.400 450.450 251.250 ;
        RECT 452.850 248.400 454.650 251.250 ;
        RECT 457.350 248.400 459.150 251.250 ;
        RECT 435.000 247.500 436.050 248.400 ;
        RECT 433.950 245.400 436.050 247.500 ;
        RECT 444.750 246.600 445.800 248.400 ;
        RECT 416.100 237.150 417.900 238.950 ;
        RECT 415.950 235.050 418.050 237.150 ;
        RECT 419.550 235.950 420.750 243.300 ;
        RECT 422.100 237.150 423.900 238.950 ;
        RECT 418.950 233.850 421.050 235.950 ;
        RECT 421.950 235.050 424.050 237.150 ;
        RECT 378.150 230.400 379.050 231.300 ;
        RECT 375.450 230.100 377.250 230.400 ;
        RECT 362.550 228.600 363.750 229.500 ;
        RECT 370.950 229.200 377.250 230.100 ;
        RECT 375.450 228.600 377.250 229.200 ;
        RECT 378.150 228.600 380.850 230.400 ;
        RECT 358.950 226.500 363.750 228.600 ;
        RECT 366.150 226.500 373.050 228.300 ;
        RECT 362.550 225.600 363.750 226.500 ;
        RECT 357.150 219.750 358.950 225.600 ;
        RECT 362.250 219.750 364.050 225.600 ;
        RECT 367.050 219.750 368.850 225.600 ;
        RECT 370.050 219.750 371.850 226.500 ;
        RECT 378.150 225.600 382.050 227.700 ;
        RECT 373.950 219.750 375.750 225.600 ;
        RECT 378.150 219.750 379.950 225.600 ;
        RECT 382.650 219.750 384.450 222.600 ;
        RECT 385.650 219.750 387.450 231.600 ;
        RECT 419.550 225.600 420.750 233.850 ;
        RECT 429.150 232.800 430.050 245.400 ;
        RECT 437.550 244.800 439.350 246.600 ;
        RECT 440.850 245.550 445.800 246.600 ;
        RECT 453.300 247.500 454.350 248.400 ;
        RECT 453.300 246.300 457.050 247.500 ;
        RECT 440.850 244.800 442.650 245.550 ;
        RECT 437.850 243.900 438.900 244.800 ;
        RECT 448.050 244.200 449.850 246.000 ;
        RECT 454.950 245.400 457.050 246.300 ;
        RECT 460.650 245.400 462.450 251.250 ;
        RECT 491.850 245.400 493.650 251.250 ;
        RECT 448.050 243.900 448.950 244.200 ;
        RECT 437.850 243.000 448.950 243.900 ;
        RECT 461.250 243.150 462.450 245.400 ;
        RECT 496.350 244.200 498.150 251.250 ;
        RECT 529.650 245.400 531.450 251.250 ;
        RECT 437.850 241.800 438.900 243.000 ;
        RECT 432.000 240.600 438.900 241.800 ;
        RECT 432.000 239.850 432.900 240.600 ;
        RECT 437.100 240.000 438.900 240.600 ;
        RECT 431.100 238.050 432.900 239.850 ;
        RECT 434.100 238.950 435.900 239.700 ;
        RECT 448.050 238.950 448.950 243.000 ;
        RECT 457.950 241.050 462.450 243.150 ;
        RECT 456.150 239.250 460.050 241.050 ;
        RECT 457.950 238.950 460.050 239.250 ;
        RECT 434.100 237.900 442.050 238.950 ;
        RECT 439.950 236.850 442.050 237.900 ;
        RECT 445.950 236.850 448.950 238.950 ;
        RECT 438.450 233.100 440.250 233.400 ;
        RECT 438.450 232.800 446.850 233.100 ;
        RECT 429.150 232.200 446.850 232.800 ;
        RECT 429.150 231.600 440.250 232.200 ;
        RECT 416.550 219.750 418.350 225.600 ;
        RECT 419.550 219.750 421.350 225.600 ;
        RECT 422.550 219.750 424.350 225.600 ;
        RECT 429.150 219.750 430.950 231.600 ;
        RECT 443.250 230.700 445.050 231.300 ;
        RECT 437.550 229.500 445.050 230.700 ;
        RECT 445.950 230.100 446.850 232.200 ;
        RECT 448.050 232.200 448.950 236.850 ;
        RECT 458.250 233.400 460.050 235.200 ;
        RECT 454.950 232.200 459.150 233.400 ;
        RECT 448.050 231.300 454.050 232.200 ;
        RECT 454.950 231.300 457.050 232.200 ;
        RECT 461.250 231.600 462.450 241.050 ;
        RECT 494.550 243.300 498.150 244.200 ;
        RECT 530.250 243.300 531.450 245.400 ;
        RECT 532.650 246.300 534.450 251.250 ;
        RECT 535.650 247.200 537.450 251.250 ;
        RECT 538.650 246.300 540.450 251.250 ;
        RECT 572.700 248.400 574.500 251.250 ;
        RECT 576.000 247.050 577.800 251.250 ;
        RECT 532.650 244.950 540.450 246.300 ;
        RECT 572.100 245.400 577.800 247.050 ;
        RECT 580.200 245.400 582.000 251.250 ;
        RECT 614.700 248.400 616.500 251.250 ;
        RECT 618.000 247.050 619.800 251.250 ;
        RECT 614.100 245.400 619.800 247.050 ;
        RECT 622.200 245.400 624.000 251.250 ;
        RECT 655.650 245.400 657.450 251.250 ;
        RECT 658.650 248.400 660.450 251.250 ;
        RECT 661.650 248.400 663.450 251.250 ;
        RECT 664.650 248.400 666.450 251.250 ;
        RECT 491.100 237.150 492.900 238.950 ;
        RECT 490.950 235.050 493.050 237.150 ;
        RECT 494.550 235.950 495.750 243.300 ;
        RECT 530.250 242.250 534.000 243.300 ;
        RECT 532.950 238.950 534.150 242.250 ;
        RECT 536.100 240.150 537.900 241.950 ;
        RECT 497.100 237.150 498.900 238.950 ;
        RECT 493.950 233.850 496.050 235.950 ;
        RECT 496.950 235.050 499.050 237.150 ;
        RECT 532.950 236.850 535.050 238.950 ;
        RECT 535.950 238.050 538.050 240.150 ;
        RECT 572.100 238.950 573.300 245.400 ;
        RECT 575.100 240.150 576.900 241.950 ;
        RECT 538.950 236.850 541.050 238.950 ;
        RECT 571.950 236.850 574.050 238.950 ;
        RECT 574.950 238.050 577.050 240.150 ;
        RECT 577.950 239.850 580.050 241.950 ;
        RECT 581.100 240.150 582.900 241.950 ;
        RECT 578.100 238.050 579.900 239.850 ;
        RECT 580.950 238.050 583.050 240.150 ;
        RECT 614.100 238.950 615.300 245.400 ;
        RECT 617.100 240.150 618.900 241.950 ;
        RECT 613.950 236.850 616.050 238.950 ;
        RECT 616.950 238.050 619.050 240.150 ;
        RECT 619.950 239.850 622.050 241.950 ;
        RECT 623.100 240.150 624.900 241.950 ;
        RECT 655.950 240.150 657.000 245.400 ;
        RECT 661.650 244.200 662.550 248.400 ;
        RECT 659.250 243.300 662.550 244.200 ;
        RECT 695.550 243.900 697.350 251.250 ;
        RECT 700.050 245.400 701.850 251.250 ;
        RECT 703.050 246.900 704.850 251.250 ;
        RECT 737.550 248.400 739.350 251.250 ;
        RECT 740.550 248.400 742.350 251.250 ;
        RECT 743.550 248.400 745.350 251.250 ;
        RECT 703.050 245.400 706.350 246.900 ;
        RECT 701.250 243.900 703.050 244.500 ;
        RECT 659.250 242.400 661.050 243.300 ;
        RECT 695.550 242.700 703.050 243.900 ;
        RECT 620.100 238.050 621.900 239.850 ;
        RECT 622.950 238.050 625.050 240.150 ;
        RECT 655.950 238.050 658.050 240.150 ;
        RECT 529.950 233.850 532.050 235.950 ;
        RECT 453.150 230.400 454.050 231.300 ;
        RECT 450.450 230.100 452.250 230.400 ;
        RECT 437.550 228.600 438.750 229.500 ;
        RECT 445.950 229.200 452.250 230.100 ;
        RECT 450.450 228.600 452.250 229.200 ;
        RECT 453.150 228.600 455.850 230.400 ;
        RECT 433.950 226.500 438.750 228.600 ;
        RECT 441.150 226.500 448.050 228.300 ;
        RECT 437.550 225.600 438.750 226.500 ;
        RECT 432.150 219.750 433.950 225.600 ;
        RECT 437.250 219.750 439.050 225.600 ;
        RECT 442.050 219.750 443.850 225.600 ;
        RECT 445.050 219.750 446.850 226.500 ;
        RECT 453.150 225.600 457.050 227.700 ;
        RECT 448.950 219.750 450.750 225.600 ;
        RECT 453.150 219.750 454.950 225.600 ;
        RECT 457.650 219.750 459.450 222.600 ;
        RECT 460.650 219.750 462.450 231.600 ;
        RECT 494.550 225.600 495.750 233.850 ;
        RECT 530.250 232.050 532.050 233.850 ;
        RECT 533.850 231.600 535.050 236.850 ;
        RECT 539.100 235.050 540.900 236.850 ;
        RECT 572.100 231.600 573.300 236.850 ;
        RECT 614.100 231.600 615.300 236.850 ;
        RECT 491.550 219.750 493.350 225.600 ;
        RECT 494.550 219.750 496.350 225.600 ;
        RECT 497.550 219.750 499.350 225.600 ;
        RECT 530.400 219.750 532.200 225.600 ;
        RECT 533.700 219.750 535.500 231.600 ;
        RECT 537.900 219.750 539.700 231.600 ;
        RECT 571.650 219.750 573.450 231.600 ;
        RECT 574.650 230.700 582.450 231.600 ;
        RECT 574.650 219.750 576.450 230.700 ;
        RECT 577.650 219.750 579.450 229.800 ;
        RECT 580.650 219.750 582.450 230.700 ;
        RECT 613.650 219.750 615.450 231.600 ;
        RECT 616.650 230.700 624.450 231.600 ;
        RECT 616.650 219.750 618.450 230.700 ;
        RECT 619.650 219.750 621.450 229.800 ;
        RECT 622.650 219.750 624.450 230.700 ;
        RECT 656.550 231.450 657.900 238.050 ;
        RECT 659.400 234.150 660.300 242.400 ;
        RECT 664.950 239.850 667.050 241.950 ;
        RECT 661.950 236.850 664.050 238.950 ;
        RECT 665.100 238.050 666.900 239.850 ;
        RECT 694.950 236.850 697.050 238.950 ;
        RECT 662.100 235.050 663.900 236.850 ;
        RECT 695.100 235.050 696.900 236.850 ;
        RECT 659.250 234.000 661.050 234.150 ;
        RECT 659.250 232.800 666.450 234.000 ;
        RECT 659.250 232.350 661.050 232.800 ;
        RECT 665.250 231.600 666.450 232.800 ;
        RECT 656.550 230.100 658.950 231.450 ;
        RECT 657.150 219.750 658.950 230.100 ;
        RECT 660.150 219.750 661.950 231.450 ;
        RECT 664.650 219.750 666.450 231.600 ;
        RECT 698.700 225.600 699.900 242.700 ;
        RECT 705.150 238.950 706.350 245.400 ;
        RECT 741.000 241.950 742.050 248.400 ;
        RECT 739.950 239.850 742.050 241.950 ;
        RECT 701.100 237.150 702.900 238.950 ;
        RECT 700.950 235.050 703.050 237.150 ;
        RECT 703.950 236.850 706.350 238.950 ;
        RECT 736.950 236.850 739.050 238.950 ;
        RECT 705.150 231.600 706.350 236.850 ;
        RECT 737.100 235.050 738.900 236.850 ;
        RECT 741.000 232.650 742.050 239.850 ;
        RECT 742.950 236.850 745.050 238.950 ;
        RECT 743.100 235.050 744.900 236.850 ;
        RECT 741.000 231.600 743.550 232.650 ;
        RECT 695.550 219.750 697.350 225.600 ;
        RECT 698.550 219.750 700.350 225.600 ;
        RECT 702.150 219.750 703.950 231.600 ;
        RECT 705.150 219.750 706.950 231.600 ;
        RECT 737.550 219.750 739.350 231.600 ;
        RECT 741.750 219.750 743.550 231.600 ;
        RECT 30.450 203.400 32.250 215.250 ;
        RECT 34.650 203.400 36.450 215.250 ;
        RECT 69.450 203.400 71.250 215.250 ;
        RECT 73.650 203.400 75.450 215.250 ;
        RECT 105.300 203.400 107.100 215.250 ;
        RECT 109.500 203.400 111.300 215.250 ;
        RECT 112.800 209.400 114.600 215.250 ;
        RECT 146.550 209.400 148.350 215.250 ;
        RECT 149.550 209.400 151.350 215.250 ;
        RECT 152.550 209.400 154.350 215.250 ;
        RECT 30.450 202.350 33.000 203.400 ;
        RECT 69.450 202.350 72.000 203.400 ;
        RECT 29.100 198.150 30.900 199.950 ;
        RECT 28.950 196.050 31.050 198.150 ;
        RECT 31.950 195.150 33.000 202.350 ;
        RECT 35.100 198.150 36.900 199.950 ;
        RECT 68.100 198.150 69.900 199.950 ;
        RECT 34.950 196.050 37.050 198.150 ;
        RECT 67.950 196.050 70.050 198.150 ;
        RECT 70.950 195.150 72.000 202.350 ;
        RECT 74.100 198.150 75.900 199.950 ;
        RECT 104.100 198.150 105.900 199.950 ;
        RECT 109.950 198.150 111.150 203.400 ;
        RECT 112.950 201.150 114.750 202.950 ;
        RECT 149.550 201.150 150.750 209.400 ;
        RECT 185.550 203.400 187.350 215.250 ;
        RECT 189.750 203.400 191.550 215.250 ;
        RECT 221.550 209.400 223.350 215.250 ;
        RECT 224.550 209.400 226.350 215.250 ;
        RECT 227.550 209.400 229.350 215.250 ;
        RECT 260.550 209.400 262.350 215.250 ;
        RECT 263.550 209.400 265.350 215.250 ;
        RECT 266.550 209.400 268.350 215.250 ;
        RECT 189.000 202.350 191.550 203.400 ;
        RECT 112.950 199.050 115.050 201.150 ;
        RECT 73.950 196.050 76.050 198.150 ;
        RECT 103.950 196.050 106.050 198.150 ;
        RECT 31.950 193.050 34.050 195.150 ;
        RECT 70.950 193.050 73.050 195.150 ;
        RECT 106.950 194.850 109.050 196.950 ;
        RECT 109.950 196.050 112.050 198.150 ;
        RECT 145.950 197.850 148.050 199.950 ;
        RECT 148.950 199.050 151.050 201.150 ;
        RECT 146.100 196.050 147.900 197.850 ;
        RECT 107.100 193.050 108.900 194.850 ;
        RECT 31.950 186.600 33.000 193.050 ;
        RECT 70.950 186.600 72.000 193.050 ;
        RECT 110.850 192.750 112.050 196.050 ;
        RECT 111.000 191.700 114.750 192.750 ;
        RECT 104.550 188.700 112.350 190.050 ;
        RECT 28.650 183.750 30.450 186.600 ;
        RECT 31.650 183.750 33.450 186.600 ;
        RECT 34.650 183.750 36.450 186.600 ;
        RECT 67.650 183.750 69.450 186.600 ;
        RECT 70.650 183.750 72.450 186.600 ;
        RECT 73.650 183.750 75.450 186.600 ;
        RECT 104.550 183.750 106.350 188.700 ;
        RECT 107.550 183.750 109.350 187.800 ;
        RECT 110.550 183.750 112.350 188.700 ;
        RECT 113.550 189.600 114.750 191.700 ;
        RECT 149.550 191.700 150.750 199.050 ;
        RECT 151.950 197.850 154.050 199.950 ;
        RECT 185.100 198.150 186.900 199.950 ;
        RECT 152.100 196.050 153.900 197.850 ;
        RECT 184.950 196.050 187.050 198.150 ;
        RECT 189.000 195.150 190.050 202.350 ;
        RECT 224.550 201.150 225.750 209.400 ;
        RECT 263.550 201.150 264.750 209.400 ;
        RECT 301.350 203.400 303.150 215.250 ;
        RECT 304.350 203.400 306.150 215.250 ;
        RECT 307.650 209.400 309.450 215.250 ;
        RECT 191.100 198.150 192.900 199.950 ;
        RECT 190.950 196.050 193.050 198.150 ;
        RECT 220.950 197.850 223.050 199.950 ;
        RECT 223.950 199.050 226.050 201.150 ;
        RECT 221.100 196.050 222.900 197.850 ;
        RECT 187.950 193.050 190.050 195.150 ;
        RECT 149.550 190.800 153.150 191.700 ;
        RECT 113.550 183.750 115.350 189.600 ;
        RECT 146.850 183.750 148.650 189.600 ;
        RECT 151.350 183.750 153.150 190.800 ;
        RECT 189.000 186.600 190.050 193.050 ;
        RECT 224.550 191.700 225.750 199.050 ;
        RECT 226.950 197.850 229.050 199.950 ;
        RECT 259.950 197.850 262.050 199.950 ;
        RECT 262.950 199.050 265.050 201.150 ;
        RECT 227.100 196.050 228.900 197.850 ;
        RECT 260.100 196.050 261.900 197.850 ;
        RECT 263.550 191.700 264.750 199.050 ;
        RECT 265.950 197.850 268.050 199.950 ;
        RECT 301.650 198.150 302.850 203.400 ;
        RECT 308.250 202.500 309.450 209.400 ;
        RECT 303.750 201.600 309.450 202.500 ;
        RECT 338.550 209.400 340.350 215.250 ;
        RECT 338.550 202.500 339.750 209.400 ;
        RECT 341.850 203.400 343.650 215.250 ;
        RECT 344.850 203.400 346.650 215.250 ;
        RECT 377.550 209.400 379.350 215.250 ;
        RECT 338.550 201.600 344.250 202.500 ;
        RECT 303.750 200.700 306.000 201.600 ;
        RECT 266.100 196.050 267.900 197.850 ;
        RECT 301.650 196.050 304.050 198.150 ;
        RECT 224.550 190.800 228.150 191.700 ;
        RECT 263.550 190.800 267.150 191.700 ;
        RECT 185.550 183.750 187.350 186.600 ;
        RECT 188.550 183.750 190.350 186.600 ;
        RECT 191.550 183.750 193.350 186.600 ;
        RECT 221.850 183.750 223.650 189.600 ;
        RECT 226.350 183.750 228.150 190.800 ;
        RECT 260.850 183.750 262.650 189.600 ;
        RECT 265.350 183.750 267.150 190.800 ;
        RECT 301.650 189.600 302.850 196.050 ;
        RECT 304.950 192.300 306.000 200.700 ;
        RECT 342.000 200.700 344.250 201.600 ;
        RECT 308.100 198.150 309.900 199.950 ;
        RECT 338.100 198.150 339.900 199.950 ;
        RECT 307.950 196.050 310.050 198.150 ;
        RECT 337.950 196.050 340.050 198.150 ;
        RECT 303.750 191.400 306.000 192.300 ;
        RECT 342.000 192.300 343.050 200.700 ;
        RECT 345.150 198.150 346.350 203.400 ;
        RECT 377.550 202.500 378.750 209.400 ;
        RECT 380.850 203.400 382.650 215.250 ;
        RECT 383.850 203.400 385.650 215.250 ;
        RECT 416.550 209.400 418.350 215.250 ;
        RECT 377.550 201.600 383.250 202.500 ;
        RECT 381.000 200.700 383.250 201.600 ;
        RECT 377.100 198.150 378.900 199.950 ;
        RECT 343.950 196.050 346.350 198.150 ;
        RECT 376.950 196.050 379.050 198.150 ;
        RECT 342.000 191.400 344.250 192.300 ;
        RECT 303.750 190.500 308.850 191.400 ;
        RECT 301.350 183.750 303.150 189.600 ;
        RECT 304.350 183.750 306.150 189.600 ;
        RECT 307.650 186.600 308.850 190.500 ;
        RECT 339.150 190.500 344.250 191.400 ;
        RECT 339.150 186.600 340.350 190.500 ;
        RECT 345.150 189.600 346.350 196.050 ;
        RECT 381.000 192.300 382.050 200.700 ;
        RECT 384.150 198.150 385.350 203.400 ;
        RECT 416.550 202.500 417.750 209.400 ;
        RECT 419.850 203.400 421.650 215.250 ;
        RECT 422.850 203.400 424.650 215.250 ;
        RECT 459.450 203.400 461.250 215.250 ;
        RECT 463.650 203.400 465.450 215.250 ;
        RECT 494.550 209.400 496.350 215.250 ;
        RECT 497.550 209.400 499.350 215.250 ;
        RECT 533.400 209.400 535.200 215.250 ;
        RECT 416.550 201.600 422.250 202.500 ;
        RECT 420.000 200.700 422.250 201.600 ;
        RECT 416.100 198.150 417.900 199.950 ;
        RECT 382.950 196.050 385.350 198.150 ;
        RECT 415.950 196.050 418.050 198.150 ;
        RECT 381.000 191.400 383.250 192.300 ;
        RECT 378.150 190.500 383.250 191.400 ;
        RECT 307.650 183.750 309.450 186.600 ;
        RECT 338.550 183.750 340.350 186.600 ;
        RECT 341.850 183.750 343.650 189.600 ;
        RECT 344.850 183.750 346.650 189.600 ;
        RECT 378.150 186.600 379.350 190.500 ;
        RECT 384.150 189.600 385.350 196.050 ;
        RECT 420.000 192.300 421.050 200.700 ;
        RECT 423.150 198.150 424.350 203.400 ;
        RECT 459.450 202.350 462.000 203.400 ;
        RECT 458.100 198.150 459.900 199.950 ;
        RECT 421.950 196.050 424.350 198.150 ;
        RECT 457.950 196.050 460.050 198.150 ;
        RECT 420.000 191.400 422.250 192.300 ;
        RECT 417.150 190.500 422.250 191.400 ;
        RECT 377.550 183.750 379.350 186.600 ;
        RECT 380.850 183.750 382.650 189.600 ;
        RECT 383.850 183.750 385.650 189.600 ;
        RECT 417.150 186.600 418.350 190.500 ;
        RECT 423.150 189.600 424.350 196.050 ;
        RECT 460.950 195.150 462.000 202.350 ;
        RECT 464.100 198.150 465.900 199.950 ;
        RECT 463.950 196.050 466.050 198.150 ;
        RECT 497.400 196.950 498.600 209.400 ;
        RECT 536.700 203.400 538.500 215.250 ;
        RECT 540.900 203.400 542.700 215.250 ;
        RECT 545.550 203.400 547.350 215.250 ;
        RECT 548.550 212.400 550.350 215.250 ;
        RECT 553.050 209.400 554.850 215.250 ;
        RECT 557.250 209.400 559.050 215.250 ;
        RECT 550.950 207.300 554.850 209.400 ;
        RECT 561.150 208.500 562.950 215.250 ;
        RECT 564.150 209.400 565.950 215.250 ;
        RECT 568.950 209.400 570.750 215.250 ;
        RECT 574.050 209.400 575.850 215.250 ;
        RECT 569.250 208.500 570.450 209.400 ;
        RECT 559.950 206.700 566.850 208.500 ;
        RECT 569.250 206.400 574.050 208.500 ;
        RECT 552.150 204.600 554.850 206.400 ;
        RECT 555.750 205.800 557.550 206.400 ;
        RECT 555.750 204.900 562.050 205.800 ;
        RECT 569.250 205.500 570.450 206.400 ;
        RECT 555.750 204.600 557.550 204.900 ;
        RECT 553.950 203.700 554.850 204.600 ;
        RECT 533.250 201.150 535.050 202.950 ;
        RECT 532.950 199.050 535.050 201.150 ;
        RECT 536.850 198.150 538.050 203.400 ;
        RECT 542.100 198.150 543.900 199.950 ;
        RECT 494.100 195.150 495.900 196.950 ;
        RECT 460.950 193.050 463.050 195.150 ;
        RECT 493.950 193.050 496.050 195.150 ;
        RECT 496.950 194.850 499.050 196.950 ;
        RECT 535.950 196.050 538.050 198.150 ;
        RECT 416.550 183.750 418.350 186.600 ;
        RECT 419.850 183.750 421.650 189.600 ;
        RECT 422.850 183.750 424.650 189.600 ;
        RECT 460.950 186.600 462.000 193.050 ;
        RECT 497.400 186.600 498.600 194.850 ;
        RECT 535.950 192.750 537.150 196.050 ;
        RECT 538.950 194.850 541.050 196.950 ;
        RECT 541.950 196.050 544.050 198.150 ;
        RECT 539.100 193.050 540.900 194.850 ;
        RECT 545.550 193.950 546.750 203.400 ;
        RECT 550.950 202.800 553.050 203.700 ;
        RECT 553.950 202.800 559.950 203.700 ;
        RECT 548.850 201.600 553.050 202.800 ;
        RECT 547.950 199.800 549.750 201.600 ;
        RECT 559.050 198.150 559.950 202.800 ;
        RECT 561.150 202.800 562.050 204.900 ;
        RECT 562.950 204.300 570.450 205.500 ;
        RECT 562.950 203.700 564.750 204.300 ;
        RECT 577.050 203.400 578.850 215.250 ;
        RECT 608.550 209.400 610.350 215.250 ;
        RECT 611.550 209.400 613.350 215.250 ;
        RECT 567.750 202.800 578.850 203.400 ;
        RECT 561.150 202.200 578.850 202.800 ;
        RECT 561.150 201.900 569.550 202.200 ;
        RECT 567.750 201.600 569.550 201.900 ;
        RECT 559.050 196.050 562.050 198.150 ;
        RECT 565.950 197.100 568.050 198.150 ;
        RECT 565.950 196.050 573.900 197.100 ;
        RECT 547.950 195.750 550.050 196.050 ;
        RECT 547.950 193.950 551.850 195.750 ;
        RECT 533.250 191.700 537.000 192.750 ;
        RECT 545.550 191.850 550.050 193.950 ;
        RECT 559.050 192.000 559.950 196.050 ;
        RECT 572.100 195.300 573.900 196.050 ;
        RECT 575.100 195.150 576.900 196.950 ;
        RECT 569.100 194.400 570.900 195.000 ;
        RECT 575.100 194.400 576.000 195.150 ;
        RECT 569.100 193.200 576.000 194.400 ;
        RECT 569.100 192.000 570.150 193.200 ;
        RECT 533.250 189.600 534.450 191.700 ;
        RECT 457.650 183.750 459.450 186.600 ;
        RECT 460.650 183.750 462.450 186.600 ;
        RECT 463.650 183.750 465.450 186.600 ;
        RECT 494.550 183.750 496.350 186.600 ;
        RECT 497.550 183.750 499.350 186.600 ;
        RECT 532.650 183.750 534.450 189.600 ;
        RECT 535.650 188.700 543.450 190.050 ;
        RECT 535.650 183.750 537.450 188.700 ;
        RECT 538.650 183.750 540.450 187.800 ;
        RECT 541.650 183.750 543.450 188.700 ;
        RECT 545.550 189.600 546.750 191.850 ;
        RECT 559.050 191.100 570.150 192.000 ;
        RECT 559.050 190.800 559.950 191.100 ;
        RECT 545.550 183.750 547.350 189.600 ;
        RECT 550.950 188.700 553.050 189.600 ;
        RECT 558.150 189.000 559.950 190.800 ;
        RECT 569.100 190.200 570.150 191.100 ;
        RECT 565.350 189.450 567.150 190.200 ;
        RECT 550.950 187.500 554.700 188.700 ;
        RECT 553.650 186.600 554.700 187.500 ;
        RECT 562.200 188.400 567.150 189.450 ;
        RECT 568.650 188.400 570.450 190.200 ;
        RECT 577.950 189.600 578.850 202.200 ;
        RECT 611.400 196.950 612.600 209.400 ;
        RECT 641.550 203.400 643.350 215.250 ;
        RECT 645.750 203.400 647.550 215.250 ;
        RECT 682.650 203.400 684.450 215.250 ;
        RECT 685.650 204.300 687.450 215.250 ;
        RECT 688.650 205.200 690.450 215.250 ;
        RECT 691.650 204.300 693.450 215.250 ;
        RECT 722.550 209.400 724.350 215.250 ;
        RECT 725.550 209.400 727.350 215.250 ;
        RECT 685.650 203.400 693.450 204.300 ;
        RECT 645.000 202.350 647.550 203.400 ;
        RECT 641.100 198.150 642.900 199.950 ;
        RECT 608.100 195.150 609.900 196.950 ;
        RECT 607.950 193.050 610.050 195.150 ;
        RECT 610.950 194.850 613.050 196.950 ;
        RECT 640.950 196.050 643.050 198.150 ;
        RECT 645.000 195.150 646.050 202.350 ;
        RECT 647.100 198.150 648.900 199.950 ;
        RECT 683.100 198.150 684.300 203.400 ;
        RECT 722.100 198.150 723.900 199.950 ;
        RECT 646.950 196.050 649.050 198.150 ;
        RECT 682.950 196.050 685.050 198.150 ;
        RECT 562.200 186.600 563.250 188.400 ;
        RECT 571.950 187.500 574.050 189.600 ;
        RECT 571.950 186.600 573.000 187.500 ;
        RECT 548.850 183.750 550.650 186.600 ;
        RECT 553.350 183.750 555.150 186.600 ;
        RECT 557.550 183.750 559.350 186.600 ;
        RECT 561.450 183.750 563.250 186.600 ;
        RECT 564.750 183.750 566.550 186.600 ;
        RECT 569.250 185.700 573.000 186.600 ;
        RECT 569.250 183.750 571.050 185.700 ;
        RECT 574.050 183.750 575.850 186.600 ;
        RECT 577.050 183.750 578.850 189.600 ;
        RECT 611.400 186.600 612.600 194.850 ;
        RECT 643.950 193.050 646.050 195.150 ;
        RECT 645.000 186.600 646.050 193.050 ;
        RECT 683.100 189.600 684.300 196.050 ;
        RECT 685.950 194.850 688.050 196.950 ;
        RECT 689.100 195.150 690.900 196.950 ;
        RECT 686.100 193.050 687.900 194.850 ;
        RECT 688.950 193.050 691.050 195.150 ;
        RECT 691.950 194.850 694.050 196.950 ;
        RECT 721.950 196.050 724.050 198.150 ;
        RECT 692.100 193.050 693.900 194.850 ;
        RECT 725.700 192.300 726.900 209.400 ;
        RECT 729.150 203.400 730.950 215.250 ;
        RECT 732.150 203.400 733.950 215.250 ;
        RECT 727.950 197.850 730.050 199.950 ;
        RECT 732.150 198.150 733.350 203.400 ;
        RECT 728.100 196.050 729.900 197.850 ;
        RECT 730.950 196.050 733.350 198.150 ;
        RECT 722.550 191.100 730.050 192.300 ;
        RECT 683.100 187.950 688.800 189.600 ;
        RECT 608.550 183.750 610.350 186.600 ;
        RECT 611.550 183.750 613.350 186.600 ;
        RECT 641.550 183.750 643.350 186.600 ;
        RECT 644.550 183.750 646.350 186.600 ;
        RECT 647.550 183.750 649.350 186.600 ;
        RECT 683.700 183.750 685.500 186.600 ;
        RECT 687.000 183.750 688.800 187.950 ;
        RECT 691.200 183.750 693.000 189.600 ;
        RECT 722.550 183.750 724.350 191.100 ;
        RECT 728.250 190.500 730.050 191.100 ;
        RECT 732.150 189.600 733.350 196.050 ;
        RECT 727.050 183.750 728.850 189.600 ;
        RECT 730.050 188.100 733.350 189.600 ;
        RECT 730.050 183.750 731.850 188.100 ;
        RECT 33.150 174.900 34.950 179.250 ;
        RECT 31.650 173.400 34.950 174.900 ;
        RECT 36.150 173.400 37.950 179.250 ;
        RECT 31.650 166.950 32.850 173.400 ;
        RECT 34.950 171.900 36.750 172.500 ;
        RECT 40.650 171.900 42.450 179.250 ;
        RECT 74.700 176.400 76.500 179.250 ;
        RECT 78.000 175.050 79.800 179.250 ;
        RECT 34.950 170.700 42.450 171.900 ;
        RECT 74.100 173.400 79.800 175.050 ;
        RECT 82.200 173.400 84.000 179.250 ;
        RECT 31.650 164.850 34.050 166.950 ;
        RECT 35.100 165.150 36.900 166.950 ;
        RECT 31.650 159.600 32.850 164.850 ;
        RECT 34.950 163.050 37.050 165.150 ;
        RECT 31.050 147.750 32.850 159.600 ;
        RECT 34.050 147.750 35.850 159.600 ;
        RECT 38.100 153.600 39.300 170.700 ;
        RECT 74.100 166.950 75.300 173.400 ;
        RECT 113.550 171.900 115.350 179.250 ;
        RECT 118.050 173.400 119.850 179.250 ;
        RECT 121.050 174.900 122.850 179.250 ;
        RECT 158.700 176.400 160.500 179.250 ;
        RECT 162.000 175.050 163.800 179.250 ;
        RECT 121.050 173.400 124.350 174.900 ;
        RECT 119.250 171.900 121.050 172.500 ;
        RECT 113.550 170.700 121.050 171.900 ;
        RECT 77.100 168.150 78.900 169.950 ;
        RECT 40.950 164.850 43.050 166.950 ;
        RECT 73.950 164.850 76.050 166.950 ;
        RECT 76.950 166.050 79.050 168.150 ;
        RECT 79.950 167.850 82.050 169.950 ;
        RECT 83.100 168.150 84.900 169.950 ;
        RECT 80.100 166.050 81.900 167.850 ;
        RECT 82.950 166.050 85.050 168.150 ;
        RECT 112.950 164.850 115.050 166.950 ;
        RECT 41.100 163.050 42.900 164.850 ;
        RECT 74.100 159.600 75.300 164.850 ;
        RECT 113.100 163.050 114.900 164.850 ;
        RECT 37.650 147.750 39.450 153.600 ;
        RECT 40.650 147.750 42.450 153.600 ;
        RECT 73.650 147.750 75.450 159.600 ;
        RECT 76.650 158.700 84.450 159.600 ;
        RECT 76.650 147.750 78.450 158.700 ;
        RECT 79.650 147.750 81.450 157.800 ;
        RECT 82.650 147.750 84.450 158.700 ;
        RECT 116.700 153.600 117.900 170.700 ;
        RECT 123.150 166.950 124.350 173.400 ;
        RECT 158.100 173.400 163.800 175.050 ;
        RECT 166.200 173.400 168.000 179.250 ;
        RECT 198.000 173.400 199.800 179.250 ;
        RECT 202.200 175.050 204.000 179.250 ;
        RECT 205.500 176.400 207.300 179.250 ;
        RECT 239.550 176.400 241.350 179.250 ;
        RECT 242.550 176.400 244.350 179.250 ;
        RECT 245.550 176.400 247.350 179.250 ;
        RECT 202.200 173.400 207.900 175.050 ;
        RECT 158.100 166.950 159.300 173.400 ;
        RECT 161.100 168.150 162.900 169.950 ;
        RECT 119.100 165.150 120.900 166.950 ;
        RECT 118.950 163.050 121.050 165.150 ;
        RECT 121.950 164.850 124.350 166.950 ;
        RECT 157.950 164.850 160.050 166.950 ;
        RECT 160.950 166.050 163.050 168.150 ;
        RECT 163.950 167.850 166.050 169.950 ;
        RECT 167.100 168.150 168.900 169.950 ;
        RECT 197.100 168.150 198.900 169.950 ;
        RECT 164.100 166.050 165.900 167.850 ;
        RECT 166.950 166.050 169.050 168.150 ;
        RECT 196.950 166.050 199.050 168.150 ;
        RECT 199.950 167.850 202.050 169.950 ;
        RECT 203.100 168.150 204.900 169.950 ;
        RECT 200.100 166.050 201.900 167.850 ;
        RECT 202.950 166.050 205.050 168.150 ;
        RECT 206.700 166.950 207.900 173.400 ;
        RECT 243.450 172.200 244.350 176.400 ;
        RECT 248.550 173.400 250.350 179.250 ;
        RECT 280.650 173.400 282.450 179.250 ;
        RECT 283.650 173.400 285.450 179.250 ;
        RECT 286.650 173.400 288.450 179.250 ;
        RECT 289.650 173.400 291.450 179.250 ;
        RECT 292.650 173.400 294.450 179.250 ;
        RECT 323.550 176.400 325.350 179.250 ;
        RECT 243.450 171.300 246.750 172.200 ;
        RECT 244.950 170.400 246.750 171.300 ;
        RECT 238.950 167.850 241.050 169.950 ;
        RECT 205.950 164.850 208.050 166.950 ;
        RECT 239.100 166.050 240.900 167.850 ;
        RECT 241.950 164.850 244.050 166.950 ;
        RECT 123.150 159.600 124.350 164.850 ;
        RECT 158.100 159.600 159.300 164.850 ;
        RECT 206.700 159.600 207.900 164.850 ;
        RECT 242.100 163.050 243.900 164.850 ;
        RECT 245.700 162.150 246.600 170.400 ;
        RECT 249.000 168.150 250.050 173.400 ;
        RECT 247.950 166.050 250.050 168.150 ;
        RECT 284.250 172.500 285.450 173.400 ;
        RECT 290.250 172.500 291.450 173.400 ;
        RECT 284.250 171.300 291.450 172.500 ;
        RECT 324.150 172.500 325.350 176.400 ;
        RECT 326.850 173.400 328.650 179.250 ;
        RECT 329.850 173.400 331.650 179.250 ;
        RECT 364.650 173.400 366.450 179.250 ;
        RECT 324.150 171.600 329.250 172.500 ;
        RECT 284.250 166.950 285.450 171.300 ;
        RECT 327.000 170.700 329.250 171.600 ;
        RECT 244.950 162.000 246.750 162.150 ;
        RECT 239.550 160.800 246.750 162.000 ;
        RECT 239.550 159.600 240.750 160.800 ;
        RECT 244.950 160.350 246.750 160.800 ;
        RECT 113.550 147.750 115.350 153.600 ;
        RECT 116.550 147.750 118.350 153.600 ;
        RECT 120.150 147.750 121.950 159.600 ;
        RECT 123.150 147.750 124.950 159.600 ;
        RECT 157.650 147.750 159.450 159.600 ;
        RECT 160.650 158.700 168.450 159.600 ;
        RECT 160.650 147.750 162.450 158.700 ;
        RECT 163.650 147.750 165.450 157.800 ;
        RECT 166.650 147.750 168.450 158.700 ;
        RECT 197.550 158.700 205.350 159.600 ;
        RECT 197.550 147.750 199.350 158.700 ;
        RECT 200.550 147.750 202.350 157.800 ;
        RECT 203.550 147.750 205.350 158.700 ;
        RECT 206.550 147.750 208.350 159.600 ;
        RECT 239.550 147.750 241.350 159.600 ;
        RECT 248.100 159.450 249.450 166.050 ;
        RECT 283.950 164.850 286.050 166.950 ;
        RECT 289.950 164.850 292.050 166.950 ;
        RECT 322.950 164.850 325.050 166.950 ;
        RECT 284.250 161.400 285.450 164.850 ;
        RECT 290.100 163.050 291.900 164.850 ;
        RECT 323.100 163.050 324.900 164.850 ;
        RECT 327.000 162.300 328.050 170.700 ;
        RECT 330.150 166.950 331.350 173.400 ;
        RECT 365.250 171.300 366.450 173.400 ;
        RECT 367.650 174.300 369.450 179.250 ;
        RECT 370.650 175.200 372.450 179.250 ;
        RECT 373.650 174.300 375.450 179.250 ;
        RECT 406.650 176.400 408.450 179.250 ;
        RECT 409.650 176.400 411.450 179.250 ;
        RECT 412.650 176.400 414.450 179.250 ;
        RECT 367.650 172.950 375.450 174.300 ;
        RECT 365.250 170.250 369.000 171.300 ;
        RECT 328.950 164.850 331.350 166.950 ;
        RECT 367.950 166.950 369.150 170.250 ;
        RECT 409.950 169.950 411.000 176.400 ;
        RECT 444.000 173.400 445.800 179.250 ;
        RECT 448.200 175.050 450.000 179.250 ;
        RECT 451.500 176.400 453.300 179.250 ;
        RECT 448.200 173.400 453.900 175.050 ;
        RECT 371.100 168.150 372.900 169.950 ;
        RECT 367.950 164.850 370.050 166.950 ;
        RECT 370.950 166.050 373.050 168.150 ;
        RECT 409.950 167.850 412.050 169.950 ;
        RECT 443.100 168.150 444.900 169.950 ;
        RECT 373.950 164.850 376.050 166.950 ;
        RECT 406.950 164.850 409.050 166.950 ;
        RECT 327.000 161.400 329.250 162.300 ;
        RECT 284.250 160.500 291.450 161.400 ;
        RECT 284.250 159.600 285.450 160.500 ;
        RECT 244.050 147.750 245.850 159.450 ;
        RECT 247.050 158.100 249.450 159.450 ;
        RECT 247.050 147.750 248.850 158.100 ;
        RECT 280.650 147.750 282.450 159.600 ;
        RECT 283.650 147.750 285.450 159.600 ;
        RECT 286.650 147.750 288.450 159.600 ;
        RECT 289.650 147.750 291.450 160.500 ;
        RECT 323.550 160.500 329.250 161.400 ;
        RECT 292.650 147.750 294.450 159.600 ;
        RECT 323.550 153.600 324.750 160.500 ;
        RECT 330.150 159.600 331.350 164.850 ;
        RECT 364.950 161.850 367.050 163.950 ;
        RECT 365.250 160.050 367.050 161.850 ;
        RECT 368.850 159.600 370.050 164.850 ;
        RECT 374.100 163.050 375.900 164.850 ;
        RECT 407.100 163.050 408.900 164.850 ;
        RECT 409.950 160.650 411.000 167.850 ;
        RECT 412.950 164.850 415.050 166.950 ;
        RECT 442.950 166.050 445.050 168.150 ;
        RECT 445.950 167.850 448.050 169.950 ;
        RECT 449.100 168.150 450.900 169.950 ;
        RECT 446.100 166.050 447.900 167.850 ;
        RECT 448.950 166.050 451.050 168.150 ;
        RECT 452.700 166.950 453.900 173.400 ;
        RECT 459.150 173.400 460.950 179.250 ;
        RECT 462.150 176.400 463.950 179.250 ;
        RECT 466.950 177.300 468.750 179.250 ;
        RECT 465.000 176.400 468.750 177.300 ;
        RECT 471.450 176.400 473.250 179.250 ;
        RECT 474.750 176.400 476.550 179.250 ;
        RECT 478.650 176.400 480.450 179.250 ;
        RECT 482.850 176.400 484.650 179.250 ;
        RECT 487.350 176.400 489.150 179.250 ;
        RECT 465.000 175.500 466.050 176.400 ;
        RECT 463.950 173.400 466.050 175.500 ;
        RECT 474.750 174.600 475.800 176.400 ;
        RECT 451.950 164.850 454.050 166.950 ;
        RECT 413.100 163.050 414.900 164.850 ;
        RECT 408.450 159.600 411.000 160.650 ;
        RECT 452.700 159.600 453.900 164.850 ;
        RECT 459.150 160.800 460.050 173.400 ;
        RECT 467.550 172.800 469.350 174.600 ;
        RECT 470.850 173.550 475.800 174.600 ;
        RECT 483.300 175.500 484.350 176.400 ;
        RECT 483.300 174.300 487.050 175.500 ;
        RECT 470.850 172.800 472.650 173.550 ;
        RECT 467.850 171.900 468.900 172.800 ;
        RECT 478.050 172.200 479.850 174.000 ;
        RECT 484.950 173.400 487.050 174.300 ;
        RECT 490.650 173.400 492.450 179.250 ;
        RECT 478.050 171.900 478.950 172.200 ;
        RECT 467.850 171.000 478.950 171.900 ;
        RECT 491.250 171.150 492.450 173.400 ;
        RECT 518.550 174.300 520.350 179.250 ;
        RECT 521.550 175.200 523.350 179.250 ;
        RECT 524.550 174.300 526.350 179.250 ;
        RECT 518.550 172.950 526.350 174.300 ;
        RECT 527.550 173.400 529.350 179.250 ;
        RECT 559.650 173.400 561.450 179.250 ;
        RECT 527.550 171.300 528.750 173.400 ;
        RECT 467.850 169.800 468.900 171.000 ;
        RECT 462.000 168.600 468.900 169.800 ;
        RECT 462.000 167.850 462.900 168.600 ;
        RECT 467.100 168.000 468.900 168.600 ;
        RECT 461.100 166.050 462.900 167.850 ;
        RECT 464.100 166.950 465.900 167.700 ;
        RECT 478.050 166.950 478.950 171.000 ;
        RECT 487.950 169.050 492.450 171.150 ;
        RECT 525.000 170.250 528.750 171.300 ;
        RECT 560.250 171.300 561.450 173.400 ;
        RECT 562.650 174.300 564.450 179.250 ;
        RECT 565.650 175.200 567.450 179.250 ;
        RECT 568.650 174.300 570.450 179.250 ;
        RECT 602.700 176.400 604.500 179.250 ;
        RECT 606.000 175.050 607.800 179.250 ;
        RECT 562.650 172.950 570.450 174.300 ;
        RECT 602.100 173.400 607.800 175.050 ;
        RECT 610.200 173.400 612.000 179.250 ;
        RECT 644.700 176.400 646.500 179.250 ;
        RECT 648.000 175.050 649.800 179.250 ;
        RECT 644.100 173.400 649.800 175.050 ;
        RECT 652.200 173.400 654.000 179.250 ;
        RECT 683.550 176.400 685.350 179.250 ;
        RECT 686.550 176.400 688.350 179.250 ;
        RECT 689.550 176.400 691.350 179.250 ;
        RECT 560.250 170.250 564.000 171.300 ;
        RECT 486.150 167.250 490.050 169.050 ;
        RECT 487.950 166.950 490.050 167.250 ;
        RECT 464.100 165.900 472.050 166.950 ;
        RECT 469.950 164.850 472.050 165.900 ;
        RECT 475.950 164.850 478.950 166.950 ;
        RECT 468.450 161.100 470.250 161.400 ;
        RECT 468.450 160.800 476.850 161.100 ;
        RECT 459.150 160.200 476.850 160.800 ;
        RECT 459.150 159.600 470.250 160.200 ;
        RECT 323.550 147.750 325.350 153.600 ;
        RECT 326.850 147.750 328.650 159.600 ;
        RECT 329.850 147.750 331.650 159.600 ;
        RECT 365.400 147.750 367.200 153.600 ;
        RECT 368.700 147.750 370.500 159.600 ;
        RECT 372.900 147.750 374.700 159.600 ;
        RECT 408.450 147.750 410.250 159.600 ;
        RECT 412.650 147.750 414.450 159.600 ;
        RECT 443.550 158.700 451.350 159.600 ;
        RECT 443.550 147.750 445.350 158.700 ;
        RECT 446.550 147.750 448.350 157.800 ;
        RECT 449.550 147.750 451.350 158.700 ;
        RECT 452.550 147.750 454.350 159.600 ;
        RECT 459.150 147.750 460.950 159.600 ;
        RECT 473.250 158.700 475.050 159.300 ;
        RECT 467.550 157.500 475.050 158.700 ;
        RECT 475.950 158.100 476.850 160.200 ;
        RECT 478.050 160.200 478.950 164.850 ;
        RECT 488.250 161.400 490.050 163.200 ;
        RECT 484.950 160.200 489.150 161.400 ;
        RECT 478.050 159.300 484.050 160.200 ;
        RECT 484.950 159.300 487.050 160.200 ;
        RECT 491.250 159.600 492.450 169.050 ;
        RECT 521.100 168.150 522.900 169.950 ;
        RECT 517.950 164.850 520.050 166.950 ;
        RECT 520.950 166.050 523.050 168.150 ;
        RECT 524.850 166.950 526.050 170.250 ;
        RECT 523.950 164.850 526.050 166.950 ;
        RECT 562.950 166.950 564.150 170.250 ;
        RECT 566.100 168.150 567.900 169.950 ;
        RECT 562.950 164.850 565.050 166.950 ;
        RECT 565.950 166.050 568.050 168.150 ;
        RECT 602.100 166.950 603.300 173.400 ;
        RECT 605.100 168.150 606.900 169.950 ;
        RECT 568.950 164.850 571.050 166.950 ;
        RECT 601.950 164.850 604.050 166.950 ;
        RECT 604.950 166.050 607.050 168.150 ;
        RECT 607.950 167.850 610.050 169.950 ;
        RECT 611.100 168.150 612.900 169.950 ;
        RECT 608.100 166.050 609.900 167.850 ;
        RECT 610.950 166.050 613.050 168.150 ;
        RECT 644.100 166.950 645.300 173.400 ;
        RECT 687.450 172.200 688.350 176.400 ;
        RECT 692.550 173.400 694.350 179.250 ;
        RECT 687.450 171.300 690.750 172.200 ;
        RECT 688.950 170.400 690.750 171.300 ;
        RECT 647.100 168.150 648.900 169.950 ;
        RECT 643.950 164.850 646.050 166.950 ;
        RECT 646.950 166.050 649.050 168.150 ;
        RECT 649.950 167.850 652.050 169.950 ;
        RECT 653.100 168.150 654.900 169.950 ;
        RECT 650.100 166.050 651.900 167.850 ;
        RECT 652.950 166.050 655.050 168.150 ;
        RECT 682.950 167.850 685.050 169.950 ;
        RECT 683.100 166.050 684.900 167.850 ;
        RECT 685.950 164.850 688.050 166.950 ;
        RECT 518.100 163.050 519.900 164.850 ;
        RECT 523.950 159.600 525.150 164.850 ;
        RECT 526.950 161.850 529.050 163.950 ;
        RECT 559.950 161.850 562.050 163.950 ;
        RECT 526.950 160.050 528.750 161.850 ;
        RECT 560.250 160.050 562.050 161.850 ;
        RECT 563.850 159.600 565.050 164.850 ;
        RECT 569.100 163.050 570.900 164.850 ;
        RECT 602.100 159.600 603.300 164.850 ;
        RECT 644.100 159.600 645.300 164.850 ;
        RECT 686.100 163.050 687.900 164.850 ;
        RECT 689.700 162.150 690.600 170.400 ;
        RECT 693.000 168.150 694.050 173.400 ;
        RECT 725.550 171.900 727.350 179.250 ;
        RECT 730.050 173.400 731.850 179.250 ;
        RECT 733.050 174.900 734.850 179.250 ;
        RECT 733.050 173.400 736.350 174.900 ;
        RECT 731.250 171.900 733.050 172.500 ;
        RECT 725.550 170.700 733.050 171.900 ;
        RECT 691.950 166.050 694.050 168.150 ;
        RECT 688.950 162.000 690.750 162.150 ;
        RECT 683.550 160.800 690.750 162.000 ;
        RECT 683.550 159.600 684.750 160.800 ;
        RECT 688.950 160.350 690.750 160.800 ;
        RECT 483.150 158.400 484.050 159.300 ;
        RECT 480.450 158.100 482.250 158.400 ;
        RECT 467.550 156.600 468.750 157.500 ;
        RECT 475.950 157.200 482.250 158.100 ;
        RECT 480.450 156.600 482.250 157.200 ;
        RECT 483.150 156.600 485.850 158.400 ;
        RECT 463.950 154.500 468.750 156.600 ;
        RECT 471.150 154.500 478.050 156.300 ;
        RECT 467.550 153.600 468.750 154.500 ;
        RECT 462.150 147.750 463.950 153.600 ;
        RECT 467.250 147.750 469.050 153.600 ;
        RECT 472.050 147.750 473.850 153.600 ;
        RECT 475.050 147.750 476.850 154.500 ;
        RECT 483.150 153.600 487.050 155.700 ;
        RECT 478.950 147.750 480.750 153.600 ;
        RECT 483.150 147.750 484.950 153.600 ;
        RECT 487.650 147.750 489.450 150.600 ;
        RECT 490.650 147.750 492.450 159.600 ;
        RECT 519.300 147.750 521.100 159.600 ;
        RECT 523.500 147.750 525.300 159.600 ;
        RECT 526.800 147.750 528.600 153.600 ;
        RECT 560.400 147.750 562.200 153.600 ;
        RECT 563.700 147.750 565.500 159.600 ;
        RECT 567.900 147.750 569.700 159.600 ;
        RECT 601.650 147.750 603.450 159.600 ;
        RECT 604.650 158.700 612.450 159.600 ;
        RECT 604.650 147.750 606.450 158.700 ;
        RECT 607.650 147.750 609.450 157.800 ;
        RECT 610.650 147.750 612.450 158.700 ;
        RECT 643.650 147.750 645.450 159.600 ;
        RECT 646.650 158.700 654.450 159.600 ;
        RECT 646.650 147.750 648.450 158.700 ;
        RECT 649.650 147.750 651.450 157.800 ;
        RECT 652.650 147.750 654.450 158.700 ;
        RECT 683.550 147.750 685.350 159.600 ;
        RECT 692.100 159.450 693.450 166.050 ;
        RECT 724.950 164.850 727.050 166.950 ;
        RECT 725.100 163.050 726.900 164.850 ;
        RECT 688.050 147.750 689.850 159.450 ;
        RECT 691.050 158.100 693.450 159.450 ;
        RECT 691.050 147.750 692.850 158.100 ;
        RECT 728.700 153.600 729.900 170.700 ;
        RECT 735.150 166.950 736.350 173.400 ;
        RECT 731.100 165.150 732.900 166.950 ;
        RECT 730.950 163.050 733.050 165.150 ;
        RECT 733.950 164.850 736.350 166.950 ;
        RECT 735.150 159.600 736.350 164.850 ;
        RECT 725.550 147.750 727.350 153.600 ;
        RECT 728.550 147.750 730.350 153.600 ;
        RECT 732.150 147.750 733.950 159.600 ;
        RECT 735.150 147.750 736.950 159.600 ;
        RECT 33.450 131.400 35.250 143.250 ;
        RECT 37.650 131.400 39.450 143.250 ;
        RECT 70.650 137.400 72.450 143.250 ;
        RECT 73.650 137.400 75.450 143.250 ;
        RECT 33.450 130.350 36.000 131.400 ;
        RECT 32.100 126.150 33.900 127.950 ;
        RECT 31.950 124.050 34.050 126.150 ;
        RECT 34.950 123.150 36.000 130.350 ;
        RECT 38.100 126.150 39.900 127.950 ;
        RECT 37.950 124.050 40.050 126.150 ;
        RECT 71.400 124.950 72.600 137.400 ;
        RECT 102.300 131.400 104.100 143.250 ;
        RECT 106.500 131.400 108.300 143.250 ;
        RECT 109.800 137.400 111.600 143.250 ;
        RECT 141.300 131.400 143.100 143.250 ;
        RECT 145.500 131.400 147.300 143.250 ;
        RECT 148.800 137.400 150.600 143.250 ;
        RECT 184.650 137.400 186.450 143.250 ;
        RECT 187.650 137.400 189.450 143.250 ;
        RECT 101.100 126.150 102.900 127.950 ;
        RECT 106.950 126.150 108.150 131.400 ;
        RECT 109.950 129.150 111.750 130.950 ;
        RECT 109.950 127.050 112.050 129.150 ;
        RECT 140.100 126.150 141.900 127.950 ;
        RECT 145.950 126.150 147.150 131.400 ;
        RECT 148.950 129.150 150.750 130.950 ;
        RECT 148.950 127.050 151.050 129.150 ;
        RECT 34.950 121.050 37.050 123.150 ;
        RECT 70.950 122.850 73.050 124.950 ;
        RECT 74.100 123.150 75.900 124.950 ;
        RECT 100.950 124.050 103.050 126.150 ;
        RECT 34.950 114.600 36.000 121.050 ;
        RECT 71.400 114.600 72.600 122.850 ;
        RECT 73.950 121.050 76.050 123.150 ;
        RECT 103.950 122.850 106.050 124.950 ;
        RECT 106.950 124.050 109.050 126.150 ;
        RECT 139.950 124.050 142.050 126.150 ;
        RECT 104.100 121.050 105.900 122.850 ;
        RECT 107.850 120.750 109.050 124.050 ;
        RECT 142.950 122.850 145.050 124.950 ;
        RECT 145.950 124.050 148.050 126.150 ;
        RECT 185.400 124.950 186.600 137.400 ;
        RECT 218.550 132.300 220.350 143.250 ;
        RECT 221.550 133.200 223.350 143.250 ;
        RECT 224.550 132.300 226.350 143.250 ;
        RECT 218.550 131.400 226.350 132.300 ;
        RECT 227.550 131.400 229.350 143.250 ;
        RECT 264.450 131.400 266.250 143.250 ;
        RECT 268.650 131.400 270.450 143.250 ;
        RECT 273.150 131.400 274.950 143.250 ;
        RECT 276.150 137.400 277.950 143.250 ;
        RECT 281.250 137.400 283.050 143.250 ;
        RECT 286.050 137.400 287.850 143.250 ;
        RECT 281.550 136.500 282.750 137.400 ;
        RECT 289.050 136.500 290.850 143.250 ;
        RECT 292.950 137.400 294.750 143.250 ;
        RECT 297.150 137.400 298.950 143.250 ;
        RECT 301.650 140.400 303.450 143.250 ;
        RECT 277.950 134.400 282.750 136.500 ;
        RECT 285.150 134.700 292.050 136.500 ;
        RECT 297.150 135.300 301.050 137.400 ;
        RECT 281.550 133.500 282.750 134.400 ;
        RECT 294.450 133.800 296.250 134.400 ;
        RECT 281.550 132.300 289.050 133.500 ;
        RECT 287.250 131.700 289.050 132.300 ;
        RECT 289.950 132.900 296.250 133.800 ;
        RECT 227.700 126.150 228.900 131.400 ;
        RECT 264.450 130.350 267.000 131.400 ;
        RECT 263.100 126.150 264.900 127.950 ;
        RECT 143.100 121.050 144.900 122.850 ;
        RECT 146.850 120.750 148.050 124.050 ;
        RECT 184.950 122.850 187.050 124.950 ;
        RECT 188.100 123.150 189.900 124.950 ;
        RECT 108.000 119.700 111.750 120.750 ;
        RECT 147.000 119.700 150.750 120.750 ;
        RECT 101.550 116.700 109.350 118.050 ;
        RECT 31.650 111.750 33.450 114.600 ;
        RECT 34.650 111.750 36.450 114.600 ;
        RECT 37.650 111.750 39.450 114.600 ;
        RECT 70.650 111.750 72.450 114.600 ;
        RECT 73.650 111.750 75.450 114.600 ;
        RECT 101.550 111.750 103.350 116.700 ;
        RECT 104.550 111.750 106.350 115.800 ;
        RECT 107.550 111.750 109.350 116.700 ;
        RECT 110.550 117.600 111.750 119.700 ;
        RECT 110.550 111.750 112.350 117.600 ;
        RECT 140.550 116.700 148.350 118.050 ;
        RECT 140.550 111.750 142.350 116.700 ;
        RECT 143.550 111.750 145.350 115.800 ;
        RECT 146.550 111.750 148.350 116.700 ;
        RECT 149.550 117.600 150.750 119.700 ;
        RECT 149.550 111.750 151.350 117.600 ;
        RECT 185.400 114.600 186.600 122.850 ;
        RECT 187.950 121.050 190.050 123.150 ;
        RECT 217.950 122.850 220.050 124.950 ;
        RECT 221.100 123.150 222.900 124.950 ;
        RECT 218.100 121.050 219.900 122.850 ;
        RECT 220.950 121.050 223.050 123.150 ;
        RECT 223.950 122.850 226.050 124.950 ;
        RECT 226.950 124.050 229.050 126.150 ;
        RECT 262.950 124.050 265.050 126.150 ;
        RECT 224.100 121.050 225.900 122.850 ;
        RECT 227.700 117.600 228.900 124.050 ;
        RECT 265.950 123.150 267.000 130.350 ;
        RECT 273.150 130.800 284.250 131.400 ;
        RECT 289.950 130.800 290.850 132.900 ;
        RECT 294.450 132.600 296.250 132.900 ;
        RECT 297.150 132.600 299.850 134.400 ;
        RECT 297.150 131.700 298.050 132.600 ;
        RECT 273.150 130.200 290.850 130.800 ;
        RECT 269.100 126.150 270.900 127.950 ;
        RECT 268.950 124.050 271.050 126.150 ;
        RECT 265.950 121.050 268.050 123.150 ;
        RECT 256.950 120.450 259.050 121.050 ;
        RECT 262.950 120.450 265.050 121.050 ;
        RECT 256.950 119.550 265.050 120.450 ;
        RECT 256.950 118.950 259.050 119.550 ;
        RECT 262.950 118.950 265.050 119.550 ;
        RECT 184.650 111.750 186.450 114.600 ;
        RECT 187.650 111.750 189.450 114.600 ;
        RECT 219.000 111.750 220.800 117.600 ;
        RECT 223.200 115.950 228.900 117.600 ;
        RECT 223.200 111.750 225.000 115.950 ;
        RECT 265.950 114.600 267.000 121.050 ;
        RECT 273.150 117.600 274.050 130.200 ;
        RECT 282.450 129.900 290.850 130.200 ;
        RECT 292.050 130.800 298.050 131.700 ;
        RECT 298.950 130.800 301.050 131.700 ;
        RECT 304.650 131.400 306.450 143.250 ;
        RECT 335.550 131.400 337.350 143.250 ;
        RECT 339.750 131.400 341.550 143.250 ;
        RECT 374.400 137.400 376.200 143.250 ;
        RECT 377.700 131.400 379.500 143.250 ;
        RECT 381.900 131.400 383.700 143.250 ;
        RECT 412.650 131.400 414.450 143.250 ;
        RECT 415.650 132.300 417.450 143.250 ;
        RECT 418.650 133.200 420.450 143.250 ;
        RECT 421.650 132.300 423.450 143.250 ;
        RECT 452.550 137.400 454.350 143.250 ;
        RECT 455.550 137.400 457.350 143.250 ;
        RECT 458.550 137.400 460.350 143.250 ;
        RECT 415.650 131.400 423.450 132.300 ;
        RECT 282.450 129.600 284.250 129.900 ;
        RECT 292.050 126.150 292.950 130.800 ;
        RECT 298.950 129.600 303.150 130.800 ;
        RECT 302.250 127.800 304.050 129.600 ;
        RECT 283.950 125.100 286.050 126.150 ;
        RECT 275.100 123.150 276.900 124.950 ;
        RECT 278.100 124.050 286.050 125.100 ;
        RECT 289.950 124.050 292.950 126.150 ;
        RECT 278.100 123.300 279.900 124.050 ;
        RECT 276.000 122.400 276.900 123.150 ;
        RECT 281.100 122.400 282.900 123.000 ;
        RECT 276.000 121.200 282.900 122.400 ;
        RECT 281.850 120.000 282.900 121.200 ;
        RECT 292.050 120.000 292.950 124.050 ;
        RECT 301.950 123.750 304.050 124.050 ;
        RECT 300.150 121.950 304.050 123.750 ;
        RECT 305.250 121.950 306.450 131.400 ;
        RECT 339.000 130.350 341.550 131.400 ;
        RECT 335.100 126.150 336.900 127.950 ;
        RECT 334.950 124.050 337.050 126.150 ;
        RECT 339.000 123.150 340.050 130.350 ;
        RECT 374.250 129.150 376.050 130.950 ;
        RECT 341.100 126.150 342.900 127.950 ;
        RECT 373.950 127.050 376.050 129.150 ;
        RECT 377.850 126.150 379.050 131.400 ;
        RECT 383.100 126.150 384.900 127.950 ;
        RECT 413.100 126.150 414.300 131.400 ;
        RECT 455.550 129.150 456.750 137.400 ;
        RECT 492.150 132.900 493.950 143.250 ;
        RECT 491.550 131.550 493.950 132.900 ;
        RECT 495.150 131.550 496.950 143.250 ;
        RECT 340.950 124.050 343.050 126.150 ;
        RECT 376.950 124.050 379.050 126.150 ;
        RECT 281.850 119.100 292.950 120.000 ;
        RECT 301.950 119.850 306.450 121.950 ;
        RECT 337.950 121.050 340.050 123.150 ;
        RECT 281.850 118.200 282.900 119.100 ;
        RECT 292.050 118.800 292.950 119.100 ;
        RECT 226.500 111.750 228.300 114.600 ;
        RECT 262.650 111.750 264.450 114.600 ;
        RECT 265.650 111.750 267.450 114.600 ;
        RECT 268.650 111.750 270.450 114.600 ;
        RECT 273.150 111.750 274.950 117.600 ;
        RECT 277.950 115.500 280.050 117.600 ;
        RECT 281.550 116.400 283.350 118.200 ;
        RECT 284.850 117.450 286.650 118.200 ;
        RECT 284.850 116.400 289.800 117.450 ;
        RECT 292.050 117.000 293.850 118.800 ;
        RECT 305.250 117.600 306.450 119.850 ;
        RECT 298.950 116.700 301.050 117.600 ;
        RECT 279.000 114.600 280.050 115.500 ;
        RECT 288.750 114.600 289.800 116.400 ;
        RECT 297.300 115.500 301.050 116.700 ;
        RECT 297.300 114.600 298.350 115.500 ;
        RECT 276.150 111.750 277.950 114.600 ;
        RECT 279.000 113.700 282.750 114.600 ;
        RECT 280.950 111.750 282.750 113.700 ;
        RECT 285.450 111.750 287.250 114.600 ;
        RECT 288.750 111.750 290.550 114.600 ;
        RECT 292.650 111.750 294.450 114.600 ;
        RECT 296.850 111.750 298.650 114.600 ;
        RECT 301.350 111.750 303.150 114.600 ;
        RECT 304.650 111.750 306.450 117.600 ;
        RECT 339.000 114.600 340.050 121.050 ;
        RECT 376.950 120.750 378.150 124.050 ;
        RECT 379.950 122.850 382.050 124.950 ;
        RECT 382.950 124.050 385.050 126.150 ;
        RECT 412.950 124.050 415.050 126.150 ;
        RECT 451.950 125.850 454.050 127.950 ;
        RECT 454.950 127.050 457.050 129.150 ;
        RECT 380.100 121.050 381.900 122.850 ;
        RECT 374.250 119.700 378.000 120.750 ;
        RECT 374.250 117.600 375.450 119.700 ;
        RECT 335.550 111.750 337.350 114.600 ;
        RECT 338.550 111.750 340.350 114.600 ;
        RECT 341.550 111.750 343.350 114.600 ;
        RECT 373.650 111.750 375.450 117.600 ;
        RECT 376.650 116.700 384.450 118.050 ;
        RECT 376.650 111.750 378.450 116.700 ;
        RECT 379.650 111.750 381.450 115.800 ;
        RECT 382.650 111.750 384.450 116.700 ;
        RECT 413.100 117.600 414.300 124.050 ;
        RECT 415.950 122.850 418.050 124.950 ;
        RECT 419.100 123.150 420.900 124.950 ;
        RECT 416.100 121.050 417.900 122.850 ;
        RECT 418.950 121.050 421.050 123.150 ;
        RECT 421.950 122.850 424.050 124.950 ;
        RECT 452.100 124.050 453.900 125.850 ;
        RECT 422.100 121.050 423.900 122.850 ;
        RECT 455.550 119.700 456.750 127.050 ;
        RECT 457.950 125.850 460.050 127.950 ;
        RECT 458.100 124.050 459.900 125.850 ;
        RECT 491.550 124.950 492.900 131.550 ;
        RECT 499.650 131.400 501.450 143.250 ;
        RECT 533.400 137.400 535.200 143.250 ;
        RECT 536.700 131.400 538.500 143.250 ;
        RECT 540.900 131.400 542.700 143.250 ;
        RECT 571.650 131.400 573.450 143.250 ;
        RECT 574.650 132.300 576.450 143.250 ;
        RECT 577.650 133.200 579.450 143.250 ;
        RECT 580.650 132.300 582.450 143.250 ;
        RECT 610.650 137.400 612.450 143.250 ;
        RECT 613.650 138.000 615.450 143.250 ;
        RECT 574.650 131.400 582.450 132.300 ;
        RECT 611.250 137.100 612.450 137.400 ;
        RECT 616.650 137.400 618.450 143.250 ;
        RECT 619.650 137.400 621.450 143.250 ;
        RECT 650.550 137.400 652.350 143.250 ;
        RECT 653.550 137.400 655.350 143.250 ;
        RECT 656.550 137.400 658.350 143.250 ;
        RECT 689.550 137.400 691.350 143.250 ;
        RECT 692.550 137.400 694.350 143.250 ;
        RECT 695.550 137.400 697.350 143.250 ;
        RECT 728.550 137.400 730.350 143.250 ;
        RECT 731.550 137.400 733.350 143.250 ;
        RECT 734.550 137.400 736.350 143.250 ;
        RECT 616.650 137.100 618.300 137.400 ;
        RECT 611.250 136.200 618.300 137.100 ;
        RECT 494.250 130.200 496.050 130.650 ;
        RECT 500.250 130.200 501.450 131.400 ;
        RECT 494.250 129.000 501.450 130.200 ;
        RECT 533.250 129.150 535.050 130.950 ;
        RECT 494.250 128.850 496.050 129.000 ;
        RECT 490.950 122.850 493.050 124.950 ;
        RECT 455.550 118.800 459.150 119.700 ;
        RECT 413.100 115.950 418.800 117.600 ;
        RECT 413.700 111.750 415.500 114.600 ;
        RECT 417.000 111.750 418.800 115.950 ;
        RECT 421.200 111.750 423.000 117.600 ;
        RECT 452.850 111.750 454.650 117.600 ;
        RECT 457.350 111.750 459.150 118.800 ;
        RECT 490.950 117.600 492.000 122.850 ;
        RECT 494.400 120.600 495.300 128.850 ;
        RECT 497.100 126.150 498.900 127.950 ;
        RECT 532.950 127.050 535.050 129.150 ;
        RECT 536.850 126.150 538.050 131.400 ;
        RECT 542.100 126.150 543.900 127.950 ;
        RECT 572.100 126.150 573.300 131.400 ;
        RECT 611.250 127.950 612.300 136.200 ;
        RECT 617.100 132.150 618.900 133.950 ;
        RECT 613.950 129.150 615.750 130.950 ;
        RECT 616.950 130.050 619.050 132.150 ;
        RECT 620.100 129.150 621.900 130.950 ;
        RECT 653.550 129.150 654.750 137.400 ;
        RECT 692.550 129.150 693.750 137.400 ;
        RECT 731.550 129.150 732.750 137.400 ;
        RECT 496.950 124.050 499.050 126.150 ;
        RECT 500.100 123.150 501.900 124.950 ;
        RECT 535.950 124.050 538.050 126.150 ;
        RECT 499.950 121.050 502.050 123.150 ;
        RECT 535.950 120.750 537.150 124.050 ;
        RECT 538.950 122.850 541.050 124.950 ;
        RECT 541.950 124.050 544.050 126.150 ;
        RECT 571.950 124.050 574.050 126.150 ;
        RECT 610.950 125.850 613.050 127.950 ;
        RECT 613.950 127.050 616.050 129.150 ;
        RECT 619.950 127.050 622.050 129.150 ;
        RECT 649.950 125.850 652.050 127.950 ;
        RECT 652.950 127.050 655.050 129.150 ;
        RECT 539.100 121.050 540.900 122.850 ;
        RECT 494.250 119.700 496.050 120.600 ;
        RECT 533.250 119.700 537.000 120.750 ;
        RECT 494.250 118.800 497.550 119.700 ;
        RECT 490.650 111.750 492.450 117.600 ;
        RECT 496.650 114.600 497.550 118.800 ;
        RECT 533.250 117.600 534.450 119.700 ;
        RECT 493.650 111.750 495.450 114.600 ;
        RECT 496.650 111.750 498.450 114.600 ;
        RECT 499.650 111.750 501.450 114.600 ;
        RECT 532.650 111.750 534.450 117.600 ;
        RECT 535.650 116.700 543.450 118.050 ;
        RECT 535.650 111.750 537.450 116.700 ;
        RECT 538.650 111.750 540.450 115.800 ;
        RECT 541.650 111.750 543.450 116.700 ;
        RECT 572.100 117.600 573.300 124.050 ;
        RECT 574.950 122.850 577.050 124.950 ;
        RECT 578.100 123.150 579.900 124.950 ;
        RECT 575.100 121.050 576.900 122.850 ;
        RECT 577.950 121.050 580.050 123.150 ;
        RECT 580.950 122.850 583.050 124.950 ;
        RECT 581.100 121.050 582.900 122.850 ;
        RECT 611.400 121.650 612.600 125.850 ;
        RECT 650.100 124.050 651.900 125.850 ;
        RECT 611.400 120.000 615.900 121.650 ;
        RECT 572.100 115.950 577.800 117.600 ;
        RECT 572.700 111.750 574.500 114.600 ;
        RECT 576.000 111.750 577.800 115.950 ;
        RECT 580.200 111.750 582.000 117.600 ;
        RECT 614.100 111.750 615.900 120.000 ;
        RECT 619.500 111.750 621.300 120.600 ;
        RECT 653.550 119.700 654.750 127.050 ;
        RECT 655.950 125.850 658.050 127.950 ;
        RECT 688.950 125.850 691.050 127.950 ;
        RECT 691.950 127.050 694.050 129.150 ;
        RECT 656.100 124.050 657.900 125.850 ;
        RECT 689.100 124.050 690.900 125.850 ;
        RECT 692.550 119.700 693.750 127.050 ;
        RECT 694.950 125.850 697.050 127.950 ;
        RECT 727.950 125.850 730.050 127.950 ;
        RECT 730.950 127.050 733.050 129.150 ;
        RECT 695.100 124.050 696.900 125.850 ;
        RECT 728.100 124.050 729.900 125.850 ;
        RECT 731.550 119.700 732.750 127.050 ;
        RECT 733.950 125.850 736.050 127.950 ;
        RECT 734.100 124.050 735.900 125.850 ;
        RECT 653.550 118.800 657.150 119.700 ;
        RECT 692.550 118.800 696.150 119.700 ;
        RECT 731.550 118.800 735.150 119.700 ;
        RECT 650.850 111.750 652.650 117.600 ;
        RECT 655.350 111.750 657.150 118.800 ;
        RECT 689.850 111.750 691.650 117.600 ;
        RECT 694.350 111.750 696.150 118.800 ;
        RECT 728.850 111.750 730.650 117.600 ;
        RECT 733.350 111.750 735.150 118.800 ;
        RECT 30.150 102.900 31.950 107.250 ;
        RECT 28.650 101.400 31.950 102.900 ;
        RECT 33.150 101.400 34.950 107.250 ;
        RECT 28.650 94.950 29.850 101.400 ;
        RECT 31.950 99.900 33.750 100.500 ;
        RECT 37.650 99.900 39.450 107.250 ;
        RECT 66.000 101.400 67.800 107.250 ;
        RECT 70.200 103.050 72.000 107.250 ;
        RECT 73.500 104.400 75.300 107.250 ;
        RECT 107.550 104.400 109.350 107.250 ;
        RECT 110.550 104.400 112.350 107.250 ;
        RECT 70.200 101.400 75.900 103.050 ;
        RECT 31.950 98.700 39.450 99.900 ;
        RECT 28.650 92.850 31.050 94.950 ;
        RECT 32.100 93.150 33.900 94.950 ;
        RECT 28.650 87.600 29.850 92.850 ;
        RECT 31.950 91.050 34.050 93.150 ;
        RECT 28.050 75.750 29.850 87.600 ;
        RECT 31.050 75.750 32.850 87.600 ;
        RECT 35.100 81.600 36.300 98.700 ;
        RECT 65.100 96.150 66.900 97.950 ;
        RECT 37.950 92.850 40.050 94.950 ;
        RECT 64.950 94.050 67.050 96.150 ;
        RECT 67.950 95.850 70.050 97.950 ;
        RECT 71.100 96.150 72.900 97.950 ;
        RECT 68.100 94.050 69.900 95.850 ;
        RECT 70.950 94.050 73.050 96.150 ;
        RECT 74.700 94.950 75.900 101.400 ;
        RECT 106.950 95.850 109.050 97.950 ;
        RECT 110.400 96.150 111.600 104.400 ;
        RECT 146.850 100.200 148.650 107.250 ;
        RECT 151.350 101.400 153.150 107.250 ;
        RECT 182.550 104.400 184.350 107.250 ;
        RECT 185.550 104.400 187.350 107.250 ;
        RECT 146.850 99.300 150.450 100.200 ;
        RECT 73.950 92.850 76.050 94.950 ;
        RECT 107.100 94.050 108.900 95.850 ;
        RECT 109.950 94.050 112.050 96.150 ;
        RECT 38.100 91.050 39.900 92.850 ;
        RECT 74.700 87.600 75.900 92.850 ;
        RECT 65.550 86.700 73.350 87.600 ;
        RECT 34.650 75.750 36.450 81.600 ;
        RECT 37.650 75.750 39.450 81.600 ;
        RECT 65.550 75.750 67.350 86.700 ;
        RECT 68.550 75.750 70.350 85.800 ;
        RECT 71.550 75.750 73.350 86.700 ;
        RECT 74.550 75.750 76.350 87.600 ;
        RECT 110.400 81.600 111.600 94.050 ;
        RECT 146.100 93.150 147.900 94.950 ;
        RECT 145.950 91.050 148.050 93.150 ;
        RECT 149.250 91.950 150.450 99.300 ;
        RECT 181.950 95.850 184.050 97.950 ;
        RECT 185.400 96.150 186.600 104.400 ;
        RECT 218.550 102.300 220.350 107.250 ;
        RECT 221.550 103.200 223.350 107.250 ;
        RECT 224.550 102.300 226.350 107.250 ;
        RECT 218.550 100.950 226.350 102.300 ;
        RECT 227.550 101.400 229.350 107.250 ;
        RECT 259.650 101.400 261.450 107.250 ;
        RECT 227.550 99.300 228.750 101.400 ;
        RECT 225.000 98.250 228.750 99.300 ;
        RECT 260.250 99.300 261.450 101.400 ;
        RECT 262.650 102.300 264.450 107.250 ;
        RECT 265.650 103.200 267.450 107.250 ;
        RECT 268.650 102.300 270.450 107.250 ;
        RECT 299.550 104.400 301.350 107.250 ;
        RECT 302.550 104.400 304.350 107.250 ;
        RECT 305.550 104.400 307.350 107.250 ;
        RECT 262.650 100.950 270.450 102.300 ;
        RECT 303.450 100.200 304.350 104.400 ;
        RECT 308.550 101.400 310.350 107.250 ;
        RECT 339.000 101.400 340.800 107.250 ;
        RECT 343.200 103.050 345.000 107.250 ;
        RECT 346.500 104.400 348.300 107.250 ;
        RECT 343.200 101.400 348.900 103.050 ;
        RECT 381.000 101.400 382.800 107.250 ;
        RECT 385.200 103.050 387.000 107.250 ;
        RECT 388.500 104.400 390.300 107.250 ;
        RECT 422.550 104.400 424.350 107.250 ;
        RECT 425.550 104.400 427.350 107.250 ;
        RECT 428.550 104.400 430.350 107.250 ;
        RECT 385.200 101.400 390.900 103.050 ;
        RECT 303.450 99.300 306.750 100.200 ;
        RECT 260.250 98.250 264.000 99.300 ;
        RECT 304.950 98.400 306.750 99.300 ;
        RECT 221.100 96.150 222.900 97.950 ;
        RECT 152.100 93.150 153.900 94.950 ;
        RECT 182.100 94.050 183.900 95.850 ;
        RECT 184.950 94.050 187.050 96.150 ;
        RECT 148.950 89.850 151.050 91.950 ;
        RECT 151.950 91.050 154.050 93.150 ;
        RECT 149.250 81.600 150.450 89.850 ;
        RECT 185.400 81.600 186.600 94.050 ;
        RECT 217.950 92.850 220.050 94.950 ;
        RECT 220.950 94.050 223.050 96.150 ;
        RECT 224.850 94.950 226.050 98.250 ;
        RECT 223.950 92.850 226.050 94.950 ;
        RECT 262.950 94.950 264.150 98.250 ;
        RECT 266.100 96.150 267.900 97.950 ;
        RECT 262.950 92.850 265.050 94.950 ;
        RECT 265.950 94.050 268.050 96.150 ;
        RECT 298.950 95.850 301.050 97.950 ;
        RECT 268.950 92.850 271.050 94.950 ;
        RECT 299.100 94.050 300.900 95.850 ;
        RECT 301.950 92.850 304.050 94.950 ;
        RECT 218.100 91.050 219.900 92.850 ;
        RECT 223.950 87.600 225.150 92.850 ;
        RECT 226.950 89.850 229.050 91.950 ;
        RECT 259.950 89.850 262.050 91.950 ;
        RECT 226.950 88.050 228.750 89.850 ;
        RECT 260.250 88.050 262.050 89.850 ;
        RECT 263.850 87.600 265.050 92.850 ;
        RECT 269.100 91.050 270.900 92.850 ;
        RECT 302.100 91.050 303.900 92.850 ;
        RECT 305.700 90.150 306.600 98.400 ;
        RECT 309.000 96.150 310.050 101.400 ;
        RECT 338.100 96.150 339.900 97.950 ;
        RECT 307.950 94.050 310.050 96.150 ;
        RECT 337.950 94.050 340.050 96.150 ;
        RECT 340.950 95.850 343.050 97.950 ;
        RECT 344.100 96.150 345.900 97.950 ;
        RECT 341.100 94.050 342.900 95.850 ;
        RECT 343.950 94.050 346.050 96.150 ;
        RECT 347.700 94.950 348.900 101.400 ;
        RECT 380.100 96.150 381.900 97.950 ;
        RECT 304.950 90.000 306.750 90.150 ;
        RECT 299.550 88.800 306.750 90.000 ;
        RECT 299.550 87.600 300.750 88.800 ;
        RECT 304.950 88.350 306.750 88.800 ;
        RECT 107.550 75.750 109.350 81.600 ;
        RECT 110.550 75.750 112.350 81.600 ;
        RECT 145.650 75.750 147.450 81.600 ;
        RECT 148.650 75.750 150.450 81.600 ;
        RECT 151.650 75.750 153.450 81.600 ;
        RECT 182.550 75.750 184.350 81.600 ;
        RECT 185.550 75.750 187.350 81.600 ;
        RECT 219.300 75.750 221.100 87.600 ;
        RECT 223.500 75.750 225.300 87.600 ;
        RECT 226.800 75.750 228.600 81.600 ;
        RECT 260.400 75.750 262.200 81.600 ;
        RECT 263.700 75.750 265.500 87.600 ;
        RECT 267.900 75.750 269.700 87.600 ;
        RECT 299.550 75.750 301.350 87.600 ;
        RECT 308.100 87.450 309.450 94.050 ;
        RECT 346.950 92.850 349.050 94.950 ;
        RECT 379.950 94.050 382.050 96.150 ;
        RECT 382.950 95.850 385.050 97.950 ;
        RECT 386.100 96.150 387.900 97.950 ;
        RECT 383.100 94.050 384.900 95.850 ;
        RECT 385.950 94.050 388.050 96.150 ;
        RECT 389.700 94.950 390.900 101.400 ;
        RECT 426.000 97.950 427.050 104.400 ;
        RECT 463.650 101.400 465.450 107.250 ;
        RECT 464.250 99.300 465.450 101.400 ;
        RECT 466.650 102.300 468.450 107.250 ;
        RECT 469.650 103.200 471.450 107.250 ;
        RECT 472.650 102.300 474.450 107.250 ;
        RECT 466.650 100.950 474.450 102.300 ;
        RECT 476.550 101.400 478.350 107.250 ;
        RECT 479.850 104.400 481.650 107.250 ;
        RECT 484.350 104.400 486.150 107.250 ;
        RECT 488.550 104.400 490.350 107.250 ;
        RECT 492.450 104.400 494.250 107.250 ;
        RECT 495.750 104.400 497.550 107.250 ;
        RECT 500.250 105.300 502.050 107.250 ;
        RECT 500.250 104.400 504.000 105.300 ;
        RECT 505.050 104.400 506.850 107.250 ;
        RECT 484.650 103.500 485.700 104.400 ;
        RECT 481.950 102.300 485.700 103.500 ;
        RECT 493.200 102.600 494.250 104.400 ;
        RECT 502.950 103.500 504.000 104.400 ;
        RECT 481.950 101.400 484.050 102.300 ;
        RECT 464.250 98.250 468.000 99.300 ;
        RECT 476.550 99.150 477.750 101.400 ;
        RECT 489.150 100.200 490.950 102.000 ;
        RECT 493.200 101.550 498.150 102.600 ;
        RECT 496.350 100.800 498.150 101.550 ;
        RECT 499.650 100.800 501.450 102.600 ;
        RECT 502.950 101.400 505.050 103.500 ;
        RECT 508.050 101.400 509.850 107.250 ;
        RECT 539.850 101.400 541.650 107.250 ;
        RECT 490.050 99.900 490.950 100.200 ;
        RECT 500.100 99.900 501.150 100.800 ;
        RECT 424.950 95.850 427.050 97.950 ;
        RECT 388.950 92.850 391.050 94.950 ;
        RECT 421.950 92.850 424.050 94.950 ;
        RECT 347.700 87.600 348.900 92.850 ;
        RECT 389.700 87.600 390.900 92.850 ;
        RECT 422.100 91.050 423.900 92.850 ;
        RECT 426.000 88.650 427.050 95.850 ;
        RECT 466.950 94.950 468.150 98.250 ;
        RECT 470.100 96.150 471.900 97.950 ;
        RECT 476.550 97.050 481.050 99.150 ;
        RECT 490.050 99.000 501.150 99.900 ;
        RECT 427.950 92.850 430.050 94.950 ;
        RECT 466.950 92.850 469.050 94.950 ;
        RECT 469.950 94.050 472.050 96.150 ;
        RECT 472.950 92.850 475.050 94.950 ;
        RECT 428.100 91.050 429.900 92.850 ;
        RECT 463.950 89.850 466.050 91.950 ;
        RECT 426.000 87.600 428.550 88.650 ;
        RECT 464.250 88.050 466.050 89.850 ;
        RECT 467.850 87.600 469.050 92.850 ;
        RECT 473.100 91.050 474.900 92.850 ;
        RECT 476.550 87.600 477.750 97.050 ;
        RECT 478.950 95.250 482.850 97.050 ;
        RECT 478.950 94.950 481.050 95.250 ;
        RECT 490.050 94.950 490.950 99.000 ;
        RECT 500.100 97.800 501.150 99.000 ;
        RECT 500.100 96.600 507.000 97.800 ;
        RECT 500.100 96.000 501.900 96.600 ;
        RECT 506.100 95.850 507.000 96.600 ;
        RECT 503.100 94.950 504.900 95.700 ;
        RECT 490.050 92.850 493.050 94.950 ;
        RECT 496.950 93.900 504.900 94.950 ;
        RECT 506.100 94.050 507.900 95.850 ;
        RECT 496.950 92.850 499.050 93.900 ;
        RECT 478.950 89.400 480.750 91.200 ;
        RECT 479.850 88.200 484.050 89.400 ;
        RECT 490.050 88.200 490.950 92.850 ;
        RECT 498.750 89.100 500.550 89.400 ;
        RECT 304.050 75.750 305.850 87.450 ;
        RECT 307.050 86.100 309.450 87.450 ;
        RECT 338.550 86.700 346.350 87.600 ;
        RECT 307.050 75.750 308.850 86.100 ;
        RECT 338.550 75.750 340.350 86.700 ;
        RECT 341.550 75.750 343.350 85.800 ;
        RECT 344.550 75.750 346.350 86.700 ;
        RECT 347.550 75.750 349.350 87.600 ;
        RECT 380.550 86.700 388.350 87.600 ;
        RECT 380.550 75.750 382.350 86.700 ;
        RECT 383.550 75.750 385.350 85.800 ;
        RECT 386.550 75.750 388.350 86.700 ;
        RECT 389.550 75.750 391.350 87.600 ;
        RECT 422.550 75.750 424.350 87.600 ;
        RECT 426.750 75.750 428.550 87.600 ;
        RECT 464.400 75.750 466.200 81.600 ;
        RECT 467.700 75.750 469.500 87.600 ;
        RECT 471.900 75.750 473.700 87.600 ;
        RECT 476.550 75.750 478.350 87.600 ;
        RECT 481.950 87.300 484.050 88.200 ;
        RECT 484.950 87.300 490.950 88.200 ;
        RECT 492.150 88.800 500.550 89.100 ;
        RECT 508.950 88.800 509.850 101.400 ;
        RECT 544.350 100.200 546.150 107.250 ;
        RECT 542.550 99.300 546.150 100.200 ;
        RECT 552.150 101.400 553.950 107.250 ;
        RECT 555.150 104.400 556.950 107.250 ;
        RECT 559.950 105.300 561.750 107.250 ;
        RECT 558.000 104.400 561.750 105.300 ;
        RECT 564.450 104.400 566.250 107.250 ;
        RECT 567.750 104.400 569.550 107.250 ;
        RECT 571.650 104.400 573.450 107.250 ;
        RECT 575.850 104.400 577.650 107.250 ;
        RECT 580.350 104.400 582.150 107.250 ;
        RECT 558.000 103.500 559.050 104.400 ;
        RECT 556.950 101.400 559.050 103.500 ;
        RECT 567.750 102.600 568.800 104.400 ;
        RECT 539.100 93.150 540.900 94.950 ;
        RECT 538.950 91.050 541.050 93.150 ;
        RECT 542.550 91.950 543.750 99.300 ;
        RECT 545.100 93.150 546.900 94.950 ;
        RECT 541.950 89.850 544.050 91.950 ;
        RECT 544.950 91.050 547.050 93.150 ;
        RECT 492.150 88.200 509.850 88.800 ;
        RECT 484.950 86.400 485.850 87.300 ;
        RECT 483.150 84.600 485.850 86.400 ;
        RECT 486.750 86.100 488.550 86.400 ;
        RECT 492.150 86.100 493.050 88.200 ;
        RECT 498.750 87.600 509.850 88.200 ;
        RECT 486.750 85.200 493.050 86.100 ;
        RECT 493.950 86.700 495.750 87.300 ;
        RECT 493.950 85.500 501.450 86.700 ;
        RECT 486.750 84.600 488.550 85.200 ;
        RECT 500.250 84.600 501.450 85.500 ;
        RECT 481.950 81.600 485.850 83.700 ;
        RECT 490.950 82.500 497.850 84.300 ;
        RECT 500.250 82.500 505.050 84.600 ;
        RECT 479.550 75.750 481.350 78.600 ;
        RECT 484.050 75.750 485.850 81.600 ;
        RECT 488.250 75.750 490.050 81.600 ;
        RECT 492.150 75.750 493.950 82.500 ;
        RECT 500.250 81.600 501.450 82.500 ;
        RECT 495.150 75.750 496.950 81.600 ;
        RECT 499.950 75.750 501.750 81.600 ;
        RECT 505.050 75.750 506.850 81.600 ;
        RECT 508.050 75.750 509.850 87.600 ;
        RECT 542.550 81.600 543.750 89.850 ;
        RECT 552.150 88.800 553.050 101.400 ;
        RECT 560.550 100.800 562.350 102.600 ;
        RECT 563.850 101.550 568.800 102.600 ;
        RECT 576.300 103.500 577.350 104.400 ;
        RECT 576.300 102.300 580.050 103.500 ;
        RECT 563.850 100.800 565.650 101.550 ;
        RECT 560.850 99.900 561.900 100.800 ;
        RECT 571.050 100.200 572.850 102.000 ;
        RECT 577.950 101.400 580.050 102.300 ;
        RECT 583.650 101.400 585.450 107.250 ;
        RECT 614.550 104.400 616.350 107.250 ;
        RECT 617.550 104.400 619.350 107.250 ;
        RECT 620.550 104.400 622.350 107.250 ;
        RECT 571.050 99.900 571.950 100.200 ;
        RECT 560.850 99.000 571.950 99.900 ;
        RECT 584.250 99.150 585.450 101.400 ;
        RECT 560.850 97.800 561.900 99.000 ;
        RECT 555.000 96.600 561.900 97.800 ;
        RECT 555.000 95.850 555.900 96.600 ;
        RECT 560.100 96.000 561.900 96.600 ;
        RECT 554.100 94.050 555.900 95.850 ;
        RECT 557.100 94.950 558.900 95.700 ;
        RECT 571.050 94.950 571.950 99.000 ;
        RECT 580.950 97.050 585.450 99.150 ;
        RECT 618.000 97.950 619.050 104.400 ;
        RECT 653.700 98.400 655.500 107.250 ;
        RECT 659.100 99.000 660.900 107.250 ;
        RECT 697.650 101.400 699.450 107.250 ;
        RECT 700.650 104.400 702.450 107.250 ;
        RECT 703.650 104.400 705.450 107.250 ;
        RECT 706.650 104.400 708.450 107.250 ;
        RECT 736.650 104.400 738.450 107.250 ;
        RECT 739.650 104.400 741.450 107.250 ;
        RECT 742.650 104.400 744.450 107.250 ;
        RECT 579.150 95.250 583.050 97.050 ;
        RECT 580.950 94.950 583.050 95.250 ;
        RECT 557.100 93.900 565.050 94.950 ;
        RECT 562.950 92.850 565.050 93.900 ;
        RECT 568.950 92.850 571.950 94.950 ;
        RECT 561.450 89.100 563.250 89.400 ;
        RECT 561.450 88.800 569.850 89.100 ;
        RECT 552.150 88.200 569.850 88.800 ;
        RECT 552.150 87.600 563.250 88.200 ;
        RECT 539.550 75.750 541.350 81.600 ;
        RECT 542.550 75.750 544.350 81.600 ;
        RECT 545.550 75.750 547.350 81.600 ;
        RECT 552.150 75.750 553.950 87.600 ;
        RECT 566.250 86.700 568.050 87.300 ;
        RECT 560.550 85.500 568.050 86.700 ;
        RECT 568.950 86.100 569.850 88.200 ;
        RECT 571.050 88.200 571.950 92.850 ;
        RECT 581.250 89.400 583.050 91.200 ;
        RECT 577.950 88.200 582.150 89.400 ;
        RECT 571.050 87.300 577.050 88.200 ;
        RECT 577.950 87.300 580.050 88.200 ;
        RECT 584.250 87.600 585.450 97.050 ;
        RECT 616.950 95.850 619.050 97.950 ;
        RECT 659.100 97.350 663.600 99.000 ;
        RECT 613.950 92.850 616.050 94.950 ;
        RECT 614.100 91.050 615.900 92.850 ;
        RECT 618.000 88.650 619.050 95.850 ;
        RECT 619.950 92.850 622.050 94.950 ;
        RECT 662.400 93.150 663.600 97.350 ;
        RECT 697.950 96.150 699.000 101.400 ;
        RECT 703.650 100.200 704.550 104.400 ;
        RECT 701.250 99.300 704.550 100.200 ;
        RECT 701.250 98.400 703.050 99.300 ;
        RECT 697.950 94.050 700.050 96.150 ;
        RECT 620.100 91.050 621.900 92.850 ;
        RECT 652.950 89.850 655.050 91.950 ;
        RECT 658.950 89.850 661.050 91.950 ;
        RECT 661.950 91.050 664.050 93.150 ;
        RECT 618.000 87.600 620.550 88.650 ;
        RECT 653.100 88.050 654.900 89.850 ;
        RECT 576.150 86.400 577.050 87.300 ;
        RECT 573.450 86.100 575.250 86.400 ;
        RECT 560.550 84.600 561.750 85.500 ;
        RECT 568.950 85.200 575.250 86.100 ;
        RECT 573.450 84.600 575.250 85.200 ;
        RECT 576.150 84.600 578.850 86.400 ;
        RECT 556.950 82.500 561.750 84.600 ;
        RECT 564.150 82.500 571.050 84.300 ;
        RECT 560.550 81.600 561.750 82.500 ;
        RECT 555.150 75.750 556.950 81.600 ;
        RECT 560.250 75.750 562.050 81.600 ;
        RECT 565.050 75.750 566.850 81.600 ;
        RECT 568.050 75.750 569.850 82.500 ;
        RECT 576.150 81.600 580.050 83.700 ;
        RECT 571.950 75.750 573.750 81.600 ;
        RECT 576.150 75.750 577.950 81.600 ;
        RECT 580.650 75.750 582.450 78.600 ;
        RECT 583.650 75.750 585.450 87.600 ;
        RECT 614.550 75.750 616.350 87.600 ;
        RECT 618.750 75.750 620.550 87.600 ;
        RECT 655.950 86.850 658.050 88.950 ;
        RECT 659.250 88.050 661.050 89.850 ;
        RECT 656.100 85.050 657.900 86.850 ;
        RECT 662.700 82.800 663.750 91.050 ;
        RECT 698.550 87.450 699.900 94.050 ;
        RECT 701.400 90.150 702.300 98.400 ;
        RECT 739.950 97.950 741.000 104.400 ;
        RECT 706.950 95.850 709.050 97.950 ;
        RECT 739.950 95.850 742.050 97.950 ;
        RECT 703.950 92.850 706.050 94.950 ;
        RECT 707.100 94.050 708.900 95.850 ;
        RECT 736.950 92.850 739.050 94.950 ;
        RECT 704.100 91.050 705.900 92.850 ;
        RECT 737.100 91.050 738.900 92.850 ;
        RECT 701.250 90.000 703.050 90.150 ;
        RECT 701.250 88.800 708.450 90.000 ;
        RECT 701.250 88.350 703.050 88.800 ;
        RECT 707.250 87.600 708.450 88.800 ;
        RECT 739.950 88.650 741.000 95.850 ;
        RECT 742.950 92.850 745.050 94.950 ;
        RECT 743.100 91.050 744.900 92.850 ;
        RECT 698.550 86.100 700.950 87.450 ;
        RECT 656.700 81.900 663.750 82.800 ;
        RECT 656.700 81.600 658.350 81.900 ;
        RECT 653.550 75.750 655.350 81.600 ;
        RECT 656.550 75.750 658.350 81.600 ;
        RECT 662.550 81.600 663.750 81.900 ;
        RECT 659.550 75.750 661.350 81.000 ;
        RECT 662.550 75.750 664.350 81.600 ;
        RECT 699.150 75.750 700.950 86.100 ;
        RECT 702.150 75.750 703.950 87.450 ;
        RECT 706.650 75.750 708.450 87.600 ;
        RECT 738.450 87.600 741.000 88.650 ;
        RECT 738.450 75.750 740.250 87.600 ;
        RECT 742.650 75.750 744.450 87.600 ;
        RECT 33.450 59.400 35.250 71.250 ;
        RECT 37.650 59.400 39.450 71.250 ;
        RECT 68.550 65.400 70.350 71.250 ;
        RECT 71.550 65.400 73.350 71.250 ;
        RECT 33.450 58.350 36.000 59.400 ;
        RECT 32.100 54.150 33.900 55.950 ;
        RECT 31.950 52.050 34.050 54.150 ;
        RECT 34.950 51.150 36.000 58.350 ;
        RECT 38.100 54.150 39.900 55.950 ;
        RECT 37.950 52.050 40.050 54.150 ;
        RECT 71.400 52.950 72.600 65.400 ;
        RECT 105.150 60.900 106.950 71.250 ;
        RECT 104.550 59.550 106.950 60.900 ;
        RECT 108.150 59.550 109.950 71.250 ;
        RECT 104.550 52.950 105.900 59.550 ;
        RECT 112.650 59.400 114.450 71.250 ;
        RECT 145.650 65.400 147.450 71.250 ;
        RECT 148.650 66.000 150.450 71.250 ;
        RECT 107.250 58.200 109.050 58.650 ;
        RECT 113.250 58.200 114.450 59.400 ;
        RECT 107.250 57.000 114.450 58.200 ;
        RECT 146.250 65.100 147.450 65.400 ;
        RECT 151.650 65.400 153.450 71.250 ;
        RECT 154.650 65.400 156.450 71.250 ;
        RECT 151.650 65.100 153.300 65.400 ;
        RECT 146.250 64.200 153.300 65.100 ;
        RECT 107.250 56.850 109.050 57.000 ;
        RECT 68.100 51.150 69.900 52.950 ;
        RECT 34.950 49.050 37.050 51.150 ;
        RECT 67.950 49.050 70.050 51.150 ;
        RECT 70.950 50.850 73.050 52.950 ;
        RECT 103.950 50.850 106.050 52.950 ;
        RECT 34.950 42.600 36.000 49.050 ;
        RECT 71.400 42.600 72.600 50.850 ;
        RECT 103.950 45.600 105.000 50.850 ;
        RECT 107.400 48.600 108.300 56.850 ;
        RECT 146.250 55.950 147.300 64.200 ;
        RECT 152.100 60.150 153.900 61.950 ;
        RECT 148.950 57.150 150.750 58.950 ;
        RECT 151.950 58.050 154.050 60.150 ;
        RECT 186.300 59.400 188.100 71.250 ;
        RECT 190.500 59.400 192.300 71.250 ;
        RECT 193.800 65.400 195.600 71.250 ;
        RECT 226.650 65.400 228.450 71.250 ;
        RECT 229.650 65.400 231.450 71.250 ;
        RECT 232.650 65.400 234.450 71.250 ;
        RECT 263.550 65.400 265.350 71.250 ;
        RECT 266.550 65.400 268.350 71.250 ;
        RECT 299.550 65.400 301.350 71.250 ;
        RECT 302.550 65.400 304.350 71.250 ;
        RECT 305.550 65.400 307.350 71.250 ;
        RECT 155.100 57.150 156.900 58.950 ;
        RECT 110.100 54.150 111.900 55.950 ;
        RECT 109.950 52.050 112.050 54.150 ;
        RECT 145.950 53.850 148.050 55.950 ;
        RECT 148.950 55.050 151.050 57.150 ;
        RECT 154.950 55.050 157.050 57.150 ;
        RECT 185.100 54.150 186.900 55.950 ;
        RECT 190.950 54.150 192.150 59.400 ;
        RECT 193.950 57.150 195.750 58.950 ;
        RECT 230.250 57.150 231.450 65.400 ;
        RECT 193.950 55.050 196.050 57.150 ;
        RECT 113.100 51.150 114.900 52.950 ;
        RECT 112.950 49.050 115.050 51.150 ;
        RECT 146.400 49.650 147.600 53.850 ;
        RECT 184.950 52.050 187.050 54.150 ;
        RECT 187.950 50.850 190.050 52.950 ;
        RECT 190.950 52.050 193.050 54.150 ;
        RECT 226.950 53.850 229.050 55.950 ;
        RECT 229.950 55.050 232.050 57.150 ;
        RECT 227.100 52.050 228.900 53.850 ;
        RECT 107.250 47.700 109.050 48.600 ;
        RECT 146.400 48.000 150.900 49.650 ;
        RECT 188.100 49.050 189.900 50.850 ;
        RECT 191.850 48.750 193.050 52.050 ;
        RECT 107.250 46.800 110.550 47.700 ;
        RECT 31.650 39.750 33.450 42.600 ;
        RECT 34.650 39.750 36.450 42.600 ;
        RECT 37.650 39.750 39.450 42.600 ;
        RECT 68.550 39.750 70.350 42.600 ;
        RECT 71.550 39.750 73.350 42.600 ;
        RECT 103.650 39.750 105.450 45.600 ;
        RECT 109.650 42.600 110.550 46.800 ;
        RECT 106.650 39.750 108.450 42.600 ;
        RECT 109.650 39.750 111.450 42.600 ;
        RECT 112.650 39.750 114.450 42.600 ;
        RECT 149.100 39.750 150.900 48.000 ;
        RECT 154.500 39.750 156.300 48.600 ;
        RECT 192.000 47.700 195.750 48.750 ;
        RECT 230.250 47.700 231.450 55.050 ;
        RECT 232.950 53.850 235.050 55.950 ;
        RECT 233.100 52.050 234.900 53.850 ;
        RECT 266.400 52.950 267.600 65.400 ;
        RECT 302.550 57.150 303.750 65.400 ;
        RECT 336.300 59.400 338.100 71.250 ;
        RECT 340.500 59.400 342.300 71.250 ;
        RECT 343.800 65.400 345.600 71.250 ;
        RECT 378.300 59.400 380.100 71.250 ;
        RECT 382.500 59.400 384.300 71.250 ;
        RECT 385.800 65.400 387.600 71.250 ;
        RECT 421.650 65.400 423.450 71.250 ;
        RECT 424.650 65.400 426.450 71.250 ;
        RECT 427.650 65.400 429.450 71.250 ;
        RECT 298.950 53.850 301.050 55.950 ;
        RECT 301.950 55.050 304.050 57.150 ;
        RECT 263.100 51.150 264.900 52.950 ;
        RECT 262.950 49.050 265.050 51.150 ;
        RECT 265.950 50.850 268.050 52.950 ;
        RECT 299.100 52.050 300.900 53.850 ;
        RECT 185.550 44.700 193.350 46.050 ;
        RECT 185.550 39.750 187.350 44.700 ;
        RECT 188.550 39.750 190.350 43.800 ;
        RECT 191.550 39.750 193.350 44.700 ;
        RECT 194.550 45.600 195.750 47.700 ;
        RECT 227.850 46.800 231.450 47.700 ;
        RECT 194.550 39.750 196.350 45.600 ;
        RECT 227.850 39.750 229.650 46.800 ;
        RECT 232.350 39.750 234.150 45.600 ;
        RECT 266.400 42.600 267.600 50.850 ;
        RECT 302.550 47.700 303.750 55.050 ;
        RECT 304.950 53.850 307.050 55.950 ;
        RECT 335.100 54.150 336.900 55.950 ;
        RECT 340.950 54.150 342.150 59.400 ;
        RECT 343.950 57.150 345.750 58.950 ;
        RECT 343.950 55.050 346.050 57.150 ;
        RECT 377.100 54.150 378.900 55.950 ;
        RECT 382.950 54.150 384.150 59.400 ;
        RECT 385.950 57.150 387.750 58.950 ;
        RECT 425.250 57.150 426.450 65.400 ;
        RECT 458.550 59.400 460.350 71.250 ;
        RECT 463.050 59.550 464.850 71.250 ;
        RECT 466.050 60.900 467.850 71.250 ;
        RECT 502.650 65.400 504.450 71.250 ;
        RECT 505.650 65.400 507.450 71.250 ;
        RECT 508.650 65.400 510.450 71.250 ;
        RECT 542.400 65.400 544.200 71.250 ;
        RECT 466.050 59.550 468.450 60.900 ;
        RECT 458.550 58.200 459.750 59.400 ;
        RECT 463.950 58.200 465.750 58.650 ;
        RECT 385.950 55.050 388.050 57.150 ;
        RECT 305.100 52.050 306.900 53.850 ;
        RECT 334.950 52.050 337.050 54.150 ;
        RECT 337.950 50.850 340.050 52.950 ;
        RECT 340.950 52.050 343.050 54.150 ;
        RECT 376.950 52.050 379.050 54.150 ;
        RECT 338.100 49.050 339.900 50.850 ;
        RECT 341.850 48.750 343.050 52.050 ;
        RECT 379.950 50.850 382.050 52.950 ;
        RECT 382.950 52.050 385.050 54.150 ;
        RECT 421.950 53.850 424.050 55.950 ;
        RECT 424.950 55.050 427.050 57.150 ;
        RECT 458.550 57.000 465.750 58.200 ;
        RECT 463.950 56.850 465.750 57.000 ;
        RECT 422.100 52.050 423.900 53.850 ;
        RECT 380.100 49.050 381.900 50.850 ;
        RECT 383.850 48.750 385.050 52.050 ;
        RECT 342.000 47.700 345.750 48.750 ;
        RECT 384.000 47.700 387.750 48.750 ;
        RECT 425.250 47.700 426.450 55.050 ;
        RECT 427.950 53.850 430.050 55.950 ;
        RECT 461.100 54.150 462.900 55.950 ;
        RECT 428.100 52.050 429.900 53.850 ;
        RECT 458.100 51.150 459.900 52.950 ;
        RECT 460.950 52.050 463.050 54.150 ;
        RECT 457.950 49.050 460.050 51.150 ;
        RECT 464.700 48.600 465.600 56.850 ;
        RECT 467.100 52.950 468.450 59.550 ;
        RECT 506.250 57.150 507.450 65.400 ;
        RECT 545.700 59.400 547.500 71.250 ;
        RECT 549.900 59.400 551.700 71.250 ;
        RECT 581.550 59.400 583.350 71.250 ;
        RECT 586.050 59.550 587.850 71.250 ;
        RECT 589.050 60.900 590.850 71.250 ;
        RECT 622.650 65.400 624.450 71.250 ;
        RECT 625.650 65.400 627.450 71.250 ;
        RECT 589.050 59.550 591.450 60.900 ;
        RECT 542.250 57.150 544.050 58.950 ;
        RECT 502.950 53.850 505.050 55.950 ;
        RECT 505.950 55.050 508.050 57.150 ;
        RECT 466.950 50.850 469.050 52.950 ;
        RECT 503.100 52.050 504.900 53.850 ;
        RECT 463.950 47.700 465.750 48.600 ;
        RECT 302.550 46.800 306.150 47.700 ;
        RECT 263.550 39.750 265.350 42.600 ;
        RECT 266.550 39.750 268.350 42.600 ;
        RECT 299.850 39.750 301.650 45.600 ;
        RECT 304.350 39.750 306.150 46.800 ;
        RECT 335.550 44.700 343.350 46.050 ;
        RECT 335.550 39.750 337.350 44.700 ;
        RECT 338.550 39.750 340.350 43.800 ;
        RECT 341.550 39.750 343.350 44.700 ;
        RECT 344.550 45.600 345.750 47.700 ;
        RECT 344.550 39.750 346.350 45.600 ;
        RECT 377.550 44.700 385.350 46.050 ;
        RECT 377.550 39.750 379.350 44.700 ;
        RECT 380.550 39.750 382.350 43.800 ;
        RECT 383.550 39.750 385.350 44.700 ;
        RECT 386.550 45.600 387.750 47.700 ;
        RECT 422.850 46.800 426.450 47.700 ;
        RECT 462.450 46.800 465.750 47.700 ;
        RECT 386.550 39.750 388.350 45.600 ;
        RECT 422.850 39.750 424.650 46.800 ;
        RECT 427.350 39.750 429.150 45.600 ;
        RECT 462.450 42.600 463.350 46.800 ;
        RECT 468.000 45.600 469.050 50.850 ;
        RECT 506.250 47.700 507.450 55.050 ;
        RECT 508.950 53.850 511.050 55.950 ;
        RECT 541.950 55.050 544.050 57.150 ;
        RECT 545.850 54.150 547.050 59.400 ;
        RECT 581.550 58.200 582.750 59.400 ;
        RECT 586.950 58.200 588.750 58.650 ;
        RECT 581.550 57.000 588.750 58.200 ;
        RECT 586.950 56.850 588.750 57.000 ;
        RECT 551.100 54.150 552.900 55.950 ;
        RECT 584.100 54.150 585.900 55.950 ;
        RECT 509.100 52.050 510.900 53.850 ;
        RECT 544.950 52.050 547.050 54.150 ;
        RECT 544.950 48.750 546.150 52.050 ;
        RECT 547.950 50.850 550.050 52.950 ;
        RECT 550.950 52.050 553.050 54.150 ;
        RECT 581.100 51.150 582.900 52.950 ;
        RECT 583.950 52.050 586.050 54.150 ;
        RECT 548.100 49.050 549.900 50.850 ;
        RECT 580.950 49.050 583.050 51.150 ;
        RECT 503.850 46.800 507.450 47.700 ;
        RECT 542.250 47.700 546.000 48.750 ;
        RECT 587.700 48.600 588.600 56.850 ;
        RECT 590.100 52.950 591.450 59.550 ;
        RECT 623.400 52.950 624.600 65.400 ;
        RECT 657.300 59.400 659.100 71.250 ;
        RECT 661.500 59.400 663.300 71.250 ;
        RECT 664.800 65.400 666.600 71.250 ;
        RECT 700.650 65.400 702.450 71.250 ;
        RECT 703.650 65.400 705.450 71.250 ;
        RECT 706.650 65.400 708.450 71.250 ;
        RECT 656.100 54.150 657.900 55.950 ;
        RECT 661.950 54.150 663.150 59.400 ;
        RECT 664.950 57.150 666.750 58.950 ;
        RECT 704.250 57.150 705.450 65.400 ;
        RECT 737.550 59.400 739.350 71.250 ;
        RECT 741.750 59.400 743.550 71.250 ;
        RECT 741.000 58.350 743.550 59.400 ;
        RECT 664.950 55.050 667.050 57.150 ;
        RECT 589.950 50.850 592.050 52.950 ;
        RECT 622.950 50.850 625.050 52.950 ;
        RECT 626.100 51.150 627.900 52.950 ;
        RECT 655.950 52.050 658.050 54.150 ;
        RECT 586.950 47.700 588.750 48.600 ;
        RECT 458.550 39.750 460.350 42.600 ;
        RECT 461.550 39.750 463.350 42.600 ;
        RECT 464.550 39.750 466.350 42.600 ;
        RECT 467.550 39.750 469.350 45.600 ;
        RECT 503.850 39.750 505.650 46.800 ;
        RECT 542.250 45.600 543.450 47.700 ;
        RECT 585.450 46.800 588.750 47.700 ;
        RECT 508.350 39.750 510.150 45.600 ;
        RECT 541.650 39.750 543.450 45.600 ;
        RECT 544.650 44.700 552.450 46.050 ;
        RECT 544.650 39.750 546.450 44.700 ;
        RECT 547.650 39.750 549.450 43.800 ;
        RECT 550.650 39.750 552.450 44.700 ;
        RECT 585.450 42.600 586.350 46.800 ;
        RECT 591.000 45.600 592.050 50.850 ;
        RECT 581.550 39.750 583.350 42.600 ;
        RECT 584.550 39.750 586.350 42.600 ;
        RECT 587.550 39.750 589.350 42.600 ;
        RECT 590.550 39.750 592.350 45.600 ;
        RECT 623.400 42.600 624.600 50.850 ;
        RECT 625.950 49.050 628.050 51.150 ;
        RECT 658.950 50.850 661.050 52.950 ;
        RECT 661.950 52.050 664.050 54.150 ;
        RECT 700.950 53.850 703.050 55.950 ;
        RECT 703.950 55.050 706.050 57.150 ;
        RECT 701.100 52.050 702.900 53.850 ;
        RECT 659.100 49.050 660.900 50.850 ;
        RECT 662.850 48.750 664.050 52.050 ;
        RECT 663.000 47.700 666.750 48.750 ;
        RECT 704.250 47.700 705.450 55.050 ;
        RECT 706.950 53.850 709.050 55.950 ;
        RECT 737.100 54.150 738.900 55.950 ;
        RECT 707.100 52.050 708.900 53.850 ;
        RECT 736.950 52.050 739.050 54.150 ;
        RECT 724.950 51.450 727.050 52.050 ;
        RECT 733.950 51.450 736.050 52.050 ;
        RECT 724.950 50.550 736.050 51.450 ;
        RECT 741.000 51.150 742.050 58.350 ;
        RECT 743.100 54.150 744.900 55.950 ;
        RECT 742.950 52.050 745.050 54.150 ;
        RECT 724.950 49.950 727.050 50.550 ;
        RECT 733.950 49.950 736.050 50.550 ;
        RECT 739.950 49.050 742.050 51.150 ;
        RECT 656.550 44.700 664.350 46.050 ;
        RECT 622.650 39.750 624.450 42.600 ;
        RECT 625.650 39.750 627.450 42.600 ;
        RECT 656.550 39.750 658.350 44.700 ;
        RECT 659.550 39.750 661.350 43.800 ;
        RECT 662.550 39.750 664.350 44.700 ;
        RECT 665.550 45.600 666.750 47.700 ;
        RECT 701.850 46.800 705.450 47.700 ;
        RECT 665.550 39.750 667.350 45.600 ;
        RECT 701.850 39.750 703.650 46.800 ;
        RECT 706.350 39.750 708.150 45.600 ;
        RECT 741.000 42.600 742.050 49.050 ;
        RECT 737.550 39.750 739.350 42.600 ;
        RECT 740.550 39.750 742.350 42.600 ;
        RECT 743.550 39.750 745.350 42.600 ;
        RECT 32.850 28.200 34.650 35.250 ;
        RECT 37.350 29.400 39.150 35.250 ;
        RECT 72.150 30.900 73.950 35.250 ;
        RECT 70.650 29.400 73.950 30.900 ;
        RECT 75.150 29.400 76.950 35.250 ;
        RECT 32.850 27.300 36.450 28.200 ;
        RECT 32.100 21.150 33.900 22.950 ;
        RECT 31.950 19.050 34.050 21.150 ;
        RECT 35.250 19.950 36.450 27.300 ;
        RECT 70.650 22.950 71.850 29.400 ;
        RECT 73.950 27.900 75.750 28.500 ;
        RECT 79.650 27.900 81.450 35.250 ;
        RECT 112.650 32.400 114.450 35.250 ;
        RECT 115.650 32.400 117.450 35.250 ;
        RECT 118.650 32.400 120.450 35.250 ;
        RECT 146.550 32.400 148.350 35.250 ;
        RECT 149.550 32.400 151.350 35.250 ;
        RECT 152.550 32.400 154.350 35.250 ;
        RECT 185.550 32.400 187.350 35.250 ;
        RECT 188.550 32.400 190.350 35.250 ;
        RECT 191.550 32.400 193.350 35.250 ;
        RECT 73.950 26.700 81.450 27.900 ;
        RECT 38.100 21.150 39.900 22.950 ;
        RECT 34.950 17.850 37.050 19.950 ;
        RECT 37.950 19.050 40.050 21.150 ;
        RECT 70.650 20.850 73.050 22.950 ;
        RECT 74.100 21.150 75.900 22.950 ;
        RECT 35.250 9.600 36.450 17.850 ;
        RECT 70.650 15.600 71.850 20.850 ;
        RECT 73.950 19.050 76.050 21.150 ;
        RECT 31.650 3.750 33.450 9.600 ;
        RECT 34.650 3.750 36.450 9.600 ;
        RECT 37.650 3.750 39.450 9.600 ;
        RECT 70.050 3.750 71.850 15.600 ;
        RECT 73.050 3.750 74.850 15.600 ;
        RECT 77.100 9.600 78.300 26.700 ;
        RECT 115.950 25.950 117.000 32.400 ;
        RECT 150.000 25.950 151.050 32.400 ;
        RECT 189.450 28.200 190.350 32.400 ;
        RECT 194.550 29.400 196.350 35.250 ;
        RECT 200.550 29.400 202.350 35.250 ;
        RECT 203.850 32.400 205.650 35.250 ;
        RECT 208.350 32.400 210.150 35.250 ;
        RECT 212.550 32.400 214.350 35.250 ;
        RECT 216.450 32.400 218.250 35.250 ;
        RECT 219.750 32.400 221.550 35.250 ;
        RECT 224.250 33.300 226.050 35.250 ;
        RECT 224.250 32.400 228.000 33.300 ;
        RECT 229.050 32.400 230.850 35.250 ;
        RECT 208.650 31.500 209.700 32.400 ;
        RECT 205.950 30.300 209.700 31.500 ;
        RECT 217.200 30.600 218.250 32.400 ;
        RECT 226.950 31.500 228.000 32.400 ;
        RECT 205.950 29.400 208.050 30.300 ;
        RECT 189.450 27.300 192.750 28.200 ;
        RECT 190.950 26.400 192.750 27.300 ;
        RECT 115.950 23.850 118.050 25.950 ;
        RECT 148.950 23.850 151.050 25.950 ;
        RECT 184.950 23.850 187.050 25.950 ;
        RECT 79.950 20.850 82.050 22.950 ;
        RECT 112.950 20.850 115.050 22.950 ;
        RECT 80.100 19.050 81.900 20.850 ;
        RECT 113.100 19.050 114.900 20.850 ;
        RECT 115.950 16.650 117.000 23.850 ;
        RECT 118.950 20.850 121.050 22.950 ;
        RECT 145.950 20.850 148.050 22.950 ;
        RECT 119.100 19.050 120.900 20.850 ;
        RECT 146.100 19.050 147.900 20.850 ;
        RECT 114.450 15.600 117.000 16.650 ;
        RECT 150.000 16.650 151.050 23.850 ;
        RECT 151.950 20.850 154.050 22.950 ;
        RECT 185.100 22.050 186.900 23.850 ;
        RECT 187.950 20.850 190.050 22.950 ;
        RECT 152.100 19.050 153.900 20.850 ;
        RECT 188.100 19.050 189.900 20.850 ;
        RECT 191.700 18.150 192.600 26.400 ;
        RECT 195.000 24.150 196.050 29.400 ;
        RECT 193.950 22.050 196.050 24.150 ;
        RECT 200.550 27.150 201.750 29.400 ;
        RECT 213.150 28.200 214.950 30.000 ;
        RECT 217.200 29.550 222.150 30.600 ;
        RECT 220.350 28.800 222.150 29.550 ;
        RECT 223.650 28.800 225.450 30.600 ;
        RECT 226.950 29.400 229.050 31.500 ;
        RECT 232.050 29.400 233.850 35.250 ;
        RECT 214.050 27.900 214.950 28.200 ;
        RECT 224.100 27.900 225.150 28.800 ;
        RECT 200.550 25.050 205.050 27.150 ;
        RECT 214.050 27.000 225.150 27.900 ;
        RECT 190.950 18.000 192.750 18.150 ;
        RECT 185.550 16.800 192.750 18.000 ;
        RECT 150.000 15.600 152.550 16.650 ;
        RECT 76.650 3.750 78.450 9.600 ;
        RECT 79.650 3.750 81.450 9.600 ;
        RECT 114.450 3.750 116.250 15.600 ;
        RECT 118.650 3.750 120.450 15.600 ;
        RECT 146.550 3.750 148.350 15.600 ;
        RECT 150.750 3.750 152.550 15.600 ;
        RECT 185.550 15.600 186.750 16.800 ;
        RECT 190.950 16.350 192.750 16.800 ;
        RECT 185.550 3.750 187.350 15.600 ;
        RECT 194.100 15.450 195.450 22.050 ;
        RECT 190.050 3.750 191.850 15.450 ;
        RECT 193.050 14.100 195.450 15.450 ;
        RECT 200.550 15.600 201.750 25.050 ;
        RECT 202.950 23.250 206.850 25.050 ;
        RECT 202.950 22.950 205.050 23.250 ;
        RECT 214.050 22.950 214.950 27.000 ;
        RECT 224.100 25.800 225.150 27.000 ;
        RECT 224.100 24.600 231.000 25.800 ;
        RECT 224.100 24.000 225.900 24.600 ;
        RECT 230.100 23.850 231.000 24.600 ;
        RECT 227.100 22.950 228.900 23.700 ;
        RECT 214.050 20.850 217.050 22.950 ;
        RECT 220.950 21.900 228.900 22.950 ;
        RECT 230.100 22.050 231.900 23.850 ;
        RECT 220.950 20.850 223.050 21.900 ;
        RECT 202.950 17.400 204.750 19.200 ;
        RECT 203.850 16.200 208.050 17.400 ;
        RECT 214.050 16.200 214.950 20.850 ;
        RECT 222.750 17.100 224.550 17.400 ;
        RECT 193.050 3.750 194.850 14.100 ;
        RECT 200.550 3.750 202.350 15.600 ;
        RECT 205.950 15.300 208.050 16.200 ;
        RECT 208.950 15.300 214.950 16.200 ;
        RECT 216.150 16.800 224.550 17.100 ;
        RECT 232.950 16.800 233.850 29.400 ;
        RECT 216.150 16.200 233.850 16.800 ;
        RECT 208.950 14.400 209.850 15.300 ;
        RECT 207.150 12.600 209.850 14.400 ;
        RECT 210.750 14.100 212.550 14.400 ;
        RECT 216.150 14.100 217.050 16.200 ;
        RECT 222.750 15.600 233.850 16.200 ;
        RECT 210.750 13.200 217.050 14.100 ;
        RECT 217.950 14.700 219.750 15.300 ;
        RECT 217.950 13.500 225.450 14.700 ;
        RECT 210.750 12.600 212.550 13.200 ;
        RECT 224.250 12.600 225.450 13.500 ;
        RECT 205.950 9.600 209.850 11.700 ;
        RECT 214.950 10.500 221.850 12.300 ;
        RECT 224.250 10.500 229.050 12.600 ;
        RECT 203.550 3.750 205.350 6.600 ;
        RECT 208.050 3.750 209.850 9.600 ;
        RECT 212.250 3.750 214.050 9.600 ;
        RECT 216.150 3.750 217.950 10.500 ;
        RECT 224.250 9.600 225.450 10.500 ;
        RECT 219.150 3.750 220.950 9.600 ;
        RECT 223.950 3.750 225.750 9.600 ;
        RECT 229.050 3.750 230.850 9.600 ;
        RECT 232.050 3.750 233.850 15.600 ;
        RECT 237.150 29.400 238.950 35.250 ;
        RECT 240.150 32.400 241.950 35.250 ;
        RECT 244.950 33.300 246.750 35.250 ;
        RECT 243.000 32.400 246.750 33.300 ;
        RECT 249.450 32.400 251.250 35.250 ;
        RECT 252.750 32.400 254.550 35.250 ;
        RECT 256.650 32.400 258.450 35.250 ;
        RECT 260.850 32.400 262.650 35.250 ;
        RECT 265.350 32.400 267.150 35.250 ;
        RECT 243.000 31.500 244.050 32.400 ;
        RECT 241.950 29.400 244.050 31.500 ;
        RECT 252.750 30.600 253.800 32.400 ;
        RECT 237.150 16.800 238.050 29.400 ;
        RECT 245.550 28.800 247.350 30.600 ;
        RECT 248.850 29.550 253.800 30.600 ;
        RECT 261.300 31.500 262.350 32.400 ;
        RECT 261.300 30.300 265.050 31.500 ;
        RECT 248.850 28.800 250.650 29.550 ;
        RECT 245.850 27.900 246.900 28.800 ;
        RECT 256.050 28.200 257.850 30.000 ;
        RECT 262.950 29.400 265.050 30.300 ;
        RECT 268.650 29.400 270.450 35.250 ;
        RECT 302.700 32.400 304.500 35.250 ;
        RECT 306.000 31.050 307.800 35.250 ;
        RECT 256.050 27.900 256.950 28.200 ;
        RECT 245.850 27.000 256.950 27.900 ;
        RECT 269.250 27.150 270.450 29.400 ;
        RECT 245.850 25.800 246.900 27.000 ;
        RECT 240.000 24.600 246.900 25.800 ;
        RECT 240.000 23.850 240.900 24.600 ;
        RECT 245.100 24.000 246.900 24.600 ;
        RECT 239.100 22.050 240.900 23.850 ;
        RECT 242.100 22.950 243.900 23.700 ;
        RECT 256.050 22.950 256.950 27.000 ;
        RECT 265.950 25.050 270.450 27.150 ;
        RECT 264.150 23.250 268.050 25.050 ;
        RECT 265.950 22.950 268.050 23.250 ;
        RECT 242.100 21.900 250.050 22.950 ;
        RECT 247.950 20.850 250.050 21.900 ;
        RECT 253.950 20.850 256.950 22.950 ;
        RECT 246.450 17.100 248.250 17.400 ;
        RECT 246.450 16.800 254.850 17.100 ;
        RECT 237.150 16.200 254.850 16.800 ;
        RECT 237.150 15.600 248.250 16.200 ;
        RECT 237.150 3.750 238.950 15.600 ;
        RECT 251.250 14.700 253.050 15.300 ;
        RECT 245.550 13.500 253.050 14.700 ;
        RECT 253.950 14.100 254.850 16.200 ;
        RECT 256.050 16.200 256.950 20.850 ;
        RECT 266.250 17.400 268.050 19.200 ;
        RECT 262.950 16.200 267.150 17.400 ;
        RECT 256.050 15.300 262.050 16.200 ;
        RECT 262.950 15.300 265.050 16.200 ;
        RECT 269.250 15.600 270.450 25.050 ;
        RECT 302.100 29.400 307.800 31.050 ;
        RECT 310.200 29.400 312.000 35.250 ;
        RECT 341.550 32.400 343.350 35.250 ;
        RECT 344.550 32.400 346.350 35.250 ;
        RECT 347.550 32.400 349.350 35.250 ;
        RECT 302.100 22.950 303.300 29.400 ;
        RECT 345.000 25.950 346.050 32.400 ;
        RECT 380.550 30.300 382.350 35.250 ;
        RECT 383.550 31.200 385.350 35.250 ;
        RECT 386.550 30.300 388.350 35.250 ;
        RECT 380.550 28.950 388.350 30.300 ;
        RECT 389.550 29.400 391.350 35.250 ;
        RECT 424.650 32.400 426.450 35.250 ;
        RECT 427.650 32.400 429.450 35.250 ;
        RECT 430.650 32.400 432.450 35.250 ;
        RECT 389.550 27.300 390.750 29.400 ;
        RECT 387.000 26.250 390.750 27.300 ;
        RECT 305.100 24.150 306.900 25.950 ;
        RECT 301.950 20.850 304.050 22.950 ;
        RECT 304.950 22.050 307.050 24.150 ;
        RECT 307.950 23.850 310.050 25.950 ;
        RECT 311.100 24.150 312.900 25.950 ;
        RECT 308.100 22.050 309.900 23.850 ;
        RECT 310.950 22.050 313.050 24.150 ;
        RECT 343.950 23.850 346.050 25.950 ;
        RECT 383.100 24.150 384.900 25.950 ;
        RECT 340.950 20.850 343.050 22.950 ;
        RECT 302.100 15.600 303.300 20.850 ;
        RECT 341.100 19.050 342.900 20.850 ;
        RECT 345.000 16.650 346.050 23.850 ;
        RECT 346.950 20.850 349.050 22.950 ;
        RECT 379.950 20.850 382.050 22.950 ;
        RECT 382.950 22.050 385.050 24.150 ;
        RECT 386.850 22.950 388.050 26.250 ;
        RECT 427.950 25.950 429.000 32.400 ;
        RECT 464.850 28.200 466.650 35.250 ;
        RECT 469.350 29.400 471.150 35.250 ;
        RECT 502.650 32.400 504.450 35.250 ;
        RECT 505.650 32.400 507.450 35.250 ;
        RECT 508.650 32.400 510.450 35.250 ;
        RECT 464.850 27.300 468.450 28.200 ;
        RECT 427.950 23.850 430.050 25.950 ;
        RECT 385.950 20.850 388.050 22.950 ;
        RECT 424.950 20.850 427.050 22.950 ;
        RECT 347.100 19.050 348.900 20.850 ;
        RECT 380.100 19.050 381.900 20.850 ;
        RECT 345.000 15.600 347.550 16.650 ;
        RECT 385.950 15.600 387.150 20.850 ;
        RECT 388.950 17.850 391.050 19.950 ;
        RECT 425.100 19.050 426.900 20.850 ;
        RECT 388.950 16.050 390.750 17.850 ;
        RECT 427.950 16.650 429.000 23.850 ;
        RECT 430.950 20.850 433.050 22.950 ;
        RECT 464.100 21.150 465.900 22.950 ;
        RECT 431.100 19.050 432.900 20.850 ;
        RECT 463.950 19.050 466.050 21.150 ;
        RECT 467.250 19.950 468.450 27.300 ;
        RECT 505.950 25.950 507.000 32.400 ;
        RECT 539.550 30.300 541.350 35.250 ;
        RECT 542.550 31.200 544.350 35.250 ;
        RECT 545.550 30.300 547.350 35.250 ;
        RECT 539.550 28.950 547.350 30.300 ;
        RECT 548.550 29.400 550.350 35.250 ;
        RECT 548.550 27.300 549.750 29.400 ;
        RECT 584.850 28.200 586.650 35.250 ;
        RECT 589.350 29.400 591.150 35.250 ;
        RECT 620.850 29.400 622.650 35.250 ;
        RECT 625.350 28.200 627.150 35.250 ;
        RECT 659.550 32.400 661.350 35.250 ;
        RECT 662.550 32.400 664.350 35.250 ;
        RECT 584.850 27.300 588.450 28.200 ;
        RECT 546.000 26.250 549.750 27.300 ;
        RECT 505.950 23.850 508.050 25.950 ;
        RECT 542.100 24.150 543.900 25.950 ;
        RECT 470.100 21.150 471.900 22.950 ;
        RECT 466.950 17.850 469.050 19.950 ;
        RECT 469.950 19.050 472.050 21.150 ;
        RECT 502.950 20.850 505.050 22.950 ;
        RECT 503.100 19.050 504.900 20.850 ;
        RECT 426.450 15.600 429.000 16.650 ;
        RECT 261.150 14.400 262.050 15.300 ;
        RECT 258.450 14.100 260.250 14.400 ;
        RECT 245.550 12.600 246.750 13.500 ;
        RECT 253.950 13.200 260.250 14.100 ;
        RECT 258.450 12.600 260.250 13.200 ;
        RECT 261.150 12.600 263.850 14.400 ;
        RECT 241.950 10.500 246.750 12.600 ;
        RECT 249.150 10.500 256.050 12.300 ;
        RECT 245.550 9.600 246.750 10.500 ;
        RECT 240.150 3.750 241.950 9.600 ;
        RECT 245.250 3.750 247.050 9.600 ;
        RECT 250.050 3.750 251.850 9.600 ;
        RECT 253.050 3.750 254.850 10.500 ;
        RECT 261.150 9.600 265.050 11.700 ;
        RECT 256.950 3.750 258.750 9.600 ;
        RECT 261.150 3.750 262.950 9.600 ;
        RECT 265.650 3.750 267.450 6.600 ;
        RECT 268.650 3.750 270.450 15.600 ;
        RECT 301.650 3.750 303.450 15.600 ;
        RECT 304.650 14.700 312.450 15.600 ;
        RECT 304.650 3.750 306.450 14.700 ;
        RECT 307.650 3.750 309.450 13.800 ;
        RECT 310.650 3.750 312.450 14.700 ;
        RECT 341.550 3.750 343.350 15.600 ;
        RECT 345.750 3.750 347.550 15.600 ;
        RECT 381.300 3.750 383.100 15.600 ;
        RECT 385.500 3.750 387.300 15.600 ;
        RECT 388.800 3.750 390.600 9.600 ;
        RECT 426.450 3.750 428.250 15.600 ;
        RECT 430.650 3.750 432.450 15.600 ;
        RECT 467.250 9.600 468.450 17.850 ;
        RECT 505.950 16.650 507.000 23.850 ;
        RECT 508.950 20.850 511.050 22.950 ;
        RECT 538.950 20.850 541.050 22.950 ;
        RECT 541.950 22.050 544.050 24.150 ;
        RECT 545.850 22.950 547.050 26.250 ;
        RECT 544.950 20.850 547.050 22.950 ;
        RECT 584.100 21.150 585.900 22.950 ;
        RECT 509.100 19.050 510.900 20.850 ;
        RECT 539.100 19.050 540.900 20.850 ;
        RECT 504.450 15.600 507.000 16.650 ;
        RECT 544.950 15.600 546.150 20.850 ;
        RECT 547.950 17.850 550.050 19.950 ;
        RECT 583.950 19.050 586.050 21.150 ;
        RECT 587.250 19.950 588.450 27.300 ;
        RECT 623.550 27.300 627.150 28.200 ;
        RECT 590.100 21.150 591.900 22.950 ;
        RECT 620.100 21.150 621.900 22.950 ;
        RECT 586.950 17.850 589.050 19.950 ;
        RECT 589.950 19.050 592.050 21.150 ;
        RECT 619.950 19.050 622.050 21.150 ;
        RECT 623.550 19.950 624.750 27.300 ;
        RECT 658.950 23.850 661.050 25.950 ;
        RECT 662.400 24.150 663.600 32.400 ;
        RECT 695.850 28.200 697.650 35.250 ;
        RECT 700.350 29.400 702.150 35.250 ;
        RECT 731.550 32.400 733.350 35.250 ;
        RECT 734.550 32.400 736.350 35.250 ;
        RECT 695.850 27.300 699.450 28.200 ;
        RECT 626.100 21.150 627.900 22.950 ;
        RECT 659.100 22.050 660.900 23.850 ;
        RECT 661.950 22.050 664.050 24.150 ;
        RECT 622.950 17.850 625.050 19.950 ;
        RECT 625.950 19.050 628.050 21.150 ;
        RECT 547.950 16.050 549.750 17.850 ;
        RECT 463.650 3.750 465.450 9.600 ;
        RECT 466.650 3.750 468.450 9.600 ;
        RECT 469.650 3.750 471.450 9.600 ;
        RECT 504.450 3.750 506.250 15.600 ;
        RECT 508.650 3.750 510.450 15.600 ;
        RECT 540.300 3.750 542.100 15.600 ;
        RECT 544.500 3.750 546.300 15.600 ;
        RECT 587.250 9.600 588.450 17.850 ;
        RECT 623.550 9.600 624.750 17.850 ;
        RECT 662.400 9.600 663.600 22.050 ;
        RECT 695.100 21.150 696.900 22.950 ;
        RECT 694.950 19.050 697.050 21.150 ;
        RECT 698.250 19.950 699.450 27.300 ;
        RECT 730.950 23.850 733.050 25.950 ;
        RECT 734.400 24.150 735.600 32.400 ;
        RECT 701.100 21.150 702.900 22.950 ;
        RECT 731.100 22.050 732.900 23.850 ;
        RECT 733.950 22.050 736.050 24.150 ;
        RECT 697.950 17.850 700.050 19.950 ;
        RECT 700.950 19.050 703.050 21.150 ;
        RECT 698.250 9.600 699.450 17.850 ;
        RECT 734.400 9.600 735.600 22.050 ;
        RECT 547.800 3.750 549.600 9.600 ;
        RECT 583.650 3.750 585.450 9.600 ;
        RECT 586.650 3.750 588.450 9.600 ;
        RECT 589.650 3.750 591.450 9.600 ;
        RECT 620.550 3.750 622.350 9.600 ;
        RECT 623.550 3.750 625.350 9.600 ;
        RECT 626.550 3.750 628.350 9.600 ;
        RECT 659.550 3.750 661.350 9.600 ;
        RECT 662.550 3.750 664.350 9.600 ;
        RECT 694.650 3.750 696.450 9.600 ;
        RECT 697.650 3.750 699.450 9.600 ;
        RECT 700.650 3.750 702.450 9.600 ;
        RECT 731.550 3.750 733.350 9.600 ;
        RECT 734.550 3.750 736.350 9.600 ;
      LAYER metal2 ;
        RECT 70.950 704.250 73.050 705.150 ;
        RECT 112.950 703.950 115.050 706.050 ;
        RECT 145.950 705.450 148.050 706.050 ;
        RECT 143.400 704.400 148.050 705.450 ;
        RECT 113.400 703.050 114.450 703.950 ;
        RECT 31.950 701.250 34.050 702.150 ;
        RECT 37.950 701.250 40.050 702.150 ;
        RECT 64.950 700.950 67.050 703.050 ;
        RECT 70.950 700.950 73.050 703.050 ;
        RECT 74.250 701.250 75.750 702.150 ;
        RECT 76.950 700.950 79.050 703.050 ;
        RECT 80.250 701.250 82.050 702.150 ;
        RECT 112.950 700.950 115.050 703.050 ;
        RECT 35.250 698.250 36.750 699.150 ;
        RECT 37.950 697.950 40.050 700.050 ;
        RECT 34.950 694.950 37.050 697.050 ;
        RECT 38.400 694.050 39.450 697.950 ;
        RECT 37.950 691.950 40.050 694.050 ;
        RECT 28.950 668.250 30.750 669.150 ;
        RECT 31.950 667.950 34.050 670.050 ;
        RECT 35.250 668.250 37.050 669.150 ;
        RECT 32.250 665.850 33.750 666.750 ;
        RECT 34.950 666.450 37.050 667.050 ;
        RECT 38.400 666.450 39.450 691.950 ;
        RECT 65.400 676.050 66.450 700.950 ;
        RECT 71.400 682.050 72.450 700.950 ;
        RECT 143.400 700.050 144.450 704.400 ;
        RECT 145.950 703.950 148.050 704.400 ;
        RECT 149.250 704.250 150.750 705.150 ;
        RECT 151.950 703.950 154.050 706.050 ;
        RECT 502.950 705.450 505.050 706.050 ;
        RECT 193.950 704.250 196.050 705.150 ;
        RECT 274.950 704.250 277.050 705.150 ;
        RECT 500.400 704.400 505.050 705.450 ;
        RECT 145.950 701.850 147.750 702.750 ;
        RECT 148.950 700.950 151.050 703.050 ;
        RECT 152.250 701.850 154.050 702.750 ;
        RECT 184.950 701.250 186.750 702.150 ;
        RECT 187.950 700.950 190.050 703.050 ;
        RECT 193.950 702.450 196.050 703.050 ;
        RECT 196.950 702.450 199.050 703.050 ;
        RECT 191.250 701.250 192.750 702.150 ;
        RECT 193.950 701.400 199.050 702.450 ;
        RECT 193.950 700.950 196.050 701.400 ;
        RECT 196.950 700.950 199.050 701.400 ;
        RECT 199.950 700.950 202.050 703.050 ;
        RECT 202.950 700.950 205.050 703.050 ;
        RECT 223.950 702.450 226.050 703.050 ;
        RECT 221.400 701.400 226.050 702.450 ;
        RECT 149.400 700.050 150.450 700.950 ;
        RECT 73.950 697.950 76.050 700.050 ;
        RECT 77.250 698.850 78.750 699.750 ;
        RECT 79.950 697.950 82.050 700.050 ;
        RECT 109.950 698.250 112.050 699.150 ;
        RECT 112.950 698.850 115.050 699.750 ;
        RECT 142.950 697.950 145.050 700.050 ;
        RECT 148.950 697.950 151.050 700.050 ;
        RECT 184.950 697.950 187.050 700.050 ;
        RECT 188.250 698.850 189.750 699.750 ;
        RECT 190.950 697.950 193.050 700.050 ;
        RECT 193.950 697.950 196.050 700.050 ;
        RECT 200.400 699.450 201.450 700.950 ;
        RECT 197.400 698.400 201.450 699.450 ;
        RECT 80.400 697.050 81.450 697.950 ;
        RECT 73.950 694.950 76.050 697.050 ;
        RECT 79.950 694.950 82.050 697.050 ;
        RECT 109.950 694.950 112.050 697.050 ;
        RECT 70.950 679.950 73.050 682.050 ;
        RECT 64.950 673.950 67.050 676.050 ;
        RECT 40.950 667.950 43.050 670.050 ;
        RECT 34.950 665.400 39.450 666.450 ;
        RECT 34.950 664.950 37.050 665.400 ;
        RECT 31.950 649.950 34.050 652.050 ;
        RECT 32.400 631.050 33.450 649.950 ;
        RECT 31.950 628.950 34.050 631.050 ;
        RECT 31.950 626.850 34.050 627.750 ;
        RECT 34.950 626.250 37.050 627.150 ;
        RECT 41.400 625.050 42.450 667.950 ;
        RECT 65.400 652.050 66.450 673.950 ;
        RECT 74.400 673.050 75.450 694.950 ;
        RECT 103.950 679.950 106.050 682.050 ;
        RECT 104.400 676.050 105.450 679.950 ;
        RECT 110.400 676.050 111.450 694.950 ;
        RECT 185.400 694.050 186.450 697.950 ;
        RECT 184.950 691.950 187.050 694.050 ;
        RECT 191.400 693.450 192.450 697.950 ;
        RECT 194.400 697.050 195.450 697.950 ;
        RECT 193.950 694.950 196.050 697.050 ;
        RECT 197.400 693.450 198.450 698.400 ;
        RECT 191.400 692.400 198.450 693.450 ;
        RECT 203.400 691.050 204.450 700.950 ;
        RECT 221.400 700.050 222.450 701.400 ;
        RECT 223.950 700.950 226.050 701.400 ;
        RECT 229.950 700.950 232.050 703.050 ;
        RECT 233.250 701.250 235.050 702.150 ;
        RECT 262.950 700.950 265.050 703.050 ;
        RECT 265.950 701.250 267.750 702.150 ;
        RECT 268.950 700.950 271.050 703.050 ;
        RECT 272.250 701.250 273.750 702.150 ;
        RECT 274.950 700.950 277.050 703.050 ;
        RECT 304.950 701.250 307.050 702.150 ;
        RECT 310.950 701.250 313.050 702.150 ;
        RECT 343.950 701.250 346.050 702.150 ;
        RECT 349.950 701.850 352.050 702.750 ;
        RECT 466.950 702.450 469.050 703.050 ;
        RECT 352.950 701.250 355.050 702.150 ;
        RECT 385.950 701.250 388.050 702.150 ;
        RECT 391.950 701.250 394.050 702.150 ;
        RECT 424.950 701.250 427.050 702.150 ;
        RECT 430.950 701.250 433.050 702.150 ;
        RECT 464.400 701.400 469.050 702.450 ;
        RECT 214.950 697.950 217.050 700.050 ;
        RECT 220.950 697.950 223.050 700.050 ;
        RECT 223.950 698.850 226.050 699.750 ;
        RECT 226.950 698.250 229.050 699.150 ;
        RECT 229.950 698.850 231.750 699.750 ;
        RECT 232.950 697.950 235.050 700.050 ;
        RECT 215.400 697.050 216.450 697.950 ;
        RECT 214.950 694.950 217.050 697.050 ;
        RECT 226.950 694.950 229.050 697.050 ;
        RECT 202.950 688.950 205.050 691.050 ;
        RECT 121.950 677.400 124.050 679.500 ;
        RECT 142.950 677.400 145.050 679.500 ;
        RECT 76.950 673.950 79.050 676.050 ;
        RECT 103.950 673.950 106.050 676.050 ;
        RECT 109.950 673.950 112.050 676.050 ;
        RECT 112.950 673.950 115.050 676.050 ;
        RECT 118.950 674.250 121.050 675.150 ;
        RECT 73.950 672.450 76.050 673.050 ;
        RECT 67.950 671.250 70.050 672.150 ;
        RECT 71.400 671.400 76.050 672.450 ;
        RECT 77.250 671.850 79.050 672.750 ;
        RECT 67.950 667.950 70.050 670.050 ;
        RECT 64.950 649.950 67.050 652.050 ;
        RECT 71.400 633.450 72.450 671.400 ;
        RECT 73.950 670.950 76.050 671.400 ;
        RECT 73.950 668.850 76.050 669.750 ;
        RECT 94.950 661.950 97.050 664.050 ;
        RECT 67.950 632.250 70.050 633.150 ;
        RECT 71.400 632.400 75.450 633.450 ;
        RECT 74.400 631.050 75.450 632.400 ;
        RECT 67.950 628.950 70.050 631.050 ;
        RECT 71.250 629.250 72.750 630.150 ;
        RECT 73.950 628.950 76.050 631.050 ;
        RECT 77.250 629.250 79.050 630.150 ;
        RECT 68.400 625.050 69.450 628.950 ;
        RECT 70.950 625.950 73.050 628.050 ;
        RECT 74.250 626.850 75.750 627.750 ;
        RECT 76.950 625.950 79.050 628.050 ;
        RECT 34.950 622.950 37.050 625.050 ;
        RECT 40.950 622.950 43.050 625.050 ;
        RECT 67.950 622.950 70.050 625.050 ;
        RECT 46.950 605.400 49.050 607.500 ;
        RECT 67.950 605.400 70.050 607.500 ;
        RECT 34.950 601.950 37.050 604.050 ;
        RECT 43.950 602.250 46.050 603.150 ;
        RECT 35.250 599.850 36.750 600.750 ;
        RECT 37.950 598.950 40.050 601.050 ;
        RECT 43.950 598.950 46.050 601.050 ;
        RECT 31.950 596.850 34.050 597.750 ;
        RECT 37.950 596.850 40.050 597.750 ;
        RECT 44.400 565.050 45.450 598.950 ;
        RECT 47.550 593.400 48.750 605.400 ;
        RECT 49.950 601.950 52.050 604.050 ;
        RECT 55.950 601.950 58.050 604.050 ;
        RECT 46.950 591.300 49.050 593.400 ;
        RECT 47.550 587.700 48.750 591.300 ;
        RECT 46.950 585.600 49.050 587.700 ;
        RECT 43.950 562.950 46.050 565.050 ;
        RECT 31.950 557.250 34.050 558.150 ;
        RECT 34.950 557.850 37.050 558.750 ;
        RECT 40.950 557.250 43.050 558.150 ;
        RECT 31.950 553.950 34.050 556.050 ;
        RECT 40.950 555.450 43.050 556.050 ;
        RECT 44.400 555.450 45.450 562.950 ;
        RECT 50.400 556.050 51.450 601.950 ;
        RECT 56.400 601.050 57.450 601.950 ;
        RECT 55.950 598.950 58.050 601.050 ;
        RECT 61.950 598.950 64.050 601.050 ;
        RECT 55.950 596.850 58.050 597.750 ;
        RECT 61.950 596.850 64.050 597.750 ;
        RECT 68.400 588.600 69.600 605.400 ;
        RECT 67.950 586.500 70.050 588.600 ;
        RECT 71.400 562.050 72.450 625.950 ;
        RECT 82.950 605.400 85.050 607.500 ;
        RECT 79.950 598.950 82.050 601.050 ;
        RECT 64.950 559.950 67.050 562.050 ;
        RECT 70.950 559.950 73.050 562.050 ;
        RECT 40.950 554.400 45.450 555.450 ;
        RECT 40.950 553.950 43.050 554.400 ;
        RECT 49.950 553.950 52.050 556.050 ;
        RECT 32.400 553.050 33.450 553.950 ;
        RECT 31.950 550.950 34.050 553.050 ;
        RECT 37.950 529.950 40.050 532.050 ;
        RECT 38.400 529.050 39.450 529.950 ;
        RECT 65.400 529.050 66.450 559.950 ;
        RECT 70.950 557.250 73.050 558.150 ;
        RECT 76.950 557.250 79.050 558.150 ;
        RECT 80.400 556.050 81.450 598.950 ;
        RECT 83.400 588.600 84.600 605.400 ;
        RECT 95.400 604.050 96.450 661.950 ;
        RECT 104.400 628.050 105.450 673.950 ;
        RECT 113.400 673.050 114.450 673.950 ;
        RECT 106.950 670.950 109.050 673.050 ;
        RECT 110.250 671.850 111.750 672.750 ;
        RECT 112.950 670.950 115.050 673.050 ;
        RECT 118.950 670.950 121.050 673.050 ;
        RECT 106.950 668.850 109.050 669.750 ;
        RECT 112.950 668.850 115.050 669.750 ;
        RECT 115.950 633.450 118.050 634.050 ;
        RECT 119.400 633.450 120.450 670.950 ;
        RECT 122.550 665.400 123.750 677.400 ;
        RECT 130.950 672.450 133.050 673.050 ;
        RECT 130.950 671.400 135.450 672.450 ;
        RECT 130.950 670.950 133.050 671.400 ;
        RECT 130.950 668.850 133.050 669.750 ;
        RECT 121.950 663.300 124.050 665.400 ;
        RECT 134.400 664.050 135.450 671.400 ;
        RECT 136.950 670.950 139.050 673.050 ;
        RECT 136.950 668.850 139.050 669.750 ;
        RECT 122.550 659.700 123.750 663.300 ;
        RECT 133.950 661.950 136.050 664.050 ;
        RECT 143.400 660.600 144.600 677.400 ;
        RECT 187.950 673.950 190.050 676.050 ;
        RECT 193.950 673.950 196.050 676.050 ;
        RECT 208.950 673.950 211.050 676.050 ;
        RECT 181.950 670.950 184.050 673.050 ;
        RECT 185.250 671.250 187.050 672.150 ;
        RECT 187.950 671.850 190.050 672.750 ;
        RECT 190.950 671.250 193.050 672.150 ;
        RECT 194.400 670.050 195.450 673.950 ;
        RECT 181.950 668.850 183.750 669.750 ;
        RECT 184.950 667.950 187.050 670.050 ;
        RECT 190.950 667.950 193.050 670.050 ;
        RECT 193.950 667.950 196.050 670.050 ;
        RECT 191.400 667.050 192.450 667.950 ;
        RECT 187.950 664.950 190.050 667.050 ;
        RECT 190.950 664.950 193.050 667.050 ;
        RECT 121.950 657.600 124.050 659.700 ;
        RECT 142.950 658.500 145.050 660.600 ;
        RECT 145.950 640.950 148.050 643.050 ;
        RECT 113.250 632.250 114.750 633.150 ;
        RECT 115.950 632.400 120.450 633.450 ;
        RECT 115.950 631.950 118.050 632.400 ;
        RECT 109.950 629.850 111.750 630.750 ;
        RECT 112.950 628.950 115.050 631.050 ;
        RECT 116.250 629.850 118.050 630.750 ;
        RECT 113.400 628.050 114.450 628.950 ;
        RECT 103.950 625.950 106.050 628.050 ;
        RECT 112.950 625.950 115.050 628.050 ;
        RECT 119.400 625.050 120.450 632.400 ;
        RECT 146.400 631.050 147.450 640.950 ;
        RECT 184.950 633.450 187.050 634.050 ;
        RECT 188.400 633.450 189.450 664.950 ;
        RECT 191.400 643.050 192.450 664.950 ;
        RECT 190.950 640.950 193.050 643.050 ;
        RECT 182.250 632.250 183.750 633.150 ;
        RECT 184.950 632.400 189.450 633.450 ;
        RECT 184.950 631.950 187.050 632.400 ;
        RECT 145.950 628.950 148.050 631.050 ;
        RECT 178.950 629.850 180.750 630.750 ;
        RECT 181.950 628.950 184.050 631.050 ;
        RECT 185.250 629.850 187.050 630.750 ;
        RECT 142.950 626.250 145.050 627.150 ;
        RECT 145.950 626.850 148.050 627.750 ;
        RECT 118.950 622.950 121.050 625.050 ;
        RECT 142.950 622.950 145.050 625.050 ;
        RECT 103.950 605.400 106.050 607.500 ;
        RECT 94.950 601.950 97.050 604.050 ;
        RECT 95.400 601.050 96.450 601.950 ;
        RECT 88.950 598.950 91.050 601.050 ;
        RECT 94.950 598.950 97.050 601.050 ;
        RECT 88.950 596.850 91.050 597.750 ;
        RECT 94.950 596.850 97.050 597.750 ;
        RECT 104.250 593.400 105.450 605.400 ;
        RECT 106.950 602.250 109.050 603.150 ;
        RECT 109.950 601.950 112.050 604.050 ;
        RECT 139.950 601.950 142.050 604.050 ;
        RECT 160.950 601.950 163.050 604.050 ;
        RECT 181.950 601.950 184.050 604.050 ;
        RECT 106.950 600.450 109.050 601.050 ;
        RECT 110.400 600.450 111.450 601.950 ;
        RECT 106.950 599.400 111.450 600.450 ;
        RECT 139.950 599.850 142.050 600.750 ;
        RECT 106.950 598.950 109.050 599.400 ;
        RECT 142.950 599.250 145.050 600.150 ;
        RECT 142.950 595.950 145.050 598.050 ;
        RECT 143.400 595.050 144.450 595.950 ;
        RECT 103.950 591.300 106.050 593.400 ;
        RECT 142.950 592.950 145.050 595.050 ;
        RECT 82.950 586.500 85.050 588.600 ;
        RECT 104.250 587.700 105.450 591.300 ;
        RECT 103.950 585.600 106.050 587.700 ;
        RECT 151.950 562.950 154.050 565.050 ;
        RECT 152.400 562.050 153.450 562.950 ;
        RECT 151.950 559.950 154.050 562.050 ;
        RECT 157.950 561.450 160.050 562.050 ;
        RECT 161.400 561.450 162.450 601.950 ;
        RECT 175.950 598.950 178.050 601.050 ;
        RECT 179.250 599.250 181.050 600.150 ;
        RECT 181.950 599.850 184.050 600.750 ;
        RECT 184.950 599.250 187.050 600.150 ;
        RECT 175.950 596.850 177.750 597.750 ;
        RECT 178.950 595.950 181.050 598.050 ;
        RECT 184.950 595.950 187.050 598.050 ;
        RECT 185.400 595.050 186.450 595.950 ;
        RECT 184.950 592.950 187.050 595.050 ;
        RECT 155.250 560.250 156.750 561.150 ;
        RECT 157.950 560.400 162.450 561.450 ;
        RECT 157.950 559.950 160.050 560.400 ;
        RECT 112.950 557.250 114.750 558.150 ;
        RECT 115.950 556.950 118.050 559.050 ;
        RECT 121.950 558.450 124.050 559.050 ;
        RECT 121.950 557.400 126.450 558.450 ;
        RECT 121.950 556.950 124.050 557.400 ;
        RECT 70.950 553.950 73.050 556.050 ;
        RECT 74.250 554.250 75.750 555.150 ;
        RECT 76.950 553.950 79.050 556.050 ;
        RECT 79.950 553.950 82.050 556.050 ;
        RECT 112.950 553.950 115.050 556.050 ;
        RECT 116.250 554.850 118.050 555.750 ;
        RECT 118.950 554.250 121.050 555.150 ;
        RECT 121.950 554.850 124.050 555.750 ;
        RECT 77.400 553.050 78.450 553.950 ;
        RECT 73.950 550.950 76.050 553.050 ;
        RECT 76.950 550.950 79.050 553.050 ;
        RECT 118.950 550.950 121.050 553.050 ;
        RECT 74.400 532.050 75.450 550.950 ;
        RECT 67.950 529.950 70.050 532.050 ;
        RECT 73.950 529.950 76.050 532.050 ;
        RECT 28.950 528.450 31.050 529.050 ;
        RECT 26.400 527.400 31.050 528.450 ;
        RECT 26.400 487.050 27.450 527.400 ;
        RECT 28.950 526.950 31.050 527.400 ;
        RECT 34.950 526.950 37.050 529.050 ;
        RECT 37.950 526.950 40.050 529.050 ;
        RECT 64.950 526.950 67.050 529.050 ;
        RECT 28.950 524.850 31.050 525.750 ;
        RECT 31.950 524.250 34.050 525.150 ;
        RECT 31.950 522.450 34.050 523.050 ;
        RECT 35.400 522.450 36.450 526.950 ;
        RECT 65.400 526.050 66.450 526.950 ;
        RECT 37.950 524.850 40.050 525.750 ;
        RECT 64.950 523.950 67.050 526.050 ;
        RECT 68.400 523.050 69.450 529.950 ;
        RECT 70.950 523.950 73.050 526.050 ;
        RECT 74.250 524.250 76.050 525.150 ;
        RECT 31.950 521.400 36.450 522.450 ;
        RECT 64.950 521.850 66.750 522.750 ;
        RECT 31.950 520.950 34.050 521.400 ;
        RECT 67.950 520.950 70.050 523.050 ;
        RECT 71.250 521.850 72.750 522.750 ;
        RECT 73.950 520.950 76.050 523.050 ;
        RECT 67.950 518.850 70.050 519.750 ;
        RECT 74.400 493.050 75.450 520.950 ;
        RECT 73.950 490.950 76.050 493.050 ;
        RECT 77.400 490.050 78.450 550.950 ;
        RECT 125.400 550.050 126.450 557.400 ;
        RECT 127.950 556.950 130.050 559.050 ;
        RECT 151.950 557.850 153.750 558.750 ;
        RECT 154.950 556.950 157.050 559.050 ;
        RECT 158.250 557.850 160.050 558.750 ;
        RECT 112.950 547.950 115.050 550.050 ;
        RECT 124.950 547.950 127.050 550.050 ;
        RECT 113.400 529.050 114.450 547.950 ;
        RECT 115.950 529.950 118.050 532.050 ;
        RECT 106.950 526.950 109.050 529.050 ;
        RECT 110.250 527.250 111.750 528.150 ;
        RECT 112.950 526.950 115.050 529.050 ;
        RECT 116.400 526.050 117.450 529.950 ;
        RECT 79.950 523.950 82.050 526.050 ;
        RECT 106.950 524.850 108.750 525.750 ;
        RECT 109.950 523.950 112.050 526.050 ;
        RECT 113.250 524.850 114.750 525.750 ;
        RECT 115.950 523.950 118.050 526.050 ;
        RECT 76.950 487.950 79.050 490.050 ;
        RECT 25.950 484.950 28.050 487.050 ;
        RECT 28.950 485.250 31.050 486.150 ;
        RECT 34.950 485.850 37.050 486.750 ;
        RECT 37.950 485.250 40.050 486.150 ;
        RECT 70.950 485.250 73.050 486.150 ;
        RECT 76.950 485.250 79.050 486.150 ;
        RECT 28.950 481.950 31.050 484.050 ;
        RECT 37.950 481.950 40.050 484.050 ;
        RECT 70.950 481.950 73.050 484.050 ;
        RECT 74.250 482.250 75.750 483.150 ;
        RECT 76.950 481.950 79.050 484.050 ;
        RECT 29.400 457.050 30.450 481.950 ;
        RECT 71.400 460.050 72.450 481.950 ;
        RECT 73.950 478.950 76.050 481.050 ;
        RECT 31.950 457.950 34.050 460.050 ;
        RECT 70.950 457.950 73.050 460.050 ;
        RECT 73.950 457.950 76.050 460.050 ;
        RECT 77.400 457.050 78.450 481.950 ;
        RECT 80.400 481.050 81.450 523.950 ;
        RECT 110.400 523.050 111.450 523.950 ;
        RECT 109.950 520.950 112.050 523.050 ;
        RECT 115.950 521.850 118.050 522.750 ;
        RECT 82.950 490.950 85.050 493.050 ;
        RECT 79.950 478.950 82.050 481.050 ;
        RECT 28.950 454.950 31.050 457.050 ;
        RECT 32.250 455.850 33.750 456.750 ;
        RECT 37.950 454.950 40.050 457.050 ;
        RECT 70.950 455.250 73.050 456.150 ;
        RECT 73.950 455.850 76.050 456.750 ;
        RECT 76.950 454.950 79.050 457.050 ;
        RECT 28.950 452.850 31.050 453.750 ;
        RECT 34.950 452.850 37.050 453.750 ;
        RECT 7.950 422.400 10.050 424.500 ;
        RECT 28.950 423.300 31.050 425.400 ;
        RECT 8.400 405.600 9.600 422.400 ;
        RECT 29.250 419.700 30.450 423.300 ;
        RECT 28.950 417.600 31.050 419.700 ;
        RECT 13.950 413.250 16.050 414.150 ;
        RECT 19.950 413.250 22.050 414.150 ;
        RECT 13.950 409.950 16.050 412.050 ;
        RECT 19.950 409.950 22.050 412.050 ;
        RECT 7.950 403.500 10.050 405.600 ;
        RECT 7.950 317.400 10.050 319.500 ;
        RECT 8.400 300.600 9.600 317.400 ;
        RECT 20.400 316.050 21.450 409.950 ;
        RECT 29.250 405.600 30.450 417.600 ;
        RECT 38.400 415.050 39.450 454.950 ;
        RECT 70.950 451.950 73.050 454.050 ;
        RECT 83.400 424.050 84.450 490.950 ;
        RECT 106.950 487.950 109.050 490.050 ;
        RECT 109.950 488.250 112.050 489.150 ;
        RECT 107.400 481.050 108.450 487.950 ;
        RECT 109.950 484.950 112.050 487.050 ;
        RECT 113.250 485.250 114.750 486.150 ;
        RECT 115.950 484.950 118.050 487.050 ;
        RECT 119.250 485.250 121.050 486.150 ;
        RECT 110.400 484.050 111.450 484.950 ;
        RECT 109.950 481.950 112.050 484.050 ;
        RECT 112.950 481.950 115.050 484.050 ;
        RECT 116.250 482.850 117.750 483.750 ;
        RECT 118.950 481.950 121.050 484.050 ;
        RECT 106.950 478.950 109.050 481.050 ;
        RECT 107.400 460.050 108.450 478.950 ;
        RECT 113.400 463.050 114.450 481.950 ;
        RECT 119.400 481.050 120.450 481.950 ;
        RECT 118.950 478.950 121.050 481.050 ;
        RECT 112.950 460.950 115.050 463.050 ;
        RECT 118.950 460.950 121.050 463.050 ;
        RECT 106.950 457.950 109.050 460.050 ;
        RECT 103.950 455.250 106.050 456.150 ;
        RECT 106.950 455.850 109.050 456.750 ;
        RECT 112.950 456.450 115.050 457.050 ;
        RECT 109.950 455.250 111.750 456.150 ;
        RECT 112.950 455.400 117.450 456.450 ;
        RECT 112.950 454.950 115.050 455.400 ;
        RECT 103.950 451.950 106.050 454.050 ;
        RECT 109.950 451.950 112.050 454.050 ;
        RECT 113.250 452.850 115.050 453.750 ;
        RECT 82.950 421.950 85.050 424.050 ;
        RECT 106.950 421.950 109.050 424.050 ;
        RECT 31.950 412.950 34.050 415.050 ;
        RECT 37.950 412.950 40.050 415.050 ;
        RECT 46.950 412.950 49.050 415.050 ;
        RECT 67.950 413.250 69.750 414.150 ;
        RECT 70.950 412.950 73.050 415.050 ;
        RECT 76.950 412.950 79.050 415.050 ;
        RECT 32.400 412.050 33.450 412.950 ;
        RECT 31.950 409.950 34.050 412.050 ;
        RECT 31.950 407.850 34.050 408.750 ;
        RECT 28.950 403.500 31.050 405.600 ;
        RECT 31.950 403.950 34.050 406.050 ;
        RECT 32.400 385.050 33.450 403.950 ;
        RECT 38.400 385.050 39.450 412.950 ;
        RECT 47.400 406.050 48.450 412.950 ;
        RECT 67.950 409.950 70.050 412.050 ;
        RECT 71.250 410.850 73.050 411.750 ;
        RECT 73.950 410.250 76.050 411.150 ;
        RECT 76.950 410.850 79.050 411.750 ;
        RECT 73.950 406.950 76.050 409.050 ;
        RECT 46.950 403.950 49.050 406.050 ;
        RECT 31.950 382.950 34.050 385.050 ;
        RECT 35.250 383.250 36.750 384.150 ;
        RECT 37.950 382.950 40.050 385.050 ;
        RECT 28.950 381.450 31.050 382.050 ;
        RECT 26.400 380.400 31.050 381.450 ;
        RECT 32.250 380.850 33.750 381.750 ;
        RECT 26.400 334.050 27.450 380.400 ;
        RECT 28.950 379.950 31.050 380.400 ;
        RECT 34.950 379.950 37.050 382.050 ;
        RECT 38.250 380.850 40.050 381.750 ;
        RECT 70.950 380.250 72.750 381.150 ;
        RECT 73.950 379.950 76.050 382.050 ;
        RECT 77.250 380.250 79.050 381.150 ;
        RECT 28.950 377.850 31.050 378.750 ;
        RECT 35.400 373.050 36.450 379.950 ;
        RECT 70.950 376.950 73.050 379.050 ;
        RECT 74.250 377.850 75.750 378.750 ;
        RECT 76.950 376.950 79.050 379.050 ;
        RECT 71.400 376.050 72.450 376.950 ;
        RECT 83.400 376.050 84.450 421.950 ;
        RECT 103.950 418.950 106.050 421.050 ;
        RECT 85.950 406.950 88.050 409.050 ;
        RECT 70.950 373.950 73.050 376.050 ;
        RECT 82.950 373.950 85.050 376.050 ;
        RECT 86.400 373.050 87.450 406.950 ;
        RECT 104.400 379.050 105.450 418.950 ;
        RECT 107.400 385.050 108.450 421.950 ;
        RECT 116.400 421.050 117.450 455.400 ;
        RECT 115.950 418.950 118.050 421.050 ;
        RECT 109.950 415.950 112.050 418.050 ;
        RECT 115.950 417.450 118.050 418.050 ;
        RECT 119.400 417.450 120.450 460.950 ;
        RECT 124.950 457.950 127.050 460.050 ;
        RECT 125.400 454.050 126.450 457.950 ;
        RECT 124.950 451.950 127.050 454.050 ;
        RECT 113.250 416.250 114.750 417.150 ;
        RECT 115.950 416.400 120.450 417.450 ;
        RECT 115.950 415.950 118.050 416.400 ;
        RECT 109.950 413.850 111.750 414.750 ;
        RECT 112.950 412.950 115.050 415.050 ;
        RECT 116.250 413.850 118.050 414.750 ;
        RECT 128.400 391.050 129.450 556.950 ;
        RECT 155.400 553.050 156.450 556.950 ;
        RECT 154.950 550.950 157.050 553.050 ;
        RECT 154.950 529.950 157.050 532.050 ;
        RECT 151.950 528.450 154.050 529.050 ;
        RECT 149.400 527.400 154.050 528.450 ;
        RECT 155.250 527.850 156.750 528.750 ;
        RECT 157.950 528.450 160.050 529.050 ;
        RECT 161.400 528.450 162.450 560.400 ;
        RECT 188.400 553.050 189.450 632.400 ;
        RECT 194.400 631.050 195.450 667.950 ;
        RECT 209.400 664.050 210.450 673.950 ;
        RECT 215.400 667.050 216.450 694.950 ;
        RECT 229.950 688.950 232.050 691.050 ;
        RECT 220.950 672.450 223.050 673.050 ;
        RECT 218.400 671.400 223.050 672.450 ;
        RECT 218.400 667.050 219.450 671.400 ;
        RECT 220.950 670.950 223.050 671.400 ;
        RECT 224.250 671.250 225.750 672.150 ;
        RECT 226.950 670.950 229.050 673.050 ;
        RECT 230.400 670.050 231.450 688.950 ;
        RECT 233.400 673.050 234.450 697.950 ;
        RECT 263.400 697.050 264.450 700.950 ;
        RECT 265.950 697.950 268.050 700.050 ;
        RECT 269.250 698.850 270.750 699.750 ;
        RECT 271.950 697.950 274.050 700.050 ;
        RECT 262.950 694.950 265.050 697.050 ;
        RECT 235.950 691.950 238.050 694.050 ;
        RECT 232.950 670.950 235.050 673.050 ;
        RECT 236.400 672.450 237.450 691.950 ;
        RECT 241.950 677.400 244.050 679.500 ;
        RECT 262.950 677.400 265.050 679.500 ;
        RECT 238.950 674.250 241.050 675.150 ;
        RECT 238.950 672.450 241.050 673.050 ;
        RECT 236.400 671.400 241.050 672.450 ;
        RECT 238.950 670.950 241.050 671.400 ;
        RECT 220.950 668.850 222.750 669.750 ;
        RECT 223.950 667.950 226.050 670.050 ;
        RECT 227.250 668.850 228.750 669.750 ;
        RECT 229.950 667.950 232.050 670.050 ;
        RECT 238.950 667.950 241.050 670.050 ;
        RECT 214.950 664.950 217.050 667.050 ;
        RECT 217.950 664.950 220.050 667.050 ;
        RECT 229.950 665.850 232.050 666.750 ;
        RECT 208.950 661.950 211.050 664.050 ;
        RECT 193.950 628.950 196.050 631.050 ;
        RECT 193.950 605.400 196.050 607.500 ;
        RECT 194.400 588.600 195.600 605.400 ;
        RECT 199.950 598.950 202.050 601.050 ;
        RECT 205.950 600.450 208.050 601.050 ;
        RECT 209.400 600.450 210.450 661.950 ;
        RECT 220.950 632.250 223.050 633.150 ;
        RECT 232.950 631.950 235.050 634.050 ;
        RECT 211.950 628.950 214.050 631.050 ;
        RECT 220.950 628.950 223.050 631.050 ;
        RECT 224.250 629.250 225.750 630.150 ;
        RECT 226.950 628.950 229.050 631.050 ;
        RECT 230.250 629.250 232.050 630.150 ;
        RECT 212.400 604.050 213.450 628.950 ;
        RECT 221.400 628.050 222.450 628.950 ;
        RECT 220.950 625.950 223.050 628.050 ;
        RECT 223.950 625.950 226.050 628.050 ;
        RECT 227.250 626.850 228.750 627.750 ;
        RECT 229.950 627.450 232.050 628.050 ;
        RECT 233.400 627.450 234.450 631.950 ;
        RECT 239.400 628.050 240.450 667.950 ;
        RECT 242.550 665.400 243.750 677.400 ;
        RECT 250.950 673.950 253.050 676.050 ;
        RECT 251.400 673.050 252.450 673.950 ;
        RECT 250.950 670.950 253.050 673.050 ;
        RECT 256.950 670.950 259.050 673.050 ;
        RECT 250.950 668.850 253.050 669.750 ;
        RECT 256.950 668.850 259.050 669.750 ;
        RECT 241.950 663.300 244.050 665.400 ;
        RECT 242.550 659.700 243.750 663.300 ;
        RECT 263.400 660.600 264.600 677.400 ;
        RECT 266.400 673.050 267.450 697.950 ;
        RECT 265.950 670.950 268.050 673.050 ;
        RECT 241.950 657.600 244.050 659.700 ;
        RECT 262.950 658.500 265.050 660.600 ;
        RECT 266.400 634.050 267.450 670.950 ;
        RECT 272.400 670.050 273.450 697.950 ;
        RECT 275.400 691.050 276.450 700.950 ;
        RECT 304.950 697.950 307.050 700.050 ;
        RECT 343.950 697.950 346.050 700.050 ;
        RECT 352.950 697.950 355.050 700.050 ;
        RECT 385.950 697.950 388.050 700.050 ;
        RECT 389.250 698.250 390.750 699.150 ;
        RECT 418.950 697.950 421.050 700.050 ;
        RECT 424.950 697.950 427.050 700.050 ;
        RECT 305.400 697.050 306.450 697.950 ;
        RECT 304.950 694.950 307.050 697.050 ;
        RECT 274.950 688.950 277.050 691.050 ;
        RECT 277.950 677.400 280.050 679.500 ;
        RECT 298.950 677.400 301.050 679.500 ;
        RECT 274.950 674.250 277.050 675.150 ;
        RECT 274.950 670.950 277.050 673.050 ;
        RECT 271.950 667.950 274.050 670.050 ;
        RECT 278.550 665.400 279.750 677.400 ;
        RECT 286.950 673.950 289.050 676.050 ;
        RECT 287.400 673.050 288.450 673.950 ;
        RECT 286.950 670.950 289.050 673.050 ;
        RECT 292.950 670.950 295.050 673.050 ;
        RECT 286.950 668.850 289.050 669.750 ;
        RECT 292.950 668.850 295.050 669.750 ;
        RECT 277.950 663.300 280.050 665.400 ;
        RECT 278.550 659.700 279.750 663.300 ;
        RECT 299.400 660.600 300.600 677.400 ;
        RECT 305.400 676.050 306.450 694.950 ;
        RECT 353.400 676.050 354.450 697.950 ;
        RECT 388.950 694.950 391.050 697.050 ;
        RECT 304.950 673.950 307.050 676.050 ;
        RECT 343.950 673.950 346.050 676.050 ;
        RECT 352.950 673.950 355.050 676.050 ;
        RECT 370.950 673.950 373.050 676.050 ;
        RECT 389.400 675.450 390.450 694.950 ;
        RECT 389.400 674.400 393.450 675.450 ;
        RECT 337.950 670.950 340.050 673.050 ;
        RECT 341.250 671.250 343.050 672.150 ;
        RECT 343.950 671.850 346.050 672.750 ;
        RECT 346.950 671.250 349.050 672.150 ;
        RECT 337.950 668.850 339.750 669.750 ;
        RECT 340.950 667.950 343.050 670.050 ;
        RECT 346.950 667.950 349.050 670.050 ;
        RECT 277.950 657.600 280.050 659.700 ;
        RECT 298.950 658.500 301.050 660.600 ;
        RECT 298.950 649.950 301.050 652.050 ;
        RECT 263.250 632.250 264.750 633.150 ;
        RECT 265.950 631.950 268.050 634.050 ;
        RECT 259.950 629.850 261.750 630.750 ;
        RECT 262.950 628.950 265.050 631.050 ;
        RECT 266.250 629.850 268.050 630.750 ;
        RECT 295.950 630.450 298.050 631.050 ;
        RECT 299.400 630.450 300.450 649.950 ;
        RECT 337.950 632.250 340.050 633.150 ;
        RECT 295.950 629.400 300.450 630.450 ;
        RECT 295.950 628.950 298.050 629.400 ;
        RECT 229.950 626.400 234.450 627.450 ;
        RECT 229.950 625.950 232.050 626.400 ;
        RECT 238.950 625.950 241.050 628.050 ;
        RECT 214.950 605.400 217.050 607.500 ;
        RECT 211.950 601.950 214.050 604.050 ;
        RECT 205.950 599.400 210.450 600.450 ;
        RECT 205.950 598.950 208.050 599.400 ;
        RECT 199.950 596.850 202.050 597.750 ;
        RECT 205.950 596.850 208.050 597.750 ;
        RECT 202.950 592.950 205.050 595.050 ;
        RECT 193.950 586.500 196.050 588.600 ;
        RECT 193.950 554.850 196.050 555.750 ;
        RECT 187.950 550.950 190.050 553.050 ;
        RECT 193.950 550.950 196.050 553.050 ;
        RECT 194.400 529.050 195.450 550.950 ;
        RECT 149.400 487.050 150.450 527.400 ;
        RECT 151.950 526.950 154.050 527.400 ;
        RECT 157.950 527.400 162.450 528.450 ;
        RECT 157.950 526.950 160.050 527.400 ;
        RECT 151.950 524.850 154.050 525.750 ;
        RECT 157.950 524.850 160.050 525.750 ;
        RECT 161.400 508.050 162.450 527.400 ;
        RECT 187.950 526.950 190.050 529.050 ;
        RECT 193.950 526.950 196.050 529.050 ;
        RECT 187.950 524.850 190.050 525.750 ;
        RECT 193.950 524.850 196.050 525.750 ;
        RECT 160.950 505.950 163.050 508.050 ;
        RECT 148.950 484.950 151.050 487.050 ;
        RECT 151.950 485.250 154.050 486.150 ;
        RECT 157.950 485.250 160.050 486.150 ;
        RECT 187.950 485.250 190.050 486.150 ;
        RECT 193.950 485.250 196.050 486.150 ;
        RECT 151.950 481.950 154.050 484.050 ;
        RECT 155.250 482.250 156.750 483.150 ;
        RECT 157.950 481.950 160.050 484.050 ;
        RECT 193.950 481.950 196.050 484.050 ;
        RECT 158.400 481.050 159.450 481.950 ;
        RECT 194.400 481.050 195.450 481.950 ;
        RECT 154.950 478.950 157.050 481.050 ;
        RECT 157.950 478.950 160.050 481.050 ;
        RECT 193.950 478.950 196.050 481.050 ;
        RECT 130.950 457.950 133.050 460.050 ;
        RECT 151.950 457.950 154.050 460.050 ;
        RECT 131.400 418.050 132.450 457.950 ;
        RECT 152.400 457.050 153.450 457.950 ;
        RECT 145.950 454.950 148.050 457.050 ;
        RECT 149.250 455.250 150.750 456.150 ;
        RECT 151.950 454.950 154.050 457.050 ;
        RECT 155.400 454.050 156.450 478.950 ;
        RECT 190.950 455.250 193.050 456.150 ;
        RECT 145.950 452.850 147.750 453.750 ;
        RECT 148.950 451.950 151.050 454.050 ;
        RECT 152.250 452.850 153.750 453.750 ;
        RECT 154.950 451.950 157.050 454.050 ;
        RECT 154.950 449.850 157.050 450.750 ;
        RECT 160.950 422.400 163.050 424.500 ;
        RECT 181.950 423.300 184.050 425.400 ;
        RECT 130.950 415.950 133.050 418.050 ;
        RECT 145.950 413.250 148.050 414.150 ;
        RECT 151.950 413.250 154.050 414.150 ;
        RECT 145.950 409.950 148.050 412.050 ;
        RECT 151.950 409.950 154.050 412.050 ;
        RECT 146.400 409.050 147.450 409.950 ;
        RECT 145.950 406.950 148.050 409.050 ;
        RECT 152.400 406.050 153.450 409.950 ;
        RECT 151.950 403.950 154.050 406.050 ;
        RECT 161.400 405.600 162.600 422.400 ;
        RECT 182.250 419.700 183.450 423.300 ;
        RECT 181.950 417.600 184.050 419.700 ;
        RECT 166.950 413.250 169.050 414.150 ;
        RECT 172.950 413.250 175.050 414.150 ;
        RECT 166.950 409.950 169.050 412.050 ;
        RECT 172.950 409.950 175.050 412.050 ;
        RECT 160.950 403.500 163.050 405.600 ;
        RECT 167.400 397.050 168.450 409.950 ;
        RECT 166.950 394.950 169.050 397.050 ;
        RECT 127.950 388.950 130.050 391.050 ;
        RECT 151.950 388.950 154.050 391.050 ;
        RECT 152.400 385.050 153.450 388.950 ;
        RECT 106.950 382.950 109.050 385.050 ;
        RECT 115.950 382.950 118.050 385.050 ;
        RECT 121.950 382.950 124.050 385.050 ;
        RECT 151.950 382.950 154.050 385.050 ;
        RECT 155.250 383.250 157.050 384.150 ;
        RECT 106.950 380.850 109.050 381.750 ;
        RECT 112.950 380.250 115.050 381.150 ;
        RECT 115.950 380.850 118.050 381.750 ;
        RECT 103.950 376.950 106.050 379.050 ;
        RECT 112.950 376.950 115.050 379.050 ;
        RECT 34.950 370.950 37.050 373.050 ;
        RECT 85.950 370.950 88.050 373.050 ;
        RECT 86.400 343.050 87.450 370.950 ;
        RECT 103.950 350.400 106.050 352.500 ;
        RECT 91.950 344.250 94.050 345.150 ;
        RECT 49.950 342.450 52.050 343.050 ;
        RECT 49.950 341.400 54.450 342.450 ;
        RECT 49.950 340.950 52.050 341.400 ;
        RECT 53.400 340.050 54.450 341.400 ;
        RECT 73.950 340.950 76.050 343.050 ;
        RECT 82.950 341.250 84.750 342.150 ;
        RECT 85.950 340.950 88.050 343.050 ;
        RECT 89.250 341.250 90.750 342.150 ;
        RECT 91.950 340.950 94.050 343.050 ;
        RECT 28.950 338.850 31.050 339.750 ;
        RECT 49.950 338.850 52.050 339.750 ;
        RECT 52.950 337.950 55.050 340.050 ;
        RECT 25.950 331.950 28.050 334.050 ;
        RECT 28.950 317.400 31.050 319.500 ;
        RECT 43.950 317.400 46.050 319.500 ;
        RECT 19.950 313.950 22.050 316.050 ;
        RECT 20.400 313.050 21.450 313.950 ;
        RECT 13.950 312.450 16.050 313.050 ;
        RECT 13.950 311.400 18.450 312.450 ;
        RECT 13.950 310.950 16.050 311.400 ;
        RECT 13.950 308.850 16.050 309.750 ;
        RECT 7.950 298.500 10.050 300.600 ;
        RECT 17.400 268.050 18.450 311.400 ;
        RECT 19.950 310.950 22.050 313.050 ;
        RECT 19.950 308.850 22.050 309.750 ;
        RECT 29.250 305.400 30.450 317.400 ;
        RECT 31.950 314.250 34.050 315.150 ;
        RECT 40.950 314.250 43.050 315.150 ;
        RECT 31.950 310.950 34.050 313.050 ;
        RECT 40.950 310.950 43.050 313.050 ;
        RECT 28.950 303.300 31.050 305.400 ;
        RECT 29.250 299.700 30.450 303.300 ;
        RECT 28.950 297.600 31.050 299.700 ;
        RECT 32.400 295.050 33.450 310.950 ;
        RECT 41.400 310.050 42.450 310.950 ;
        RECT 40.950 307.950 43.050 310.050 ;
        RECT 31.950 292.950 34.050 295.050 ;
        RECT 41.400 280.050 42.450 307.950 ;
        RECT 44.550 305.400 45.750 317.400 ;
        RECT 53.400 316.050 54.450 337.950 ;
        RECT 64.950 317.400 67.050 319.500 ;
        RECT 52.950 313.950 55.050 316.050 ;
        RECT 53.400 313.050 54.450 313.950 ;
        RECT 52.950 310.950 55.050 313.050 ;
        RECT 58.950 310.950 61.050 313.050 ;
        RECT 52.950 308.850 55.050 309.750 ;
        RECT 58.950 308.850 61.050 309.750 ;
        RECT 43.950 303.300 46.050 305.400 ;
        RECT 44.550 299.700 45.750 303.300 ;
        RECT 65.400 300.600 66.600 317.400 ;
        RECT 43.950 297.600 46.050 299.700 ;
        RECT 64.950 298.500 67.050 300.600 ;
        RECT 43.950 292.950 46.050 295.050 ;
        RECT 40.950 277.950 43.050 280.050 ;
        RECT 34.950 271.950 37.050 274.050 ;
        RECT 35.400 271.050 36.450 271.950 ;
        RECT 31.950 269.250 33.750 270.150 ;
        RECT 34.950 268.950 37.050 271.050 ;
        RECT 40.950 268.950 43.050 271.050 ;
        RECT 44.400 268.050 45.450 292.950 ;
        RECT 46.950 277.950 49.050 280.050 ;
        RECT 16.950 265.950 19.050 268.050 ;
        RECT 31.950 265.950 34.050 268.050 ;
        RECT 35.250 266.850 37.050 267.750 ;
        RECT 37.950 266.250 40.050 267.150 ;
        RECT 40.950 266.850 43.050 267.750 ;
        RECT 43.950 265.950 46.050 268.050 ;
        RECT 37.950 264.450 40.050 265.050 ;
        RECT 35.400 263.400 40.050 264.450 ;
        RECT 35.400 238.050 36.450 263.400 ;
        RECT 37.950 262.950 40.050 263.400 ;
        RECT 31.950 236.250 33.750 237.150 ;
        RECT 34.950 235.950 37.050 238.050 ;
        RECT 38.250 236.250 40.050 237.150 ;
        RECT 31.950 232.950 34.050 235.050 ;
        RECT 35.250 233.850 36.750 234.750 ;
        RECT 37.950 232.950 40.050 235.050 ;
        RECT 32.400 232.050 33.450 232.950 ;
        RECT 31.950 229.950 34.050 232.050 ;
        RECT 28.950 197.250 31.050 198.150 ;
        RECT 34.950 197.250 37.050 198.150 ;
        RECT 32.250 194.250 33.750 195.150 ;
        RECT 34.950 193.950 37.050 196.050 ;
        RECT 40.950 193.950 43.050 196.050 ;
        RECT 31.950 190.950 34.050 193.050 ;
        RECT 31.950 187.950 34.050 190.050 ;
        RECT 32.400 169.050 33.450 187.950 ;
        RECT 41.400 169.050 42.450 193.950 ;
        RECT 31.950 166.950 34.050 169.050 ;
        RECT 40.950 166.950 43.050 169.050 ;
        RECT 31.950 164.850 34.050 165.750 ;
        RECT 34.950 164.250 37.050 165.150 ;
        RECT 40.950 164.850 43.050 165.750 ;
        RECT 44.400 147.450 45.450 265.950 ;
        RECT 47.400 196.050 48.450 277.950 ;
        RECT 74.400 274.050 75.450 340.950 ;
        RECT 82.950 337.950 85.050 340.050 ;
        RECT 86.250 338.850 87.750 339.750 ;
        RECT 88.950 337.950 91.050 340.050 ;
        RECT 83.400 310.050 84.450 337.950 ;
        RECT 89.400 310.050 90.450 337.950 ;
        RECT 92.400 334.050 93.450 340.950 ;
        RECT 91.950 331.950 94.050 334.050 ;
        RECT 104.400 333.600 105.600 350.400 ;
        RECT 106.950 340.950 109.050 343.050 ;
        RECT 109.950 341.250 112.050 342.150 ;
        RECT 115.950 341.250 118.050 342.150 ;
        RECT 82.950 307.950 85.050 310.050 ;
        RECT 88.950 307.950 91.050 310.050 ;
        RECT 73.950 271.950 76.050 274.050 ;
        RECT 79.950 272.250 82.050 273.150 ;
        RECT 74.400 271.050 75.450 271.950 ;
        RECT 92.400 271.050 93.450 331.950 ;
        RECT 103.950 331.500 106.050 333.600 ;
        RECT 107.400 315.450 108.450 340.950 ;
        RECT 109.950 337.950 112.050 340.050 ;
        RECT 115.950 337.950 118.050 340.050 ;
        RECT 110.400 319.050 111.450 337.950 ;
        RECT 109.950 316.950 112.050 319.050 ;
        RECT 109.950 315.450 112.050 316.050 ;
        RECT 107.400 314.400 112.050 315.450 ;
        RECT 109.950 313.950 112.050 314.400 ;
        RECT 103.950 310.950 106.050 313.050 ;
        RECT 107.250 311.250 109.050 312.150 ;
        RECT 109.950 311.850 112.050 312.750 ;
        RECT 112.950 311.250 115.050 312.150 ;
        RECT 103.950 308.850 105.750 309.750 ;
        RECT 106.950 307.950 109.050 310.050 ;
        RECT 112.950 309.450 115.050 310.050 ;
        RECT 110.400 308.400 115.050 309.450 ;
        RECT 70.950 269.250 72.750 270.150 ;
        RECT 73.950 268.950 76.050 271.050 ;
        RECT 77.250 269.250 78.750 270.150 ;
        RECT 79.950 268.950 82.050 271.050 ;
        RECT 91.950 268.950 94.050 271.050 ;
        RECT 70.950 265.950 73.050 268.050 ;
        RECT 74.250 266.850 75.750 267.750 ;
        RECT 76.950 265.950 79.050 268.050 ;
        RECT 73.950 262.950 76.050 265.050 ;
        RECT 74.400 244.050 75.450 262.950 ;
        RECT 73.950 241.950 76.050 244.050 ;
        RECT 64.950 238.950 67.050 241.050 ;
        RECT 70.950 238.950 73.050 241.050 ;
        RECT 74.250 239.850 75.750 240.750 ;
        RECT 76.950 238.950 79.050 241.050 ;
        RECT 79.950 238.950 82.050 241.050 ;
        RECT 65.400 232.050 66.450 238.950 ;
        RECT 70.950 236.850 73.050 237.750 ;
        RECT 76.950 236.850 79.050 237.750 ;
        RECT 80.400 235.050 81.450 238.950 ;
        RECT 110.400 238.050 111.450 308.400 ;
        RECT 112.950 307.950 115.050 308.400 ;
        RECT 112.950 269.250 115.050 270.150 ;
        RECT 118.950 269.250 121.050 270.150 ;
        RECT 112.950 265.950 115.050 268.050 ;
        RECT 116.250 266.250 117.750 267.150 ;
        RECT 118.950 265.950 121.050 268.050 ;
        RECT 113.400 265.050 114.450 265.950 ;
        RECT 119.400 265.050 120.450 265.950 ;
        RECT 112.950 262.950 115.050 265.050 ;
        RECT 115.950 262.950 118.050 265.050 ;
        RECT 118.950 262.950 121.050 265.050 ;
        RECT 116.400 262.050 117.450 262.950 ;
        RECT 115.950 259.950 118.050 262.050 ;
        RECT 106.950 236.250 108.750 237.150 ;
        RECT 109.950 235.950 112.050 238.050 ;
        RECT 113.250 236.250 115.050 237.150 ;
        RECT 115.950 235.950 118.050 238.050 ;
        RECT 79.950 232.950 82.050 235.050 ;
        RECT 106.950 232.950 109.050 235.050 ;
        RECT 110.250 233.850 111.750 234.750 ;
        RECT 112.950 234.450 115.050 235.050 ;
        RECT 116.400 234.450 117.450 235.950 ;
        RECT 112.950 233.400 117.450 234.450 ;
        RECT 112.950 232.950 115.050 233.400 ;
        RECT 64.950 229.950 67.050 232.050 ;
        RECT 46.950 193.950 49.050 196.050 ;
        RECT 65.400 187.050 66.450 229.950 ;
        RECT 107.400 208.050 108.450 232.950 ;
        RECT 122.400 208.050 123.450 382.950 ;
        RECT 151.950 380.850 153.750 381.750 ;
        RECT 154.950 379.950 157.050 382.050 ;
        RECT 163.950 379.950 166.050 382.050 ;
        RECT 124.950 351.300 127.050 353.400 ;
        RECT 155.400 352.050 156.450 379.950 ;
        RECT 125.250 347.700 126.450 351.300 ;
        RECT 145.950 349.950 148.050 352.050 ;
        RECT 154.950 349.950 157.050 352.050 ;
        RECT 124.950 345.600 127.050 347.700 ;
        RECT 125.250 333.600 126.450 345.600 ;
        RECT 127.950 339.450 130.050 340.050 ;
        RECT 127.950 338.400 132.450 339.450 ;
        RECT 127.950 337.950 130.050 338.400 ;
        RECT 131.400 337.050 132.450 338.400 ;
        RECT 142.950 337.950 145.050 340.050 ;
        RECT 127.950 335.850 130.050 336.750 ;
        RECT 130.950 334.950 133.050 337.050 ;
        RECT 124.950 331.500 127.050 333.600 ;
        RECT 127.950 278.400 130.050 280.500 ;
        RECT 128.400 261.600 129.600 278.400 ;
        RECT 143.400 277.050 144.450 337.950 ;
        RECT 146.400 334.050 147.450 349.950 ;
        RECT 160.950 340.950 163.050 343.050 ;
        RECT 157.950 338.250 160.050 339.150 ;
        RECT 160.950 338.850 163.050 339.750 ;
        RECT 157.950 334.950 160.050 337.050 ;
        RECT 145.950 331.950 148.050 334.050 ;
        RECT 146.400 313.050 147.450 331.950 ;
        RECT 145.950 310.950 148.050 313.050 ;
        RECT 145.950 308.850 148.050 309.750 ;
        RECT 151.950 308.850 154.050 309.750 ;
        RECT 148.950 279.300 151.050 281.400 ;
        RECT 142.950 274.950 145.050 277.050 ;
        RECT 149.250 275.700 150.450 279.300 ;
        RECT 133.950 269.250 136.050 270.150 ;
        RECT 139.950 269.250 142.050 270.150 ;
        RECT 133.950 265.950 136.050 268.050 ;
        RECT 136.950 265.950 139.050 268.050 ;
        RECT 139.950 267.450 142.050 268.050 ;
        RECT 143.400 267.450 144.450 274.950 ;
        RECT 148.950 273.600 151.050 275.700 ;
        RECT 139.950 266.400 144.450 267.450 ;
        RECT 139.950 265.950 142.050 266.400 ;
        RECT 134.400 262.050 135.450 265.950 ;
        RECT 127.950 259.500 130.050 261.600 ;
        RECT 133.950 259.950 136.050 262.050 ;
        RECT 100.950 205.950 103.050 208.050 ;
        RECT 106.950 205.950 109.050 208.050 ;
        RECT 115.950 205.950 118.050 208.050 ;
        RECT 121.950 205.950 124.050 208.050 ;
        RECT 67.950 197.250 70.050 198.150 ;
        RECT 73.950 197.250 76.050 198.150 ;
        RECT 97.950 196.950 100.050 199.050 ;
        RECT 67.950 193.950 70.050 196.050 ;
        RECT 71.250 194.250 72.750 195.150 ;
        RECT 73.950 193.950 76.050 196.050 ;
        RECT 68.400 190.050 69.450 193.950 ;
        RECT 74.400 193.050 75.450 193.950 ;
        RECT 98.400 193.050 99.450 196.950 ;
        RECT 101.400 196.050 102.450 205.950 ;
        RECT 112.950 200.250 115.050 201.150 ;
        RECT 103.950 197.250 105.750 198.150 ;
        RECT 106.950 196.950 109.050 199.050 ;
        RECT 112.950 198.450 115.050 199.050 ;
        RECT 116.400 198.450 117.450 205.950 ;
        RECT 118.950 202.950 121.050 205.050 ;
        RECT 110.250 197.250 111.750 198.150 ;
        RECT 112.950 197.400 117.450 198.450 ;
        RECT 112.950 196.950 115.050 197.400 ;
        RECT 100.950 193.950 103.050 196.050 ;
        RECT 103.950 193.950 106.050 196.050 ;
        RECT 107.250 194.850 108.750 195.750 ;
        RECT 109.950 193.950 112.050 196.050 ;
        RECT 70.950 190.950 73.050 193.050 ;
        RECT 73.950 190.950 76.050 193.050 ;
        RECT 97.950 190.950 100.050 193.050 ;
        RECT 67.950 187.950 70.050 190.050 ;
        RECT 64.950 184.950 67.050 187.050 ;
        RECT 68.400 166.050 69.450 187.950 ;
        RECT 71.400 172.050 72.450 190.950 ;
        RECT 104.400 190.050 105.450 193.950 ;
        RECT 103.950 187.950 106.050 190.050 ;
        RECT 73.950 184.950 76.050 187.050 ;
        RECT 70.950 169.950 73.050 172.050 ;
        RECT 74.400 169.050 75.450 184.950 ;
        RECT 119.400 175.050 120.450 202.950 ;
        RECT 79.950 172.950 82.050 175.050 ;
        RECT 112.950 172.950 115.050 175.050 ;
        RECT 118.950 172.950 121.050 175.050 ;
        RECT 121.950 172.950 124.050 175.050 ;
        RECT 80.400 172.050 81.450 172.950 ;
        RECT 79.950 169.950 82.050 172.050 ;
        RECT 85.950 169.950 88.050 172.050 ;
        RECT 73.950 166.950 76.050 169.050 ;
        RECT 77.250 167.250 79.050 168.150 ;
        RECT 79.950 167.850 82.050 168.750 ;
        RECT 82.950 167.250 85.050 168.150 ;
        RECT 67.950 163.950 70.050 166.050 ;
        RECT 73.950 164.850 75.750 165.750 ;
        RECT 76.950 163.950 79.050 166.050 ;
        RECT 82.950 165.450 85.050 166.050 ;
        RECT 86.400 165.450 87.450 169.950 ;
        RECT 113.400 169.050 114.450 172.950 ;
        RECT 122.400 169.050 123.450 172.950 ;
        RECT 112.950 166.950 115.050 169.050 ;
        RECT 121.950 166.950 124.050 169.050 ;
        RECT 82.950 164.400 87.450 165.450 ;
        RECT 112.950 164.850 115.050 165.750 ;
        RECT 82.950 163.950 85.050 164.400 ;
        RECT 118.950 164.250 121.050 165.150 ;
        RECT 121.950 164.850 124.050 165.750 ;
        RECT 41.400 146.400 45.450 147.450 ;
        RECT 31.950 125.250 34.050 126.150 ;
        RECT 37.950 125.250 40.050 126.150 ;
        RECT 31.950 123.450 34.050 124.050 ;
        RECT 29.400 122.400 34.050 123.450 ;
        RECT 29.400 100.050 30.450 122.400 ;
        RECT 31.950 121.950 34.050 122.400 ;
        RECT 35.250 122.250 36.750 123.150 ;
        RECT 37.950 121.950 40.050 124.050 ;
        RECT 34.950 118.950 37.050 121.050 ;
        RECT 35.400 118.050 36.450 118.950 ;
        RECT 34.950 115.950 37.050 118.050 ;
        RECT 28.950 97.950 31.050 100.050 ;
        RECT 29.400 97.050 30.450 97.950 ;
        RECT 28.950 94.950 31.050 97.050 ;
        RECT 37.950 96.450 40.050 97.050 ;
        RECT 41.400 96.450 42.450 146.400 ;
        RECT 68.400 121.050 69.450 163.950 ;
        RECT 118.950 160.950 121.050 163.050 ;
        RECT 109.950 128.250 112.050 129.150 ;
        RECT 70.950 124.950 73.050 127.050 ;
        RECT 100.950 125.250 102.750 126.150 ;
        RECT 103.950 124.950 106.050 127.050 ;
        RECT 109.950 126.450 112.050 127.050 ;
        RECT 107.250 125.250 108.750 126.150 ;
        RECT 109.950 125.400 114.450 126.450 ;
        RECT 109.950 124.950 112.050 125.400 ;
        RECT 70.950 122.850 73.050 123.750 ;
        RECT 73.950 122.250 76.050 123.150 ;
        RECT 100.950 121.950 103.050 124.050 ;
        RECT 104.250 122.850 105.750 123.750 ;
        RECT 106.950 121.950 109.050 124.050 ;
        RECT 67.950 118.950 70.050 121.050 ;
        RECT 73.950 118.950 76.050 121.050 ;
        RECT 68.400 100.050 69.450 118.950 ;
        RECT 67.950 97.950 70.050 100.050 ;
        RECT 37.950 95.400 42.450 96.450 ;
        RECT 37.950 94.950 40.050 95.400 ;
        RECT 28.950 92.850 31.050 93.750 ;
        RECT 31.950 92.250 34.050 93.150 ;
        RECT 37.950 92.850 40.050 93.750 ;
        RECT 31.950 53.250 34.050 54.150 ;
        RECT 37.950 53.250 40.050 54.150 ;
        RECT 37.950 51.450 40.050 52.050 ;
        RECT 41.400 51.450 42.450 95.400 ;
        RECT 64.950 95.250 67.050 96.150 ;
        RECT 67.950 95.850 70.050 96.750 ;
        RECT 70.950 95.250 72.750 96.150 ;
        RECT 73.950 94.950 76.050 97.050 ;
        RECT 64.950 91.950 67.050 94.050 ;
        RECT 70.950 91.950 73.050 94.050 ;
        RECT 74.250 92.850 76.050 93.750 ;
        RECT 65.400 91.050 66.450 91.950 ;
        RECT 64.950 88.950 67.050 91.050 ;
        RECT 70.950 88.950 73.050 91.050 ;
        RECT 71.400 55.050 72.450 88.950 ;
        RECT 70.950 52.950 73.050 55.050 ;
        RECT 35.250 50.250 36.750 51.150 ;
        RECT 37.950 50.400 42.450 51.450 ;
        RECT 37.950 49.950 40.050 50.400 ;
        RECT 67.950 50.250 70.050 51.150 ;
        RECT 70.950 50.850 73.050 51.750 ;
        RECT 101.400 49.050 102.450 121.950 ;
        RECT 106.950 97.950 109.050 100.050 ;
        RECT 106.950 95.850 109.050 96.750 ;
        RECT 109.950 95.250 112.050 96.150 ;
        RECT 109.950 93.450 112.050 94.050 ;
        RECT 113.400 93.450 114.450 125.400 ;
        RECT 119.400 118.050 120.450 160.950 ;
        RECT 124.950 130.950 127.050 133.050 ;
        RECT 125.400 124.050 126.450 130.950 ;
        RECT 124.950 121.950 127.050 124.050 ;
        RECT 118.950 115.950 121.050 118.050 ;
        RECT 109.950 92.400 114.450 93.450 ;
        RECT 109.950 91.950 112.050 92.400 ;
        RECT 103.950 55.950 106.050 58.050 ;
        RECT 104.400 55.050 105.450 55.950 ;
        RECT 103.950 52.950 106.050 55.050 ;
        RECT 109.950 53.250 112.050 54.150 ;
        RECT 103.950 50.850 106.050 51.750 ;
        RECT 113.250 50.250 115.050 51.150 ;
        RECT 34.950 46.950 37.050 49.050 ;
        RECT 67.950 46.950 70.050 49.050 ;
        RECT 100.950 46.950 103.050 49.050 ;
        RECT 112.950 46.950 115.050 49.050 ;
        RECT 113.400 46.050 114.450 46.950 ;
        RECT 137.400 46.050 138.450 265.950 ;
        RECT 149.250 261.600 150.450 273.600 ;
        RECT 151.950 265.950 154.050 268.050 ;
        RECT 151.950 263.850 154.050 264.750 ;
        RECT 148.950 259.500 151.050 261.600 ;
        RECT 139.950 238.950 142.050 241.050 ;
        RECT 140.400 202.050 141.450 238.950 ;
        RECT 142.950 236.250 144.750 237.150 ;
        RECT 145.950 235.950 148.050 238.050 ;
        RECT 149.250 236.250 151.050 237.150 ;
        RECT 164.400 235.050 165.450 379.950 ;
        RECT 173.400 340.050 174.450 409.950 ;
        RECT 182.250 405.600 183.450 417.600 ;
        RECT 184.950 409.950 187.050 412.050 ;
        RECT 184.950 407.850 187.050 408.750 ;
        RECT 181.950 403.500 184.050 405.600 ;
        RECT 190.950 394.950 193.050 397.050 ;
        RECT 187.950 388.950 190.050 391.050 ;
        RECT 188.400 385.050 189.450 388.950 ;
        RECT 191.400 388.050 192.450 394.950 ;
        RECT 203.400 388.050 204.450 592.950 ;
        RECT 209.400 583.050 210.450 599.400 ;
        RECT 215.250 593.400 216.450 605.400 ;
        RECT 217.950 602.250 220.050 603.150 ;
        RECT 217.950 598.950 220.050 601.050 ;
        RECT 214.950 591.300 217.050 593.400 ;
        RECT 215.250 587.700 216.450 591.300 ;
        RECT 214.950 585.600 217.050 587.700 ;
        RECT 208.950 580.950 211.050 583.050 ;
        RECT 214.950 580.950 217.050 583.050 ;
        RECT 215.400 559.050 216.450 580.950 ;
        RECT 214.950 556.950 217.050 559.050 ;
        RECT 214.950 554.850 217.050 555.750 ;
        RECT 218.400 550.050 219.450 598.950 ;
        RECT 217.950 547.950 220.050 550.050 ;
        RECT 221.400 547.050 222.450 625.950 ;
        RECT 224.400 598.050 225.450 625.950 ;
        RECT 263.400 607.050 264.450 628.950 ;
        RECT 295.950 626.850 298.050 627.750 ;
        RECT 262.950 604.950 265.050 607.050 ;
        RECT 259.950 601.950 262.050 604.050 ;
        RECT 253.950 598.950 256.050 601.050 ;
        RECT 257.250 599.250 259.050 600.150 ;
        RECT 259.950 599.850 262.050 600.750 ;
        RECT 262.950 599.250 265.050 600.150 ;
        RECT 299.400 598.050 300.450 629.400 ;
        RECT 301.950 629.250 304.050 630.150 ;
        RECT 307.950 628.950 310.050 631.050 ;
        RECT 337.950 628.950 340.050 631.050 ;
        RECT 341.250 629.250 342.750 630.150 ;
        RECT 343.950 628.950 346.050 631.050 ;
        RECT 347.250 629.250 349.050 630.150 ;
        RECT 301.950 625.950 304.050 628.050 ;
        RECT 305.250 626.250 307.050 627.150 ;
        RECT 304.950 624.450 307.050 625.050 ;
        RECT 308.400 624.450 309.450 628.950 ;
        RECT 304.950 623.400 309.450 624.450 ;
        RECT 304.950 622.950 307.050 623.400 ;
        RECT 338.400 607.050 339.450 628.950 ;
        RECT 340.950 625.950 343.050 628.050 ;
        RECT 344.250 626.850 345.750 627.750 ;
        RECT 346.950 625.950 349.050 628.050 ;
        RECT 341.400 607.050 342.450 625.950 ;
        RECT 304.950 604.950 307.050 607.050 ;
        RECT 337.950 604.950 340.050 607.050 ;
        RECT 340.950 604.950 343.050 607.050 ;
        RECT 346.950 604.950 349.050 607.050 ;
        RECT 305.400 598.050 306.450 604.950 ;
        RECT 334.950 601.950 337.050 604.050 ;
        RECT 340.950 601.950 343.050 604.050 ;
        RECT 335.400 601.050 336.450 601.950 ;
        RECT 334.950 598.950 337.050 601.050 ;
        RECT 338.250 599.250 340.050 600.150 ;
        RECT 340.950 599.850 343.050 600.750 ;
        RECT 343.950 599.250 346.050 600.150 ;
        RECT 223.950 595.950 226.050 598.050 ;
        RECT 253.950 596.850 255.750 597.750 ;
        RECT 256.950 597.450 259.050 598.050 ;
        RECT 256.950 596.400 261.450 597.450 ;
        RECT 256.950 595.950 259.050 596.400 ;
        RECT 256.950 560.250 259.050 561.150 ;
        RECT 232.950 556.950 235.050 559.050 ;
        RECT 247.950 557.250 249.750 558.150 ;
        RECT 250.950 556.950 253.050 559.050 ;
        RECT 254.250 557.250 255.750 558.150 ;
        RECT 256.950 556.950 259.050 559.050 ;
        RECT 220.950 544.950 223.050 547.050 ;
        RECT 233.400 529.050 234.450 556.950 ;
        RECT 247.950 553.950 250.050 556.050 ;
        RECT 251.250 554.850 252.750 555.750 ;
        RECT 253.950 553.950 256.050 556.050 ;
        RECT 248.400 550.050 249.450 553.950 ;
        RECT 247.950 547.950 250.050 550.050 ;
        RECT 257.400 547.050 258.450 556.950 ;
        RECT 260.400 556.050 261.450 596.400 ;
        RECT 262.950 595.950 265.050 598.050 ;
        RECT 295.950 596.250 297.750 597.150 ;
        RECT 298.950 595.950 301.050 598.050 ;
        RECT 304.950 595.950 307.050 598.050 ;
        RECT 334.950 596.850 336.750 597.750 ;
        RECT 337.950 595.950 340.050 598.050 ;
        RECT 343.950 597.450 346.050 598.050 ;
        RECT 347.400 597.450 348.450 604.950 ;
        RECT 343.950 596.400 348.450 597.450 ;
        RECT 343.950 595.950 346.050 596.400 ;
        RECT 263.400 595.050 264.450 595.950 ;
        RECT 262.950 592.950 265.050 595.050 ;
        RECT 295.950 592.950 298.050 595.050 ;
        RECT 299.250 593.850 300.750 594.750 ;
        RECT 301.950 592.950 304.050 595.050 ;
        RECT 305.250 593.850 307.050 594.750 ;
        RECT 301.950 590.850 304.050 591.750 ;
        RECT 313.950 568.950 316.050 571.050 ;
        RECT 314.400 559.050 315.450 568.950 ;
        RECT 313.950 556.950 316.050 559.050 ;
        RECT 259.950 553.950 262.050 556.050 ;
        RECT 292.950 554.850 295.050 555.750 ;
        RECT 313.950 554.850 316.050 555.750 ;
        RECT 277.950 547.950 280.050 550.050 ;
        RECT 256.950 544.950 259.050 547.050 ;
        RECT 226.950 528.450 229.050 529.050 ;
        RECT 226.950 527.400 231.450 528.450 ;
        RECT 226.950 526.950 229.050 527.400 ;
        RECT 226.950 524.850 229.050 525.750 ;
        RECT 230.400 523.050 231.450 527.400 ;
        RECT 232.950 526.950 235.050 529.050 ;
        RECT 257.400 526.050 258.450 544.950 ;
        RECT 278.400 529.050 279.450 547.950 ;
        RECT 313.950 529.950 316.050 532.050 ;
        RECT 265.950 526.950 268.050 529.050 ;
        RECT 271.950 526.950 274.050 529.050 ;
        RECT 275.250 527.250 276.750 528.150 ;
        RECT 277.950 526.950 280.050 529.050 ;
        RECT 310.950 527.250 313.050 528.150 ;
        RECT 313.950 527.850 316.050 528.750 ;
        RECT 232.950 524.850 235.050 525.750 ;
        RECT 256.950 523.950 259.050 526.050 ;
        RECT 229.950 520.950 232.050 523.050 ;
        RECT 205.950 494.400 208.050 496.500 ;
        RECT 226.950 495.300 229.050 497.400 ;
        RECT 206.400 477.600 207.600 494.400 ;
        RECT 227.250 491.700 228.450 495.300 ;
        RECT 226.950 489.600 229.050 491.700 ;
        RECT 257.400 490.050 258.450 523.950 ;
        RECT 211.950 485.250 214.050 486.150 ;
        RECT 217.950 485.250 220.050 486.150 ;
        RECT 211.950 481.950 214.050 484.050 ;
        RECT 217.950 481.950 220.050 484.050 ;
        RECT 205.950 475.500 208.050 477.600 ;
        RECT 218.400 457.050 219.450 481.950 ;
        RECT 227.250 477.600 228.450 489.600 ;
        RECT 256.950 487.950 259.050 490.050 ;
        RECT 266.400 489.450 267.450 526.950 ;
        RECT 268.950 523.950 271.050 526.050 ;
        RECT 272.250 524.850 273.750 525.750 ;
        RECT 274.950 523.950 277.050 526.050 ;
        RECT 278.250 524.850 280.050 525.750 ;
        RECT 310.950 523.950 313.050 526.050 ;
        RECT 268.950 521.850 271.050 522.750 ;
        RECT 275.400 508.050 276.450 523.950 ;
        RECT 316.950 520.950 319.050 523.050 ;
        RECT 274.950 505.950 277.050 508.050 ;
        RECT 286.950 505.950 289.050 508.050 ;
        RECT 266.400 488.400 270.450 489.450 ;
        RECT 250.950 484.950 253.050 487.050 ;
        RECT 229.950 483.450 232.050 484.050 ;
        RECT 229.950 482.400 234.450 483.450 ;
        RECT 229.950 481.950 232.050 482.400 ;
        RECT 229.950 479.850 232.050 480.750 ;
        RECT 233.400 478.050 234.450 482.400 ;
        RECT 226.950 475.500 229.050 477.600 ;
        RECT 232.950 475.950 235.050 478.050 ;
        RECT 244.950 475.950 247.050 478.050 ;
        RECT 245.400 460.050 246.450 475.950 ;
        RECT 244.950 457.950 247.050 460.050 ;
        RECT 211.950 455.250 214.050 456.150 ;
        RECT 217.950 454.950 220.050 457.050 ;
        RECT 244.950 455.850 247.050 456.750 ;
        RECT 247.950 455.250 250.050 456.150 ;
        RECT 218.400 454.050 219.450 454.950 ;
        RECT 211.950 451.950 214.050 454.050 ;
        RECT 217.950 451.950 220.050 454.050 ;
        RECT 247.950 453.450 250.050 454.050 ;
        RECT 251.400 453.450 252.450 484.950 ;
        RECT 257.400 481.050 258.450 487.950 ;
        RECT 269.400 487.050 270.450 488.400 ;
        RECT 265.950 485.250 267.750 486.150 ;
        RECT 268.950 484.950 271.050 487.050 ;
        RECT 274.950 484.950 277.050 487.050 ;
        RECT 277.950 484.950 280.050 487.050 ;
        RECT 265.950 481.950 268.050 484.050 ;
        RECT 269.250 482.850 271.050 483.750 ;
        RECT 271.950 482.250 274.050 483.150 ;
        RECT 274.950 482.850 277.050 483.750 ;
        RECT 256.950 478.950 259.050 481.050 ;
        RECT 271.950 478.950 274.050 481.050 ;
        RECT 247.950 452.400 252.450 453.450 ;
        RECT 247.950 451.950 250.050 452.400 ;
        RECT 220.950 415.950 223.050 418.050 ;
        RECT 250.950 415.950 253.050 418.050 ;
        RECT 221.400 415.050 222.450 415.950 ;
        RECT 220.950 412.950 223.050 415.050 ;
        RECT 217.950 410.250 220.050 411.150 ;
        RECT 220.950 410.850 223.050 411.750 ;
        RECT 217.950 406.950 220.050 409.050 ;
        RECT 229.950 391.950 232.050 394.050 ;
        RECT 190.950 385.950 193.050 388.050 ;
        RECT 202.950 385.950 205.050 388.050 ;
        RECT 187.950 382.950 190.050 385.050 ;
        RECT 191.250 383.850 192.750 384.750 ;
        RECT 193.950 382.950 196.050 385.050 ;
        RECT 230.400 382.050 231.450 391.950 ;
        RECT 187.950 380.850 190.050 381.750 ;
        RECT 193.950 380.850 196.050 381.750 ;
        RECT 226.950 380.250 228.750 381.150 ;
        RECT 229.950 379.950 232.050 382.050 ;
        RECT 233.250 380.250 235.050 381.150 ;
        RECT 226.950 376.950 229.050 379.050 ;
        RECT 230.250 377.850 231.750 378.750 ;
        RECT 232.950 376.950 235.050 379.050 ;
        RECT 196.950 343.950 199.050 346.050 ;
        RECT 202.950 344.250 205.050 345.150 ;
        RECT 197.400 343.050 198.450 343.950 ;
        RECT 181.950 340.950 184.050 343.050 ;
        RECT 193.950 341.250 195.750 342.150 ;
        RECT 196.950 340.950 199.050 343.050 ;
        RECT 200.250 341.250 201.750 342.150 ;
        RECT 202.950 340.950 205.050 343.050 ;
        RECT 182.400 340.050 183.450 340.950 ;
        RECT 227.400 340.050 228.450 376.950 ;
        RECT 235.950 349.950 238.050 352.050 ;
        RECT 236.400 343.050 237.450 349.950 ;
        RECT 251.400 346.050 252.450 415.950 ;
        RECT 256.950 414.450 259.050 415.050 ;
        RECT 254.400 413.400 259.050 414.450 ;
        RECT 254.400 385.050 255.450 413.400 ;
        RECT 256.950 412.950 259.050 413.400 ;
        RECT 256.950 410.850 259.050 411.750 ;
        RECT 259.950 410.250 262.050 411.150 ;
        RECT 259.950 406.950 262.050 409.050 ;
        RECT 260.400 397.050 261.450 406.950 ;
        RECT 259.950 394.950 262.050 397.050 ;
        RECT 274.950 394.950 277.050 397.050 ;
        RECT 268.950 391.950 271.050 394.050 ;
        RECT 259.950 385.950 262.050 388.050 ;
        RECT 260.400 385.050 261.450 385.950 ;
        RECT 253.950 382.950 256.050 385.050 ;
        RECT 259.950 382.950 262.050 385.050 ;
        RECT 263.250 383.250 264.750 384.150 ;
        RECT 265.950 382.950 268.050 385.050 ;
        RECT 254.400 382.050 255.450 382.950 ;
        RECT 269.400 382.050 270.450 391.950 ;
        RECT 253.950 379.950 256.050 382.050 ;
        RECT 259.950 380.850 261.750 381.750 ;
        RECT 262.950 379.950 265.050 382.050 ;
        RECT 266.250 380.850 267.750 381.750 ;
        RECT 268.950 379.950 271.050 382.050 ;
        RECT 254.400 379.050 255.450 379.950 ;
        RECT 253.950 376.950 256.050 379.050 ;
        RECT 268.950 377.850 271.050 378.750 ;
        RECT 238.950 344.250 241.050 345.150 ;
        RECT 250.950 343.950 253.050 346.050 ;
        RECT 235.950 342.450 238.050 343.050 ;
        RECT 238.950 342.450 241.050 343.050 ;
        RECT 235.950 341.400 241.050 342.450 ;
        RECT 235.950 340.950 238.050 341.400 ;
        RECT 238.950 340.950 241.050 341.400 ;
        RECT 242.250 341.250 243.750 342.150 ;
        RECT 244.950 340.950 247.050 343.050 ;
        RECT 248.250 341.250 250.050 342.150 ;
        RECT 172.950 337.950 175.050 340.050 ;
        RECT 181.950 337.950 184.050 340.050 ;
        RECT 193.950 337.950 196.050 340.050 ;
        RECT 197.250 338.850 198.750 339.750 ;
        RECT 199.950 337.950 202.050 340.050 ;
        RECT 226.950 337.950 229.050 340.050 ;
        RECT 241.950 337.950 244.050 340.050 ;
        RECT 245.250 338.850 246.750 339.750 ;
        RECT 247.950 339.450 250.050 340.050 ;
        RECT 251.400 339.450 252.450 343.950 ;
        RECT 259.950 340.950 262.050 343.050 ;
        RECT 247.950 338.400 252.450 339.450 ;
        RECT 247.950 337.950 250.050 338.400 ;
        RECT 182.400 310.050 183.450 337.950 ;
        RECT 196.950 331.950 199.050 334.050 ;
        RECT 226.950 331.950 229.050 334.050 ;
        RECT 184.950 316.950 187.050 319.050 ;
        RECT 185.400 313.050 186.450 316.950 ;
        RECT 190.950 313.950 193.050 316.050 ;
        RECT 184.950 310.950 187.050 313.050 ;
        RECT 188.250 311.250 190.050 312.150 ;
        RECT 190.950 311.850 193.050 312.750 ;
        RECT 193.950 311.250 196.050 312.150 ;
        RECT 181.950 307.950 184.050 310.050 ;
        RECT 184.950 308.850 186.750 309.750 ;
        RECT 187.950 307.950 190.050 310.050 ;
        RECT 193.950 307.950 196.050 310.050 ;
        RECT 188.400 307.050 189.450 307.950 ;
        RECT 187.950 304.950 190.050 307.050 ;
        RECT 181.950 271.950 184.050 274.050 ;
        RECT 187.950 271.950 190.050 274.050 ;
        RECT 193.950 272.250 196.050 273.150 ;
        RECT 182.400 247.050 183.450 271.950 ;
        RECT 188.400 271.050 189.450 271.950 ;
        RECT 184.950 269.250 186.750 270.150 ;
        RECT 187.950 268.950 190.050 271.050 ;
        RECT 193.950 270.450 196.050 271.050 ;
        RECT 197.400 270.450 198.450 331.950 ;
        RECT 202.950 313.950 205.050 316.050 ;
        RECT 199.950 310.950 202.050 313.050 ;
        RECT 200.400 307.050 201.450 310.950 ;
        RECT 203.400 310.050 204.450 313.950 ;
        RECT 227.400 310.050 228.450 331.950 ;
        RECT 247.950 313.950 250.050 316.050 ;
        RECT 229.950 310.950 232.050 313.050 ;
        RECT 235.950 312.450 238.050 313.050 ;
        RECT 233.250 311.250 234.750 312.150 ;
        RECT 235.950 311.400 240.450 312.450 ;
        RECT 235.950 310.950 238.050 311.400 ;
        RECT 202.950 307.950 205.050 310.050 ;
        RECT 226.950 307.950 229.050 310.050 ;
        RECT 230.250 308.850 231.750 309.750 ;
        RECT 232.950 307.950 235.050 310.050 ;
        RECT 236.250 308.850 238.050 309.750 ;
        RECT 199.950 304.950 202.050 307.050 ;
        RECT 226.950 305.850 229.050 306.750 ;
        RECT 239.400 304.050 240.450 311.400 ;
        RECT 238.950 301.950 241.050 304.050 ;
        RECT 205.950 278.400 208.050 280.500 ;
        RECT 226.950 279.300 229.050 281.400 ;
        RECT 191.250 269.250 192.750 270.150 ;
        RECT 193.950 269.400 198.450 270.450 ;
        RECT 193.950 268.950 196.050 269.400 ;
        RECT 184.950 265.950 187.050 268.050 ;
        RECT 188.250 266.850 189.750 267.750 ;
        RECT 190.950 265.950 193.050 268.050 ;
        RECT 184.950 259.950 187.050 262.050 ;
        RECT 181.950 244.950 184.050 247.050 ;
        RECT 185.400 241.050 186.450 259.950 ;
        RECT 191.400 249.450 192.450 265.950 ;
        RECT 206.400 261.600 207.600 278.400 ;
        RECT 214.950 274.950 217.050 277.050 ;
        RECT 227.250 275.700 228.450 279.300 ;
        RECT 211.950 269.250 214.050 270.150 ;
        RECT 211.950 265.950 214.050 268.050 ;
        RECT 215.400 267.450 216.450 274.950 ;
        RECT 226.950 273.600 229.050 275.700 ;
        RECT 217.950 269.250 220.050 270.150 ;
        RECT 217.950 267.450 220.050 268.050 ;
        RECT 215.400 266.400 220.050 267.450 ;
        RECT 217.950 265.950 220.050 266.400 ;
        RECT 212.400 262.050 213.450 265.950 ;
        RECT 205.950 259.500 208.050 261.600 ;
        RECT 211.950 259.950 214.050 262.050 ;
        RECT 227.250 261.600 228.450 273.600 ;
        RECT 248.400 268.050 249.450 313.950 ;
        RECT 256.950 307.950 259.050 310.050 ;
        RECT 260.400 309.450 261.450 340.950 ;
        RECT 275.400 339.450 276.450 394.950 ;
        RECT 278.400 382.050 279.450 484.950 ;
        RECT 287.400 481.050 288.450 505.950 ;
        RECT 292.950 490.950 295.050 493.050 ;
        RECT 310.950 490.950 313.050 493.050 ;
        RECT 286.950 478.950 289.050 481.050 ;
        RECT 287.400 457.050 288.450 478.950 ;
        RECT 280.950 456.450 283.050 457.050 ;
        RECT 280.950 455.400 285.450 456.450 ;
        RECT 280.950 454.950 283.050 455.400 ;
        RECT 280.950 452.850 283.050 453.750 ;
        RECT 277.950 379.950 280.050 382.050 ;
        RECT 284.400 346.050 285.450 455.400 ;
        RECT 286.950 454.950 289.050 457.050 ;
        RECT 286.950 452.850 289.050 453.750 ;
        RECT 293.400 418.050 294.450 490.950 ;
        RECT 311.400 490.050 312.450 490.950 ;
        RECT 304.950 487.950 307.050 490.050 ;
        RECT 308.250 488.250 309.750 489.150 ;
        RECT 310.950 487.950 313.050 490.050 ;
        RECT 304.950 485.850 306.750 486.750 ;
        RECT 307.950 484.950 310.050 487.050 ;
        RECT 311.250 485.850 313.050 486.750 ;
        RECT 298.950 461.400 301.050 463.500 ;
        RECT 299.400 444.600 300.600 461.400 ;
        RECT 308.400 459.450 309.450 484.950 ;
        RECT 305.400 458.400 309.450 459.450 ;
        RECT 317.400 483.450 318.450 520.950 ;
        RECT 322.950 495.300 325.050 497.400 ;
        RECT 323.550 491.700 324.750 495.300 ;
        RECT 338.400 493.050 339.450 595.950 ;
        RECT 346.950 561.450 349.050 562.050 ;
        RECT 344.400 560.400 349.050 561.450 ;
        RECT 344.400 529.050 345.450 560.400 ;
        RECT 346.950 559.950 349.050 560.400 ;
        RECT 350.250 560.250 351.750 561.150 ;
        RECT 346.950 557.850 348.750 558.750 ;
        RECT 349.950 556.950 352.050 559.050 ;
        RECT 353.250 557.850 355.050 558.750 ;
        RECT 346.950 544.950 349.050 547.050 ;
        RECT 347.400 532.050 348.450 544.950 ;
        RECT 371.400 532.050 372.450 673.950 ;
        RECT 388.950 670.950 391.050 673.050 ;
        RECT 379.950 668.250 381.750 669.150 ;
        RECT 382.950 667.950 385.050 670.050 ;
        RECT 386.250 668.250 388.050 669.150 ;
        RECT 379.950 664.950 382.050 667.050 ;
        RECT 383.250 665.850 384.750 666.750 ;
        RECT 385.950 666.450 388.050 667.050 ;
        RECT 389.400 666.450 390.450 670.950 ;
        RECT 392.400 670.050 393.450 674.400 ;
        RECT 419.400 673.050 420.450 697.950 ;
        RECT 442.950 676.950 445.050 679.050 ;
        RECT 427.950 673.950 430.050 676.050 ;
        RECT 428.400 673.050 429.450 673.950 ;
        RECT 418.950 670.950 421.050 673.050 ;
        RECT 421.950 670.950 424.050 673.050 ;
        RECT 425.250 671.250 426.750 672.150 ;
        RECT 427.950 670.950 430.050 673.050 ;
        RECT 391.950 667.950 394.050 670.050 ;
        RECT 418.950 669.450 421.050 670.050 ;
        RECT 416.400 668.400 421.050 669.450 ;
        RECT 422.250 668.850 423.750 669.750 ;
        RECT 385.950 665.400 390.450 666.450 ;
        RECT 385.950 664.950 388.050 665.400 ;
        RECT 380.400 652.050 381.450 664.950 ;
        RECT 388.950 652.950 391.050 655.050 ;
        RECT 379.950 649.950 382.050 652.050 ;
        RECT 379.950 629.250 382.050 630.150 ;
        RECT 385.950 629.250 388.050 630.150 ;
        RECT 379.950 627.450 382.050 628.050 ;
        RECT 377.400 626.400 382.050 627.450 ;
        RECT 385.950 627.450 388.050 628.050 ;
        RECT 389.400 627.450 390.450 652.950 ;
        RECT 416.400 631.050 417.450 668.400 ;
        RECT 418.950 667.950 421.050 668.400 ;
        RECT 424.950 667.950 427.050 670.050 ;
        RECT 428.250 668.850 430.050 669.750 ;
        RECT 418.950 665.850 421.050 666.750 ;
        RECT 418.950 658.950 421.050 661.050 ;
        RECT 419.400 634.050 420.450 658.950 ;
        RECT 418.950 631.950 421.050 634.050 ;
        RECT 443.400 631.050 444.450 676.950 ;
        RECT 460.950 671.250 463.050 672.150 ;
        RECT 460.950 667.950 463.050 670.050 ;
        RECT 461.400 655.050 462.450 667.950 ;
        RECT 464.400 667.050 465.450 701.400 ;
        RECT 466.950 700.950 469.050 701.400 ;
        RECT 472.950 701.250 475.050 702.150 ;
        RECT 466.950 698.850 469.050 699.750 ;
        RECT 476.250 698.250 478.050 699.150 ;
        RECT 500.400 697.050 501.450 704.400 ;
        RECT 502.950 703.950 505.050 704.400 ;
        RECT 506.250 704.250 507.750 705.150 ;
        RECT 541.950 704.250 544.050 705.150 ;
        RECT 610.950 703.950 613.050 706.050 ;
        RECT 616.950 703.950 619.050 706.050 ;
        RECT 691.950 705.450 694.050 706.050 ;
        RECT 620.250 704.250 621.750 705.150 ;
        RECT 689.400 704.400 694.050 705.450 ;
        RECT 502.950 701.850 504.750 702.750 ;
        RECT 505.950 700.950 508.050 703.050 ;
        RECT 509.250 701.850 511.050 702.750 ;
        RECT 535.950 700.950 538.050 703.050 ;
        RECT 541.950 700.950 544.050 703.050 ;
        RECT 545.250 701.250 546.750 702.150 ;
        RECT 547.950 700.950 550.050 703.050 ;
        RECT 551.250 701.250 553.050 702.150 ;
        RECT 580.950 701.250 583.050 702.150 ;
        RECT 586.950 701.250 589.050 702.150 ;
        RECT 475.950 694.950 478.050 697.050 ;
        RECT 499.950 694.950 502.050 697.050 ;
        RECT 532.950 694.950 535.050 697.050 ;
        RECT 469.950 679.950 472.050 682.050 ;
        RECT 505.950 679.950 508.050 682.050 ;
        RECT 470.400 676.050 471.450 679.950 ;
        RECT 469.950 673.950 472.050 676.050 ;
        RECT 475.950 673.950 478.050 676.050 ;
        RECT 502.950 673.950 505.050 676.050 ;
        RECT 466.950 670.950 469.050 673.050 ;
        RECT 470.250 671.850 472.050 672.750 ;
        RECT 466.950 668.850 469.050 669.750 ;
        RECT 463.950 664.950 466.050 667.050 ;
        RECT 460.950 652.950 463.050 655.050 ;
        RECT 415.950 628.950 418.050 631.050 ;
        RECT 418.950 629.250 420.750 630.150 ;
        RECT 421.950 628.950 424.050 631.050 ;
        RECT 427.950 630.450 430.050 631.050 ;
        RECT 427.950 629.400 432.450 630.450 ;
        RECT 427.950 628.950 430.050 629.400 ;
        RECT 377.400 604.050 378.450 626.400 ;
        RECT 379.950 625.950 382.050 626.400 ;
        RECT 383.250 626.250 384.750 627.150 ;
        RECT 385.950 626.400 390.450 627.450 ;
        RECT 416.400 627.450 417.450 628.950 ;
        RECT 418.950 627.450 421.050 628.050 ;
        RECT 416.400 626.400 421.050 627.450 ;
        RECT 422.250 626.850 424.050 627.750 ;
        RECT 385.950 625.950 388.050 626.400 ;
        RECT 418.950 625.950 421.050 626.400 ;
        RECT 424.950 626.250 427.050 627.150 ;
        RECT 427.950 626.850 430.050 627.750 ;
        RECT 431.400 625.050 432.450 629.400 ;
        RECT 442.950 628.950 445.050 631.050 ;
        RECT 460.950 629.250 463.050 630.150 ;
        RECT 466.950 629.250 469.050 630.150 ;
        RECT 472.950 628.950 475.050 631.050 ;
        RECT 460.950 625.950 463.050 628.050 ;
        RECT 464.250 626.250 465.750 627.150 ;
        RECT 466.950 625.950 469.050 628.050 ;
        RECT 382.950 622.950 385.050 625.050 ;
        RECT 424.950 622.950 427.050 625.050 ;
        RECT 427.950 622.950 430.050 625.050 ;
        RECT 430.950 622.950 433.050 625.050 ;
        RECT 463.950 622.950 466.050 625.050 ;
        RECT 376.950 601.950 379.050 604.050 ;
        RECT 377.400 598.050 378.450 601.950 ;
        RECT 383.400 601.050 384.450 622.950 ;
        RECT 425.400 622.050 426.450 622.950 ;
        RECT 415.950 619.950 418.050 622.050 ;
        RECT 424.950 619.950 427.050 622.050 ;
        RECT 382.950 598.950 385.050 601.050 ;
        RECT 412.950 598.950 415.050 601.050 ;
        RECT 373.950 596.250 375.750 597.150 ;
        RECT 376.950 595.950 379.050 598.050 ;
        RECT 380.250 596.250 382.050 597.150 ;
        RECT 412.950 596.850 415.050 597.750 ;
        RECT 373.950 592.950 376.050 595.050 ;
        RECT 377.250 593.850 378.750 594.750 ;
        RECT 379.950 592.950 382.050 595.050 ;
        RECT 416.400 594.450 417.450 619.950 ;
        RECT 421.950 600.450 424.050 601.050 ;
        RECT 421.950 599.400 426.450 600.450 ;
        RECT 421.950 598.950 424.050 599.400 ;
        RECT 418.950 596.250 421.050 597.150 ;
        RECT 421.950 596.850 424.050 597.750 ;
        RECT 418.950 594.450 421.050 595.050 ;
        RECT 416.400 593.400 421.050 594.450 ;
        RECT 418.950 592.950 421.050 593.400 ;
        RECT 374.400 559.050 375.450 592.950 ;
        RECT 376.950 586.950 379.050 589.050 ;
        RECT 373.950 556.950 376.050 559.050 ;
        RECT 373.950 532.950 376.050 535.050 ;
        RECT 346.950 529.950 349.050 532.050 ;
        RECT 370.950 529.950 373.050 532.050 ;
        RECT 343.950 526.950 346.050 529.050 ;
        RECT 347.250 527.850 348.750 528.750 ;
        RECT 374.400 526.050 375.450 532.950 ;
        RECT 343.950 524.850 346.050 525.750 ;
        RECT 349.950 524.850 352.050 525.750 ;
        RECT 373.950 523.950 376.050 526.050 ;
        RECT 343.950 494.400 346.050 496.500 ;
        RECT 322.950 489.600 325.050 491.700 ;
        RECT 337.950 490.950 340.050 493.050 ;
        RECT 319.950 483.450 322.050 484.050 ;
        RECT 317.400 482.400 322.050 483.450 ;
        RECT 305.400 457.050 306.450 458.400 ;
        RECT 304.950 454.950 307.050 457.050 ;
        RECT 310.950 454.950 313.050 457.050 ;
        RECT 313.950 454.950 316.050 457.050 ;
        RECT 304.950 452.850 307.050 453.750 ;
        RECT 310.950 452.850 313.050 453.750 ;
        RECT 298.950 442.500 301.050 444.600 ;
        RECT 307.950 423.300 310.050 425.400 ;
        RECT 308.550 419.700 309.750 423.300 ;
        RECT 292.950 415.950 295.050 418.050 ;
        RECT 296.250 416.250 297.750 417.150 ;
        RECT 298.950 415.950 301.050 418.050 ;
        RECT 307.950 417.600 310.050 419.700 ;
        RECT 292.950 413.850 294.750 414.750 ;
        RECT 295.950 412.950 298.050 415.050 ;
        RECT 299.250 413.850 301.050 414.750 ;
        RECT 296.400 352.050 297.450 412.950 ;
        RECT 304.950 411.450 307.050 412.050 ;
        RECT 302.400 410.400 307.050 411.450 ;
        RECT 302.400 397.050 303.450 410.400 ;
        RECT 304.950 409.950 307.050 410.400 ;
        RECT 304.950 407.850 307.050 408.750 ;
        RECT 308.550 405.600 309.750 417.600 ;
        RECT 314.400 411.450 315.450 454.950 ;
        RECT 317.400 438.450 318.450 482.400 ;
        RECT 319.950 481.950 322.050 482.400 ;
        RECT 319.950 479.850 322.050 480.750 ;
        RECT 323.550 477.600 324.750 489.600 ;
        RECT 331.950 485.250 334.050 486.150 ;
        RECT 337.950 485.250 340.050 486.150 ;
        RECT 331.950 481.950 334.050 484.050 ;
        RECT 337.950 481.950 340.050 484.050 ;
        RECT 322.950 475.500 325.050 477.600 ;
        RECT 319.950 461.400 322.050 463.500 ;
        RECT 332.400 463.050 333.450 481.950 ;
        RECT 338.400 481.050 339.450 481.950 ;
        RECT 337.950 478.950 340.050 481.050 ;
        RECT 344.400 477.600 345.600 494.400 ;
        RECT 377.400 483.450 378.450 586.950 ;
        RECT 380.400 535.050 381.450 592.950 ;
        RECT 415.950 589.950 418.050 592.050 ;
        RECT 412.950 559.950 415.050 562.050 ;
        RECT 382.950 557.250 385.050 558.150 ;
        RECT 388.950 557.250 391.050 558.150 ;
        RECT 382.950 553.950 385.050 556.050 ;
        RECT 386.250 554.250 387.750 555.150 ;
        RECT 388.950 553.950 391.050 556.050 ;
        RECT 383.400 547.050 384.450 553.950 ;
        RECT 385.950 550.950 388.050 553.050 ;
        RECT 389.400 547.050 390.450 553.950 ;
        RECT 413.400 553.050 414.450 559.950 ;
        RECT 412.950 550.950 415.050 553.050 ;
        RECT 382.950 544.950 385.050 547.050 ;
        RECT 388.950 544.950 391.050 547.050 ;
        RECT 391.950 544.950 394.050 547.050 ;
        RECT 379.950 532.950 382.050 535.050 ;
        RECT 382.950 529.950 385.050 532.050 ;
        RECT 379.950 527.250 382.050 528.150 ;
        RECT 382.950 527.850 385.050 528.750 ;
        RECT 385.950 527.250 387.750 528.150 ;
        RECT 388.950 526.950 391.050 529.050 ;
        RECT 392.400 526.050 393.450 544.950 ;
        RECT 379.950 523.950 382.050 526.050 ;
        RECT 385.950 523.950 388.050 526.050 ;
        RECT 389.250 524.850 391.050 525.750 ;
        RECT 391.950 523.950 394.050 526.050 ;
        RECT 379.950 485.250 382.050 486.150 ;
        RECT 385.950 485.250 388.050 486.150 ;
        RECT 379.950 483.450 382.050 484.050 ;
        RECT 377.400 482.400 382.050 483.450 ;
        RECT 343.950 475.500 346.050 477.600 ;
        RECT 346.950 472.950 349.050 475.050 ;
        RECT 320.250 449.400 321.450 461.400 ;
        RECT 331.950 460.950 334.050 463.050 ;
        RECT 322.950 458.250 325.050 459.150 ;
        RECT 325.950 457.950 328.050 460.050 ;
        RECT 322.950 456.450 325.050 457.050 ;
        RECT 326.400 456.450 327.450 457.950 ;
        RECT 332.400 457.050 333.450 460.950 ;
        RECT 322.950 455.400 327.450 456.450 ;
        RECT 322.950 454.950 325.050 455.400 ;
        RECT 331.950 454.950 334.050 457.050 ;
        RECT 319.950 447.300 322.050 449.400 ;
        RECT 320.250 443.700 321.450 447.300 ;
        RECT 319.950 441.600 322.050 443.700 ;
        RECT 317.400 437.400 321.450 438.450 ;
        RECT 316.950 413.250 319.050 414.150 ;
        RECT 316.950 411.450 319.050 412.050 ;
        RECT 314.400 410.400 319.050 411.450 ;
        RECT 316.950 409.950 319.050 410.400 ;
        RECT 320.400 408.450 321.450 437.400 ;
        RECT 328.950 422.400 331.050 424.500 ;
        RECT 343.950 422.400 346.050 424.500 ;
        RECT 322.950 413.250 325.050 414.150 ;
        RECT 325.950 412.950 328.050 415.050 ;
        RECT 322.950 409.950 325.050 412.050 ;
        RECT 317.400 407.400 321.450 408.450 ;
        RECT 317.400 406.050 318.450 407.400 ;
        RECT 307.950 403.500 310.050 405.600 ;
        RECT 316.950 403.950 319.050 406.050 ;
        RECT 301.950 394.950 304.050 397.050 ;
        RECT 304.950 394.950 307.050 397.050 ;
        RECT 305.400 388.050 306.450 394.950 ;
        RECT 304.950 385.950 307.050 388.050 ;
        RECT 298.950 382.950 301.050 385.050 ;
        RECT 301.950 383.250 304.050 384.150 ;
        RECT 304.950 383.850 307.050 384.750 ;
        RECT 307.950 383.250 309.750 384.150 ;
        RECT 310.950 382.950 313.050 385.050 ;
        RECT 299.400 379.050 300.450 382.950 ;
        RECT 301.950 379.950 304.050 382.050 ;
        RECT 304.950 379.950 307.050 382.050 ;
        RECT 307.950 379.950 310.050 382.050 ;
        RECT 311.250 380.850 313.050 381.750 ;
        RECT 298.950 376.950 301.050 379.050 ;
        RECT 295.950 349.950 298.050 352.050 ;
        RECT 283.950 343.950 286.050 346.050 ;
        RECT 286.950 344.250 289.050 345.150 ;
        RECT 298.950 343.950 301.050 346.050 ;
        RECT 277.950 341.250 279.750 342.150 ;
        RECT 280.950 340.950 283.050 343.050 ;
        RECT 284.250 341.250 285.750 342.150 ;
        RECT 286.950 340.950 289.050 343.050 ;
        RECT 277.950 339.450 280.050 340.050 ;
        RECT 275.400 338.400 280.050 339.450 ;
        RECT 281.250 338.850 282.750 339.750 ;
        RECT 277.950 337.950 280.050 338.400 ;
        RECT 283.950 337.950 286.050 340.050 ;
        RECT 299.400 319.050 300.450 343.950 ;
        RECT 305.400 343.050 306.450 379.950 ;
        RECT 304.950 340.950 307.050 343.050 ;
        RECT 308.400 328.050 309.450 379.950 ;
        RECT 307.950 325.950 310.050 328.050 ;
        RECT 298.950 316.950 301.050 319.050 ;
        RECT 262.950 313.950 265.050 316.050 ;
        RECT 299.400 313.050 300.450 316.950 ;
        RECT 262.950 311.850 265.050 312.750 ;
        RECT 265.950 311.250 268.050 312.150 ;
        RECT 283.950 310.950 286.050 313.050 ;
        RECT 298.950 310.950 301.050 313.050 ;
        RECT 304.950 310.950 307.050 313.050 ;
        RECT 310.950 310.950 313.050 313.050 ;
        RECT 265.950 309.450 268.050 310.050 ;
        RECT 260.400 308.400 268.050 309.450 ;
        RECT 229.950 265.950 232.050 268.050 ;
        RECT 247.950 265.950 250.050 268.050 ;
        RECT 257.400 265.050 258.450 307.950 ;
        RECT 263.400 271.050 264.450 308.400 ;
        RECT 265.950 307.950 268.050 308.400 ;
        RECT 262.950 268.950 265.050 271.050 ;
        RECT 268.950 268.950 271.050 271.050 ;
        RECT 272.250 269.250 274.050 270.150 ;
        RECT 262.950 266.850 265.050 267.750 ;
        RECT 265.950 266.250 268.050 267.150 ;
        RECT 268.950 266.850 270.750 267.750 ;
        RECT 271.950 265.950 274.050 268.050 ;
        RECT 229.950 263.850 232.050 264.750 ;
        RECT 256.950 262.950 259.050 265.050 ;
        RECT 265.950 262.950 268.050 265.050 ;
        RECT 272.400 262.050 273.450 265.950 ;
        RECT 226.950 259.500 229.050 261.600 ;
        RECT 271.950 259.950 274.050 262.050 ;
        RECT 229.950 256.950 232.050 259.050 ;
        RECT 188.400 248.400 192.450 249.450 ;
        RECT 188.400 244.050 189.450 248.400 ;
        RECT 190.950 244.950 193.050 247.050 ;
        RECT 191.400 244.050 192.450 244.950 ;
        RECT 187.950 241.950 190.050 244.050 ;
        RECT 190.950 241.950 193.050 244.050 ;
        RECT 230.400 241.050 231.450 256.950 ;
        RECT 184.950 238.950 187.050 241.050 ;
        RECT 188.250 239.250 190.050 240.150 ;
        RECT 190.950 239.850 193.050 240.750 ;
        RECT 193.950 239.250 196.050 240.150 ;
        RECT 217.950 238.950 220.050 241.050 ;
        RECT 223.950 238.950 226.050 241.050 ;
        RECT 227.250 239.250 228.750 240.150 ;
        RECT 229.950 238.950 232.050 241.050 ;
        RECT 268.950 239.250 271.050 240.150 ;
        RECT 184.950 236.850 186.750 237.750 ;
        RECT 187.950 235.950 190.050 238.050 ;
        RECT 193.950 235.950 196.050 238.050 ;
        RECT 142.950 232.950 145.050 235.050 ;
        RECT 146.250 233.850 147.750 234.750 ;
        RECT 148.950 232.950 151.050 235.050 ;
        RECT 163.950 232.950 166.050 235.050 ;
        RECT 143.400 205.050 144.450 232.950 ;
        RECT 142.950 202.950 145.050 205.050 ;
        RECT 145.950 202.950 148.050 205.050 ;
        RECT 146.400 202.050 147.450 202.950 ;
        RECT 139.950 199.950 142.050 202.050 ;
        RECT 145.950 199.950 148.050 202.050 ;
        RECT 149.250 200.250 150.750 201.150 ;
        RECT 151.950 199.950 154.050 202.050 ;
        RECT 140.400 163.050 141.450 199.950 ;
        RECT 145.950 197.850 147.750 198.750 ;
        RECT 148.950 196.950 151.050 199.050 ;
        RECT 152.250 197.850 154.050 198.750 ;
        RECT 149.400 196.050 150.450 196.950 ;
        RECT 148.950 193.950 151.050 196.050 ;
        RECT 142.950 190.950 145.050 193.050 ;
        RECT 139.950 160.950 142.050 163.050 ;
        RECT 143.400 127.050 144.450 190.950 ;
        RECT 157.950 178.950 160.050 181.050 ;
        RECT 158.400 169.050 159.450 178.950 ;
        RECT 164.400 172.050 165.450 232.950 ;
        RECT 184.950 197.250 187.050 198.150 ;
        RECT 190.950 197.250 193.050 198.150 ;
        RECT 194.400 196.050 195.450 235.950 ;
        RECT 199.950 199.950 202.050 202.050 ;
        RECT 184.950 193.950 187.050 196.050 ;
        RECT 188.250 194.250 189.750 195.150 ;
        RECT 190.950 193.950 193.050 196.050 ;
        RECT 193.950 193.950 196.050 196.050 ;
        RECT 191.400 193.050 192.450 193.950 ;
        RECT 187.950 190.950 190.050 193.050 ;
        RECT 190.950 190.950 193.050 193.050 ;
        RECT 163.950 169.950 166.050 172.050 ;
        RECT 157.950 166.950 160.050 169.050 ;
        RECT 161.250 167.250 163.050 168.150 ;
        RECT 163.950 167.850 166.050 168.750 ;
        RECT 166.950 167.250 169.050 168.150 ;
        RECT 188.400 166.050 189.450 190.950 ;
        RECT 200.400 175.050 201.450 199.950 ;
        RECT 218.400 199.050 219.450 238.950 ;
        RECT 223.950 236.850 225.750 237.750 ;
        RECT 226.950 235.950 229.050 238.050 ;
        RECT 230.250 236.850 231.750 237.750 ;
        RECT 232.950 237.450 235.050 238.050 ;
        RECT 232.950 236.400 237.450 237.450 ;
        RECT 232.950 235.950 235.050 236.400 ;
        RECT 227.400 208.050 228.450 235.950 ;
        RECT 232.950 233.850 235.050 234.750 ;
        RECT 226.950 205.950 229.050 208.050 ;
        RECT 220.950 202.950 223.050 205.050 ;
        RECT 229.950 202.950 232.050 205.050 ;
        RECT 221.400 202.050 222.450 202.950 ;
        RECT 220.950 199.950 223.050 202.050 ;
        RECT 224.250 200.250 225.750 201.150 ;
        RECT 226.950 199.950 229.050 202.050 ;
        RECT 217.950 196.950 220.050 199.050 ;
        RECT 220.950 197.850 222.750 198.750 ;
        RECT 223.950 196.950 226.050 199.050 ;
        RECT 227.250 197.850 229.050 198.750 ;
        RECT 199.950 172.950 202.050 175.050 ;
        RECT 200.400 172.050 201.450 172.950 ;
        RECT 193.950 169.950 196.050 172.050 ;
        RECT 199.950 169.950 202.050 172.050 ;
        RECT 205.950 169.950 208.050 172.050 ;
        RECT 157.950 164.850 159.750 165.750 ;
        RECT 160.950 163.950 163.050 166.050 ;
        RECT 166.950 163.950 169.050 166.050 ;
        RECT 187.950 163.950 190.050 166.050 ;
        RECT 194.400 165.450 195.450 169.950 ;
        RECT 206.400 169.050 207.450 169.950 ;
        RECT 196.950 167.250 199.050 168.150 ;
        RECT 199.950 167.850 202.050 168.750 ;
        RECT 202.950 167.250 204.750 168.150 ;
        RECT 205.950 166.950 208.050 169.050 ;
        RECT 196.950 165.450 199.050 166.050 ;
        RECT 194.400 164.400 199.050 165.450 ;
        RECT 196.950 163.950 199.050 164.400 ;
        RECT 202.950 163.950 205.050 166.050 ;
        RECT 206.250 164.850 208.050 165.750 ;
        RECT 148.950 128.250 151.050 129.150 ;
        RECT 139.950 125.250 141.750 126.150 ;
        RECT 142.950 124.950 145.050 127.050 ;
        RECT 146.250 125.250 147.750 126.150 ;
        RECT 148.950 124.950 151.050 127.050 ;
        RECT 161.400 124.050 162.450 163.950 ;
        RECT 203.400 133.050 204.450 163.950 ;
        RECT 202.950 130.950 205.050 133.050 ;
        RECT 196.950 127.950 199.050 130.050 ;
        RECT 184.950 124.950 187.050 127.050 ;
        RECT 139.950 121.950 142.050 124.050 ;
        RECT 143.250 122.850 144.750 123.750 ;
        RECT 145.950 121.950 148.050 124.050 ;
        RECT 160.950 121.950 163.050 124.050 ;
        RECT 184.950 122.850 187.050 123.750 ;
        RECT 187.950 122.250 190.050 123.150 ;
        RECT 140.400 97.050 141.450 121.950 ;
        RECT 197.400 121.050 198.450 127.950 ;
        RECT 203.400 121.050 204.450 130.950 ;
        RECT 223.950 127.950 226.050 130.050 ;
        RECT 224.400 127.050 225.450 127.950 ;
        RECT 230.400 127.050 231.450 202.950 ;
        RECT 217.950 124.950 220.050 127.050 ;
        RECT 223.950 124.950 226.050 127.050 ;
        RECT 227.250 125.250 229.050 126.150 ;
        RECT 229.950 124.950 232.050 127.050 ;
        RECT 217.950 122.850 220.050 123.750 ;
        RECT 220.950 122.250 223.050 123.150 ;
        RECT 223.950 122.850 225.750 123.750 ;
        RECT 226.950 121.950 229.050 124.050 ;
        RECT 230.400 121.050 231.450 124.950 ;
        RECT 236.400 124.050 237.450 236.400 ;
        RECT 268.950 235.950 271.050 238.050 ;
        RECT 250.950 199.950 253.050 202.050 ;
        RECT 259.950 201.450 262.050 202.050 ;
        RECT 257.400 200.400 262.050 201.450 ;
        RECT 238.950 169.950 241.050 172.050 ;
        RECT 238.950 167.850 240.750 168.750 ;
        RECT 241.950 168.450 244.050 169.050 ;
        RECT 241.950 167.400 246.450 168.450 ;
        RECT 241.950 166.950 244.050 167.400 ;
        RECT 241.950 164.850 244.050 165.750 ;
        RECT 245.400 124.050 246.450 167.400 ;
        RECT 247.950 167.250 250.050 168.150 ;
        RECT 247.950 165.450 250.050 166.050 ;
        RECT 251.400 165.450 252.450 199.950 ;
        RECT 247.950 164.400 252.450 165.450 ;
        RECT 247.950 163.950 250.050 164.400 ;
        RECT 253.950 127.950 256.050 130.050 ;
        RECT 235.950 121.950 238.050 124.050 ;
        RECT 244.950 121.950 247.050 124.050 ;
        RECT 142.950 118.950 145.050 121.050 ;
        RECT 187.950 118.950 190.050 121.050 ;
        RECT 196.950 118.950 199.050 121.050 ;
        RECT 202.950 118.950 205.050 121.050 ;
        RECT 220.950 118.950 223.050 121.050 ;
        RECT 229.950 118.950 232.050 121.050 ;
        RECT 139.950 94.950 142.050 97.050 ;
        RECT 143.400 57.450 144.450 118.950 ;
        RECT 181.950 99.450 184.050 100.050 ;
        RECT 179.400 98.400 184.050 99.450 ;
        RECT 148.950 94.950 151.050 97.050 ;
        RECT 149.400 94.050 150.450 94.950 ;
        RECT 145.950 92.250 147.750 93.150 ;
        RECT 148.950 91.950 151.050 94.050 ;
        RECT 152.250 92.250 154.050 93.150 ;
        RECT 179.400 91.050 180.450 98.400 ;
        RECT 181.950 97.950 184.050 98.400 ;
        RECT 181.950 95.850 184.050 96.750 ;
        RECT 184.950 95.250 187.050 96.150 ;
        RECT 184.950 91.950 187.050 94.050 ;
        RECT 145.950 88.950 148.050 91.050 ;
        RECT 149.250 89.850 150.750 90.750 ;
        RECT 151.950 88.950 154.050 91.050 ;
        RECT 178.950 88.950 181.050 91.050 ;
        RECT 146.400 61.050 147.450 88.950 ;
        RECT 152.400 76.050 153.450 88.950 ;
        RECT 151.950 73.950 154.050 76.050 ;
        RECT 157.950 73.950 160.050 76.050 ;
        RECT 145.950 58.950 148.050 61.050 ;
        RECT 151.950 59.250 154.050 60.150 ;
        RECT 145.950 57.450 148.050 58.050 ;
        RECT 143.400 56.400 148.050 57.450 ;
        RECT 145.950 55.950 148.050 56.400 ;
        RECT 149.250 56.250 150.750 57.150 ;
        RECT 151.950 55.950 154.050 58.050 ;
        RECT 155.250 56.250 157.050 57.150 ;
        RECT 145.950 53.850 147.750 54.750 ;
        RECT 148.950 52.950 151.050 55.050 ;
        RECT 151.950 52.950 154.050 55.050 ;
        RECT 154.950 52.950 157.050 55.050 ;
        RECT 40.950 43.950 43.050 46.050 ;
        RECT 112.950 43.950 115.050 46.050 ;
        RECT 136.950 43.950 139.050 46.050 ;
        RECT 31.950 20.250 33.750 21.150 ;
        RECT 34.950 19.950 37.050 22.050 ;
        RECT 38.250 20.250 40.050 21.150 ;
        RECT 35.250 17.850 36.750 18.750 ;
        RECT 37.950 18.450 40.050 19.050 ;
        RECT 41.400 18.450 42.450 43.950 ;
        RECT 149.400 43.050 150.450 52.950 ;
        RECT 115.950 40.950 118.050 43.050 ;
        RECT 148.950 40.950 151.050 43.050 ;
        RECT 79.950 28.950 82.050 31.050 ;
        RECT 80.400 25.050 81.450 28.950 ;
        RECT 116.400 28.050 117.450 40.950 ;
        RECT 145.950 28.950 148.050 31.050 ;
        RECT 115.950 25.950 118.050 28.050 ;
        RECT 118.950 25.950 121.050 28.050 ;
        RECT 119.400 25.050 120.450 25.950 ;
        RECT 146.400 25.050 147.450 28.950 ;
        RECT 148.950 27.450 151.050 28.050 ;
        RECT 152.400 27.450 153.450 52.950 ;
        RECT 155.400 52.050 156.450 52.950 ;
        RECT 158.400 52.050 159.450 73.950 ;
        RECT 193.950 56.250 196.050 57.150 ;
        RECT 184.950 53.250 186.750 54.150 ;
        RECT 187.950 52.950 190.050 55.050 ;
        RECT 191.250 53.250 192.750 54.150 ;
        RECT 193.950 52.950 196.050 55.050 ;
        RECT 197.400 52.050 198.450 118.950 ;
        RECT 223.950 100.950 226.050 103.050 ;
        RECT 217.950 97.950 220.050 100.050 ;
        RECT 218.400 97.050 219.450 97.950 ;
        RECT 224.400 97.050 225.450 100.950 ;
        RECT 245.400 97.050 246.450 121.950 ;
        RECT 217.950 96.450 220.050 97.050 ;
        RECT 215.400 95.400 220.050 96.450 ;
        RECT 215.400 94.050 216.450 95.400 ;
        RECT 217.950 94.950 220.050 95.400 ;
        RECT 221.250 95.250 222.750 96.150 ;
        RECT 223.950 94.950 226.050 97.050 ;
        RECT 244.950 94.950 247.050 97.050 ;
        RECT 214.950 91.950 217.050 94.050 ;
        RECT 217.950 92.850 219.750 93.750 ;
        RECT 220.950 91.950 223.050 94.050 ;
        RECT 224.250 92.850 225.750 93.750 ;
        RECT 226.950 93.450 229.050 94.050 ;
        RECT 226.950 92.400 231.450 93.450 ;
        RECT 226.950 91.950 229.050 92.400 ;
        RECT 226.950 89.850 229.050 90.750 ;
        RECT 230.400 76.050 231.450 92.400 ;
        RECT 229.950 73.950 232.050 76.050 ;
        RECT 199.950 55.950 202.050 58.050 ;
        RECT 230.250 56.250 231.750 57.150 ;
        RECT 232.950 55.950 235.050 58.050 ;
        RECT 154.950 49.950 157.050 52.050 ;
        RECT 157.950 49.950 160.050 52.050 ;
        RECT 184.950 49.950 187.050 52.050 ;
        RECT 188.250 50.850 189.750 51.750 ;
        RECT 190.950 49.950 193.050 52.050 ;
        RECT 196.950 49.950 199.050 52.050 ;
        RECT 148.950 26.400 153.450 27.450 ;
        RECT 148.950 25.950 151.050 26.400 ;
        RECT 70.950 22.950 73.050 25.050 ;
        RECT 79.950 22.950 82.050 25.050 ;
        RECT 112.950 22.950 115.050 25.050 ;
        RECT 116.250 23.850 117.750 24.750 ;
        RECT 118.950 22.950 121.050 25.050 ;
        RECT 145.950 22.950 148.050 25.050 ;
        RECT 149.250 23.850 150.750 24.750 ;
        RECT 155.400 22.050 156.450 49.950 ;
        RECT 185.400 46.050 186.450 49.950 ;
        RECT 196.950 46.950 199.050 49.050 ;
        RECT 184.950 43.950 187.050 46.050 ;
        RECT 184.950 28.950 187.050 31.050 ;
        RECT 185.400 28.050 186.450 28.950 ;
        RECT 184.950 25.950 187.050 28.050 ;
        RECT 184.950 23.850 186.750 24.750 ;
        RECT 193.950 23.250 196.050 24.150 ;
        RECT 70.950 20.850 73.050 21.750 ;
        RECT 73.950 20.250 76.050 21.150 ;
        RECT 79.950 20.850 82.050 21.750 ;
        RECT 112.950 20.850 115.050 21.750 ;
        RECT 118.950 20.850 121.050 21.750 ;
        RECT 145.950 20.850 148.050 21.750 ;
        RECT 151.950 20.850 154.050 21.750 ;
        RECT 154.950 19.950 157.050 22.050 ;
        RECT 187.950 20.850 190.050 21.750 ;
        RECT 193.950 21.450 196.050 22.050 ;
        RECT 197.400 21.450 198.450 46.950 ;
        RECT 200.400 28.050 201.450 55.950 ;
        RECT 226.950 53.850 228.750 54.750 ;
        RECT 229.950 52.950 232.050 55.050 ;
        RECT 233.250 53.850 235.050 54.750 ;
        RECT 220.950 31.950 223.050 34.050 ;
        RECT 205.950 29.400 208.050 31.500 ;
        RECT 199.950 25.950 202.050 28.050 ;
        RECT 202.950 26.250 205.050 27.150 ;
        RECT 200.400 24.450 201.450 25.950 ;
        RECT 202.950 24.450 205.050 25.050 ;
        RECT 200.400 23.400 205.050 24.450 ;
        RECT 202.950 22.950 205.050 23.400 ;
        RECT 193.950 20.400 198.450 21.450 ;
        RECT 193.950 19.950 196.050 20.400 ;
        RECT 37.950 17.400 42.450 18.450 ;
        RECT 206.550 17.400 207.750 29.400 ;
        RECT 214.950 25.950 217.050 28.050 ;
        RECT 215.400 25.050 216.450 25.950 ;
        RECT 221.400 25.050 222.450 31.950 ;
        RECT 226.950 29.400 229.050 31.500 ;
        RECT 241.950 29.400 244.050 31.500 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 220.950 22.950 223.050 25.050 ;
        RECT 214.950 20.850 217.050 21.750 ;
        RECT 220.950 20.850 223.050 21.750 ;
        RECT 37.950 16.950 40.050 17.400 ;
        RECT 205.950 15.300 208.050 17.400 ;
        RECT 206.550 11.700 207.750 15.300 ;
        RECT 227.400 12.600 228.600 29.400 ;
        RECT 242.400 12.600 243.600 29.400 ;
        RECT 254.400 28.050 255.450 127.950 ;
        RECT 257.400 121.050 258.450 200.400 ;
        RECT 259.950 199.950 262.050 200.400 ;
        RECT 263.250 200.250 264.750 201.150 ;
        RECT 265.950 199.950 268.050 202.050 ;
        RECT 259.950 197.850 261.750 198.750 ;
        RECT 262.950 196.950 265.050 199.050 ;
        RECT 266.250 197.850 268.050 198.750 ;
        RECT 263.400 196.050 264.450 196.950 ;
        RECT 262.950 193.950 265.050 196.050 ;
        RECT 269.400 178.050 270.450 235.950 ;
        RECT 268.950 175.950 271.050 178.050 ;
        RECT 259.950 169.950 262.050 172.050 ;
        RECT 256.950 118.950 259.050 121.050 ;
        RECT 260.400 94.050 261.450 169.950 ;
        RECT 269.400 130.050 270.450 175.950 ;
        RECT 284.400 172.050 285.450 310.950 ;
        RECT 311.400 310.050 312.450 310.950 ;
        RECT 298.950 308.850 301.050 309.750 ;
        RECT 304.950 308.850 307.050 309.750 ;
        RECT 310.950 307.950 313.050 310.050 ;
        RECT 311.400 277.050 312.450 307.950 ;
        RECT 310.950 274.950 313.050 277.050 ;
        RECT 304.950 272.250 307.050 273.150 ;
        RECT 311.400 271.050 312.450 274.950 ;
        RECT 304.950 268.950 307.050 271.050 ;
        RECT 308.250 269.250 309.750 270.150 ;
        RECT 310.950 268.950 313.050 271.050 ;
        RECT 314.250 269.250 316.050 270.150 ;
        RECT 289.950 239.250 292.050 240.150 ;
        RECT 301.950 197.250 304.050 198.150 ;
        RECT 301.950 193.950 304.050 196.050 ;
        RECT 283.950 169.950 286.050 172.050 ;
        RECT 284.400 169.050 285.450 169.950 ;
        RECT 302.400 169.050 303.450 193.950 ;
        RECT 305.400 190.050 306.450 268.950 ;
        RECT 307.950 265.950 310.050 268.050 ;
        RECT 311.250 266.850 312.750 267.750 ;
        RECT 313.950 265.950 316.050 268.050 ;
        RECT 314.400 256.050 315.450 265.950 ;
        RECT 313.950 253.950 316.050 256.050 ;
        RECT 307.950 197.250 310.050 198.150 ;
        RECT 307.950 193.950 310.050 196.050 ;
        RECT 308.400 193.050 309.450 193.950 ;
        RECT 317.400 193.050 318.450 403.950 ;
        RECT 323.400 400.050 324.450 409.950 ;
        RECT 322.950 397.950 325.050 400.050 ;
        RECT 319.950 344.250 322.050 345.150 ;
        RECT 326.400 343.050 327.450 412.950 ;
        RECT 329.400 405.600 330.600 422.400 ;
        RECT 344.400 405.600 345.600 422.400 ;
        RECT 328.950 403.500 331.050 405.600 ;
        RECT 343.950 403.500 346.050 405.600 ;
        RECT 343.950 397.950 346.050 400.050 ;
        RECT 344.400 388.050 345.450 397.950 ;
        RECT 347.400 391.050 348.450 472.950 ;
        RECT 370.950 461.400 373.050 463.500 ;
        RECT 355.950 457.950 358.050 460.050 ;
        RECT 367.950 458.250 370.050 459.150 ;
        RECT 355.950 455.850 358.050 456.750 ;
        RECT 358.950 455.250 361.050 456.150 ;
        RECT 367.950 454.950 370.050 457.050 ;
        RECT 358.950 451.950 361.050 454.050 ;
        RECT 364.950 423.300 367.050 425.400 ;
        RECT 365.250 419.700 366.450 423.300 ;
        RECT 364.950 417.600 367.050 419.700 ;
        RECT 368.400 418.050 369.450 454.950 ;
        RECT 371.550 449.400 372.750 461.400 ;
        RECT 377.400 454.050 378.450 482.400 ;
        RECT 379.950 481.950 382.050 482.400 ;
        RECT 383.250 482.250 384.750 483.150 ;
        RECT 385.950 481.950 388.050 484.050 ;
        RECT 382.950 478.950 385.050 481.050 ;
        RECT 386.400 475.050 387.450 481.950 ;
        RECT 385.950 472.950 388.050 475.050 ;
        RECT 379.950 460.950 382.050 463.050 ;
        RECT 385.950 460.950 388.050 463.050 ;
        RECT 391.950 461.400 394.050 463.500 ;
        RECT 380.400 457.050 381.450 460.950 ;
        RECT 386.400 457.050 387.450 460.950 ;
        RECT 379.950 454.950 382.050 457.050 ;
        RECT 385.950 454.950 388.050 457.050 ;
        RECT 376.950 451.950 379.050 454.050 ;
        RECT 379.950 452.850 382.050 453.750 ;
        RECT 385.950 452.850 388.050 453.750 ;
        RECT 370.950 447.300 373.050 449.400 ;
        RECT 371.550 443.700 372.750 447.300 ;
        RECT 392.400 444.600 393.600 461.400 ;
        RECT 370.950 441.600 373.050 443.700 ;
        RECT 391.950 442.500 394.050 444.600 ;
        RECT 349.950 413.250 352.050 414.150 ;
        RECT 355.950 413.250 358.050 414.150 ;
        RECT 349.950 409.950 352.050 412.050 ;
        RECT 355.950 409.950 358.050 412.050 ;
        RECT 350.400 409.050 351.450 409.950 ;
        RECT 349.950 406.950 352.050 409.050 ;
        RECT 365.250 405.600 366.450 417.600 ;
        RECT 367.950 415.950 370.050 418.050 ;
        RECT 403.950 414.450 406.050 415.050 ;
        RECT 406.950 414.450 409.050 415.050 ;
        RECT 403.950 413.400 409.050 414.450 ;
        RECT 403.950 412.950 406.050 413.400 ;
        RECT 406.950 412.950 409.050 413.400 ;
        RECT 367.950 411.450 370.050 412.050 ;
        RECT 367.950 410.400 372.450 411.450 ;
        RECT 367.950 409.950 370.050 410.400 ;
        RECT 371.400 409.050 372.450 410.400 ;
        RECT 400.950 410.250 403.050 411.150 ;
        RECT 403.950 410.850 406.050 411.750 ;
        RECT 367.950 407.850 370.050 408.750 ;
        RECT 370.950 406.950 373.050 409.050 ;
        RECT 400.950 406.950 403.050 409.050 ;
        RECT 364.950 403.500 367.050 405.600 ;
        RECT 346.950 388.950 349.050 391.050 ;
        RECT 343.950 385.950 346.050 388.050 ;
        RECT 347.400 385.050 348.450 388.950 ;
        RECT 340.950 382.950 343.050 385.050 ;
        RECT 344.250 383.850 345.750 384.750 ;
        RECT 346.950 382.950 349.050 385.050 ;
        RECT 349.950 382.950 352.050 385.050 ;
        RECT 382.950 382.950 385.050 385.050 ;
        RECT 400.950 382.950 403.050 385.050 ;
        RECT 340.950 380.850 343.050 381.750 ;
        RECT 346.950 380.850 349.050 381.750 ;
        RECT 350.400 376.050 351.450 382.950 ;
        RECT 376.950 380.850 379.050 381.750 ;
        RECT 382.950 380.850 385.050 381.750 ;
        RECT 349.950 373.950 352.050 376.050 ;
        RECT 337.950 351.300 340.050 353.400 ;
        RECT 338.550 347.700 339.750 351.300 ;
        RECT 337.950 345.600 340.050 347.700 ;
        RECT 319.950 340.950 322.050 343.050 ;
        RECT 323.250 341.250 324.750 342.150 ;
        RECT 325.950 340.950 328.050 343.050 ;
        RECT 329.250 341.250 331.050 342.150 ;
        RECT 320.400 340.050 321.450 340.950 ;
        RECT 319.950 337.950 322.050 340.050 ;
        RECT 322.950 337.950 325.050 340.050 ;
        RECT 326.250 338.850 327.750 339.750 ;
        RECT 328.950 337.950 331.050 340.050 ;
        RECT 334.950 339.450 337.050 340.050 ;
        RECT 332.400 338.400 337.050 339.450 ;
        RECT 323.400 307.050 324.450 337.950 ;
        RECT 329.400 310.050 330.450 337.950 ;
        RECT 332.400 328.050 333.450 338.400 ;
        RECT 334.950 337.950 337.050 338.400 ;
        RECT 334.950 335.850 337.050 336.750 ;
        RECT 338.550 333.600 339.750 345.600 ;
        RECT 346.950 341.250 349.050 342.150 ;
        RECT 350.400 340.050 351.450 373.950 ;
        RECT 358.950 350.400 361.050 352.500 ;
        RECT 352.950 341.250 355.050 342.150 ;
        RECT 346.950 339.450 349.050 340.050 ;
        RECT 344.400 338.400 349.050 339.450 ;
        RECT 337.950 331.500 340.050 333.600 ;
        RECT 331.950 325.950 334.050 328.050 ;
        RECT 337.950 325.950 340.050 328.050 ;
        RECT 338.400 316.050 339.450 325.950 ;
        RECT 337.950 313.950 340.050 316.050 ;
        RECT 337.950 311.850 340.050 312.750 ;
        RECT 340.950 311.250 343.050 312.150 ;
        RECT 328.950 307.950 331.050 310.050 ;
        RECT 340.950 307.950 343.050 310.050 ;
        RECT 322.950 304.950 325.050 307.050 ;
        RECT 325.950 239.250 328.050 240.150 ;
        RECT 344.400 238.050 345.450 338.400 ;
        RECT 346.950 337.950 349.050 338.400 ;
        RECT 349.950 337.950 352.050 340.050 ;
        RECT 352.950 337.950 355.050 340.050 ;
        RECT 359.400 333.600 360.600 350.400 ;
        RECT 401.400 346.050 402.450 382.950 ;
        RECT 416.400 375.450 417.450 589.950 ;
        RECT 425.400 568.050 426.450 599.400 ;
        RECT 428.400 592.050 429.450 622.950 ;
        RECT 464.400 622.050 465.450 622.950 ;
        RECT 463.950 619.950 466.050 622.050 ;
        RECT 460.950 597.450 463.050 598.050 ;
        RECT 464.400 597.450 465.450 619.950 ;
        RECT 467.400 619.050 468.450 625.950 ;
        RECT 466.950 616.950 469.050 619.050 ;
        RECT 457.950 596.250 459.750 597.150 ;
        RECT 460.950 596.400 465.450 597.450 ;
        RECT 460.950 595.950 463.050 596.400 ;
        RECT 466.950 595.950 469.050 598.050 ;
        RECT 454.950 592.950 457.050 595.050 ;
        RECT 457.950 592.950 460.050 595.050 ;
        RECT 461.250 593.850 462.750 594.750 ;
        RECT 463.950 592.950 466.050 595.050 ;
        RECT 467.250 593.850 469.050 594.750 ;
        RECT 427.950 589.950 430.050 592.050 ;
        RECT 424.950 565.950 427.050 568.050 ;
        RECT 433.950 559.950 436.050 562.050 ;
        RECT 418.950 556.950 421.050 559.050 ;
        RECT 424.950 558.450 427.050 559.050 ;
        RECT 424.950 557.400 429.450 558.450 ;
        RECT 424.950 556.950 427.050 557.400 ;
        RECT 419.400 552.450 420.450 556.950 ;
        RECT 421.950 554.250 424.050 555.150 ;
        RECT 424.950 554.850 427.050 555.750 ;
        RECT 421.950 552.450 424.050 553.050 ;
        RECT 419.400 551.400 424.050 552.450 ;
        RECT 421.950 550.950 424.050 551.400 ;
        RECT 428.400 547.050 429.450 557.400 ;
        RECT 430.950 553.950 433.050 556.050 ;
        RECT 427.950 544.950 430.050 547.050 ;
        RECT 421.950 526.950 424.050 529.050 ;
        RECT 424.950 526.950 427.050 529.050 ;
        RECT 422.400 523.050 423.450 526.950 ;
        RECT 424.950 524.850 427.050 525.750 ;
        RECT 427.950 524.250 430.050 525.150 ;
        RECT 421.950 520.950 424.050 523.050 ;
        RECT 427.950 520.950 430.050 523.050 ;
        RECT 427.950 490.950 430.050 493.050 ;
        RECT 421.950 488.250 424.050 489.150 ;
        RECT 428.400 487.050 429.450 490.950 ;
        RECT 431.400 489.450 432.450 553.950 ;
        RECT 434.400 529.050 435.450 559.950 ;
        RECT 455.400 559.050 456.450 592.950 ;
        RECT 458.400 565.050 459.450 592.950 ;
        RECT 463.950 590.850 466.050 591.750 ;
        RECT 457.950 562.950 460.050 565.050 ;
        RECT 466.950 563.250 469.050 564.150 ;
        RECT 457.950 559.950 460.050 562.050 ;
        RECT 460.950 559.950 463.050 562.050 ;
        RECT 464.250 560.250 465.750 561.150 ;
        RECT 466.950 559.950 469.050 562.050 ;
        RECT 470.250 560.250 472.050 561.150 ;
        RECT 454.950 556.950 457.050 559.050 ;
        RECT 436.950 550.950 439.050 553.050 ;
        RECT 433.950 526.950 436.050 529.050 ;
        RECT 433.950 524.850 436.050 525.750 ;
        RECT 431.400 488.400 435.450 489.450 ;
        RECT 421.950 484.950 424.050 487.050 ;
        RECT 425.250 485.250 426.750 486.150 ;
        RECT 427.950 484.950 430.050 487.050 ;
        RECT 431.250 485.250 433.050 486.150 ;
        RECT 422.400 454.050 423.450 484.950 ;
        RECT 424.950 481.950 427.050 484.050 ;
        RECT 428.250 482.850 429.750 483.750 ;
        RECT 430.950 481.950 433.050 484.050 ;
        RECT 421.950 451.950 424.050 454.050 ;
        RECT 422.400 385.050 423.450 451.950 ;
        RECT 425.400 415.050 426.450 481.950 ;
        RECT 430.950 457.950 433.050 460.050 ;
        RECT 434.400 457.050 435.450 488.400 ;
        RECT 437.400 484.050 438.450 550.950 ;
        RECT 458.400 520.050 459.450 559.950 ;
        RECT 460.950 557.850 462.750 558.750 ;
        RECT 463.950 556.950 466.050 559.050 ;
        RECT 469.950 558.450 472.050 559.050 ;
        RECT 473.400 558.450 474.450 628.950 ;
        RECT 476.400 598.050 477.450 673.950 ;
        RECT 506.400 673.050 507.450 679.950 ;
        RECT 499.950 670.950 502.050 673.050 ;
        RECT 503.250 671.850 504.750 672.750 ;
        RECT 505.950 670.950 508.050 673.050 ;
        RECT 499.950 668.850 502.050 669.750 ;
        RECT 502.950 667.950 505.050 670.050 ;
        RECT 505.950 668.850 508.050 669.750 ;
        RECT 493.950 628.950 496.050 631.050 ;
        RECT 499.950 628.950 502.050 631.050 ;
        RECT 475.950 595.950 478.050 598.050 ;
        RECT 494.400 597.450 495.450 628.950 ;
        RECT 503.400 628.050 504.450 667.950 ;
        RECT 505.950 629.250 508.050 630.150 ;
        RECT 511.950 628.950 514.050 631.050 ;
        RECT 499.950 626.850 502.050 627.750 ;
        RECT 502.950 627.450 505.050 628.050 ;
        RECT 505.950 627.450 508.050 628.050 ;
        RECT 502.950 626.400 508.050 627.450 ;
        RECT 502.950 625.950 505.050 626.400 ;
        RECT 505.950 625.950 508.050 626.400 ;
        RECT 509.250 626.250 511.050 627.150 ;
        RECT 506.400 622.050 507.450 625.950 ;
        RECT 508.950 624.450 511.050 625.050 ;
        RECT 512.400 624.450 513.450 628.950 ;
        RECT 508.950 623.400 513.450 624.450 ;
        RECT 508.950 622.950 511.050 623.400 ;
        RECT 505.950 619.950 508.050 622.050 ;
        RECT 499.950 604.950 502.050 607.050 ;
        RECT 517.950 605.400 520.050 607.500 ;
        RECT 500.400 604.050 501.450 604.950 ;
        RECT 499.950 601.950 502.050 604.050 ;
        RECT 496.950 599.250 499.050 600.150 ;
        RECT 499.950 599.850 502.050 600.750 ;
        RECT 502.950 599.250 504.750 600.150 ;
        RECT 505.950 598.950 508.050 601.050 ;
        RECT 496.950 597.450 499.050 598.050 ;
        RECT 494.400 596.400 499.050 597.450 ;
        RECT 496.950 595.950 499.050 596.400 ;
        RECT 502.950 595.950 505.050 598.050 ;
        RECT 506.250 596.850 508.050 597.750 ;
        RECT 476.400 562.050 477.450 595.950 ;
        RECT 503.400 595.050 504.450 595.950 ;
        RECT 496.950 592.950 499.050 595.050 ;
        RECT 502.950 592.950 505.050 595.050 ;
        RECT 490.950 562.950 493.050 565.050 ;
        RECT 475.950 559.950 478.050 562.050 ;
        RECT 469.950 557.400 474.450 558.450 ;
        RECT 469.950 556.950 472.050 557.400 ;
        RECT 475.950 526.950 478.050 529.050 ;
        RECT 463.950 524.250 465.750 525.150 ;
        RECT 466.950 523.950 469.050 526.050 ;
        RECT 470.250 524.250 472.050 525.150 ;
        RECT 463.950 520.950 466.050 523.050 ;
        RECT 467.250 521.850 468.750 522.750 ;
        RECT 469.950 520.950 472.050 523.050 ;
        RECT 470.400 520.050 471.450 520.950 ;
        RECT 457.950 517.950 460.050 520.050 ;
        RECT 469.950 517.950 472.050 520.050 ;
        RECT 463.950 484.950 466.050 487.050 ;
        RECT 472.950 484.950 475.050 487.050 ;
        RECT 436.950 481.950 439.050 484.050 ;
        RECT 460.950 482.250 463.050 483.150 ;
        RECT 463.950 482.850 466.050 483.750 ;
        RECT 460.950 478.950 463.050 481.050 ;
        RECT 466.950 460.950 469.050 463.050 ;
        RECT 467.400 460.050 468.450 460.950 ;
        RECT 463.950 457.950 466.050 460.050 ;
        RECT 466.950 457.950 469.050 460.050 ;
        RECT 469.950 457.950 472.050 460.050 ;
        RECT 464.400 457.050 465.450 457.950 ;
        RECT 470.400 457.050 471.450 457.950 ;
        RECT 427.950 454.950 430.050 457.050 ;
        RECT 431.250 455.850 432.750 456.750 ;
        RECT 433.950 454.950 436.050 457.050 ;
        RECT 463.950 454.950 466.050 457.050 ;
        RECT 467.250 455.850 468.750 456.750 ;
        RECT 469.950 454.950 472.050 457.050 ;
        RECT 427.950 452.850 430.050 453.750 ;
        RECT 433.950 452.850 436.050 453.750 ;
        RECT 463.950 452.850 466.050 453.750 ;
        RECT 469.950 452.850 472.050 453.750 ;
        RECT 424.950 412.950 427.050 415.050 ;
        RECT 433.950 414.450 436.050 415.050 ;
        RECT 436.950 414.450 439.050 415.050 ;
        RECT 433.950 413.400 439.050 414.450 ;
        RECT 433.950 412.950 436.050 413.400 ;
        RECT 436.950 412.950 439.050 413.400 ;
        RECT 442.950 412.950 445.050 415.050 ;
        RECT 446.250 413.250 448.050 414.150 ;
        RECT 436.950 410.850 439.050 411.750 ;
        RECT 439.950 410.250 442.050 411.150 ;
        RECT 442.950 410.850 444.750 411.750 ;
        RECT 445.950 409.950 448.050 412.050 ;
        RECT 439.950 406.950 442.050 409.050 ;
        RECT 473.400 385.050 474.450 484.950 ;
        RECT 476.400 414.450 477.450 526.950 ;
        RECT 487.950 523.950 490.050 526.050 ;
        RECT 488.400 490.050 489.450 523.950 ;
        RECT 487.950 487.950 490.050 490.050 ;
        RECT 491.400 459.450 492.450 562.950 ;
        RECT 493.950 556.950 496.050 559.050 ;
        RECT 494.400 526.050 495.450 556.950 ;
        RECT 497.400 555.450 498.450 592.950 ;
        RECT 518.400 588.600 519.600 605.400 ;
        RECT 533.400 601.050 534.450 694.950 ;
        RECT 536.400 666.450 537.450 700.950 ;
        RECT 544.950 697.950 547.050 700.050 ;
        RECT 548.250 698.850 549.750 699.750 ;
        RECT 550.950 697.950 553.050 700.050 ;
        RECT 580.950 697.950 583.050 700.050 ;
        RECT 584.250 698.250 585.750 699.150 ;
        RECT 545.400 679.050 546.450 697.950 ;
        RECT 551.400 685.050 552.450 697.950 ;
        RECT 581.400 697.050 582.450 697.950 ;
        RECT 580.950 694.950 583.050 697.050 ;
        RECT 583.950 694.950 586.050 697.050 ;
        RECT 550.950 682.950 553.050 685.050 ;
        RECT 586.950 682.950 589.050 685.050 ;
        RECT 544.950 676.950 547.050 679.050 ;
        RECT 550.950 670.950 553.050 673.050 ;
        RECT 577.950 672.450 580.050 673.050 ;
        RECT 575.400 671.400 580.050 672.450 ;
        RECT 538.950 668.250 540.750 669.150 ;
        RECT 541.950 667.950 544.050 670.050 ;
        RECT 545.250 668.250 547.050 669.150 ;
        RECT 538.950 666.450 541.050 667.050 ;
        RECT 536.400 665.400 541.050 666.450 ;
        RECT 542.250 665.850 543.750 666.750 ;
        RECT 538.950 664.950 541.050 665.400 ;
        RECT 544.950 664.950 547.050 667.050 ;
        RECT 535.950 631.950 538.050 634.050 ;
        RECT 544.950 631.950 547.050 634.050 ;
        RECT 523.950 598.950 526.050 601.050 ;
        RECT 529.950 600.450 532.050 601.050 ;
        RECT 527.400 599.400 532.050 600.450 ;
        RECT 523.950 596.850 526.050 597.750 ;
        RECT 517.950 586.500 520.050 588.600 ;
        RECT 527.400 571.050 528.450 599.400 ;
        RECT 529.950 598.950 532.050 599.400 ;
        RECT 532.950 598.950 535.050 601.050 ;
        RECT 529.950 596.850 532.050 597.750 ;
        RECT 526.950 568.950 529.050 571.050 ;
        RECT 529.950 568.950 532.050 571.050 ;
        RECT 499.950 560.250 502.050 561.150 ;
        RECT 511.950 559.950 514.050 562.050 ;
        RECT 499.950 556.950 502.050 559.050 ;
        RECT 503.250 557.250 504.750 558.150 ;
        RECT 505.950 556.950 508.050 559.050 ;
        RECT 509.250 557.250 511.050 558.150 ;
        RECT 502.950 555.450 505.050 556.050 ;
        RECT 497.400 554.400 505.050 555.450 ;
        RECT 506.250 554.850 507.750 555.750 ;
        RECT 502.950 553.950 505.050 554.400 ;
        RECT 508.950 553.950 511.050 556.050 ;
        RECT 509.400 553.050 510.450 553.950 ;
        RECT 508.950 550.950 511.050 553.050 ;
        RECT 512.400 529.050 513.450 559.950 ;
        RECT 520.950 533.400 523.050 535.500 ;
        RECT 517.950 530.250 520.050 531.150 ;
        RECT 499.950 526.950 502.050 529.050 ;
        RECT 505.950 526.950 508.050 529.050 ;
        RECT 509.250 527.250 510.750 528.150 ;
        RECT 511.950 526.950 514.050 529.050 ;
        RECT 517.950 526.950 520.050 529.050 ;
        RECT 493.950 523.950 496.050 526.050 ;
        RECT 496.950 484.950 499.050 487.050 ;
        RECT 500.400 486.450 501.450 526.950 ;
        RECT 502.950 523.950 505.050 526.050 ;
        RECT 506.250 524.850 507.750 525.750 ;
        RECT 508.950 523.950 511.050 526.050 ;
        RECT 512.250 524.850 514.050 525.750 ;
        RECT 509.400 523.050 510.450 523.950 ;
        RECT 502.950 521.850 505.050 522.750 ;
        RECT 508.950 520.950 511.050 523.050 ;
        RECT 521.550 521.400 522.750 533.400 ;
        RECT 530.400 529.050 531.450 568.950 ;
        RECT 533.400 553.050 534.450 598.950 ;
        RECT 536.400 582.450 537.450 631.950 ;
        RECT 545.400 631.050 546.450 631.950 ;
        RECT 551.400 631.050 552.450 670.950 ;
        RECT 575.400 634.050 576.450 671.400 ;
        RECT 577.950 670.950 580.050 671.400 ;
        RECT 581.250 671.250 582.750 672.150 ;
        RECT 583.950 670.950 586.050 673.050 ;
        RECT 587.400 670.050 588.450 682.950 ;
        RECT 611.400 676.050 612.450 703.950 ;
        RECT 616.950 701.850 618.750 702.750 ;
        RECT 619.950 700.950 622.050 703.050 ;
        RECT 623.250 701.850 625.050 702.750 ;
        RECT 658.950 701.250 661.050 702.150 ;
        RECT 664.950 701.250 667.050 702.150 ;
        RECT 610.950 673.950 613.050 676.050 ;
        RECT 577.950 668.850 579.750 669.750 ;
        RECT 580.950 667.950 583.050 670.050 ;
        RECT 584.250 668.850 585.750 669.750 ;
        RECT 586.950 667.950 589.050 670.050 ;
        RECT 581.400 666.450 582.450 667.950 ;
        RECT 581.400 665.400 585.450 666.450 ;
        RECT 586.950 665.850 589.050 666.750 ;
        RECT 574.950 631.950 577.050 634.050 ;
        RECT 541.950 629.250 543.750 630.150 ;
        RECT 544.950 628.950 547.050 631.050 ;
        RECT 550.950 628.950 553.050 631.050 ;
        RECT 541.950 625.950 544.050 628.050 ;
        RECT 545.250 626.850 547.050 627.750 ;
        RECT 547.950 626.250 550.050 627.150 ;
        RECT 550.950 626.850 553.050 627.750 ;
        RECT 538.950 605.400 541.050 607.500 ;
        RECT 542.400 607.050 543.450 625.950 ;
        RECT 547.950 622.950 550.050 625.050 ;
        RECT 548.400 622.050 549.450 622.950 ;
        RECT 547.950 619.950 550.050 622.050 ;
        RECT 575.400 619.050 576.450 631.950 ;
        RECT 584.400 631.050 585.450 665.400 ;
        RECT 583.950 628.950 586.050 631.050 ;
        RECT 583.950 626.850 586.050 627.750 ;
        RECT 586.950 626.250 589.050 627.150 ;
        RECT 586.950 622.950 589.050 625.050 ;
        RECT 574.950 616.950 577.050 619.050 ;
        RECT 539.250 593.400 540.450 605.400 ;
        RECT 541.950 604.950 544.050 607.050 ;
        RECT 541.950 602.250 544.050 603.150 ;
        RECT 575.400 601.050 576.450 616.950 ;
        RECT 577.950 601.950 580.050 604.050 ;
        RECT 587.400 601.050 588.450 622.950 ;
        RECT 592.950 605.400 595.050 607.500 ;
        RECT 541.950 598.950 544.050 601.050 ;
        RECT 568.950 598.950 571.050 601.050 ;
        RECT 574.950 598.950 577.050 601.050 ;
        RECT 578.250 599.850 579.750 600.750 ;
        RECT 580.950 598.950 583.050 601.050 ;
        RECT 586.950 598.950 589.050 601.050 ;
        RECT 538.950 591.300 541.050 593.400 ;
        RECT 539.250 587.700 540.450 591.300 ;
        RECT 538.950 585.600 541.050 587.700 ;
        RECT 536.400 581.400 540.450 582.450 ;
        RECT 539.400 561.450 540.450 581.400 ;
        RECT 541.950 561.450 544.050 562.050 ;
        RECT 539.400 560.400 544.050 561.450 ;
        RECT 532.950 550.950 535.050 553.050 ;
        RECT 535.950 529.950 538.050 532.050 ;
        RECT 536.400 529.050 537.450 529.950 ;
        RECT 523.950 526.950 526.050 529.050 ;
        RECT 529.950 526.950 532.050 529.050 ;
        RECT 535.950 526.950 538.050 529.050 ;
        RECT 509.400 493.050 510.450 520.950 ;
        RECT 520.950 519.300 523.050 521.400 ;
        RECT 521.550 515.700 522.750 519.300 ;
        RECT 520.950 513.600 523.050 515.700 ;
        RECT 517.950 495.300 520.050 497.400 ;
        RECT 508.950 490.950 511.050 493.050 ;
        RECT 518.550 491.700 519.750 495.300 ;
        RECT 502.950 486.450 505.050 487.050 ;
        RECT 500.400 485.400 505.050 486.450 ;
        RECT 502.950 484.950 505.050 485.400 ;
        RECT 506.250 485.250 508.050 486.150 ;
        RECT 496.950 482.850 499.050 483.750 ;
        RECT 499.950 482.250 502.050 483.150 ;
        RECT 502.950 482.850 504.750 483.750 ;
        RECT 505.950 481.950 508.050 484.050 ;
        RECT 499.950 478.950 502.050 481.050 ;
        RECT 509.400 480.450 510.450 490.950 ;
        RECT 517.950 489.600 520.050 491.700 ;
        RECT 514.950 483.450 517.050 484.050 ;
        RECT 512.400 482.400 517.050 483.450 ;
        RECT 512.400 481.050 513.450 482.400 ;
        RECT 514.950 481.950 517.050 482.400 ;
        RECT 506.400 479.400 510.450 480.450 ;
        RECT 500.400 478.050 501.450 478.950 ;
        RECT 499.950 475.950 502.050 478.050 ;
        RECT 491.400 458.400 495.450 459.450 ;
        RECT 490.950 454.950 493.050 457.050 ;
        RECT 478.950 416.250 481.050 417.150 ;
        RECT 478.950 414.450 481.050 415.050 ;
        RECT 476.400 413.400 481.050 414.450 ;
        RECT 478.950 412.950 481.050 413.400 ;
        RECT 482.250 413.250 483.750 414.150 ;
        RECT 484.950 412.950 487.050 415.050 ;
        RECT 488.250 413.250 490.050 414.150 ;
        RECT 481.950 409.950 484.050 412.050 ;
        RECT 485.250 410.850 486.750 411.750 ;
        RECT 487.950 409.950 490.050 412.050 ;
        RECT 421.950 382.950 424.050 385.050 ;
        RECT 445.950 382.950 448.050 385.050 ;
        RECT 460.950 382.950 463.050 385.050 ;
        RECT 464.250 383.250 465.750 384.150 ;
        RECT 466.950 382.950 469.050 385.050 ;
        RECT 472.950 382.950 475.050 385.050 ;
        RECT 418.950 380.250 420.750 381.150 ;
        RECT 421.950 379.950 424.050 382.050 ;
        RECT 425.250 380.250 427.050 381.150 ;
        RECT 418.950 376.950 421.050 379.050 ;
        RECT 422.250 377.850 423.750 378.750 ;
        RECT 424.950 376.950 427.050 379.050 ;
        RECT 425.400 376.050 426.450 376.950 ;
        RECT 416.400 374.400 420.450 375.450 ;
        RECT 400.950 343.950 403.050 346.050 ;
        RECT 397.950 341.250 400.050 342.150 ;
        RECT 400.950 341.850 403.050 342.750 ;
        RECT 406.950 341.250 409.050 342.150 ;
        RECT 397.950 337.950 400.050 340.050 ;
        RECT 406.950 337.950 409.050 340.050 ;
        RECT 407.400 337.050 408.450 337.950 ;
        RECT 373.950 334.950 376.050 337.050 ;
        RECT 385.950 334.950 388.050 337.050 ;
        RECT 406.950 334.950 409.050 337.050 ;
        RECT 358.950 331.500 361.050 333.600 ;
        RECT 374.400 313.050 375.450 334.950 ;
        RECT 373.950 310.950 376.050 313.050 ;
        RECT 377.250 311.250 378.750 312.150 ;
        RECT 379.950 310.950 382.050 313.050 ;
        RECT 373.950 308.850 375.750 309.750 ;
        RECT 376.950 307.950 379.050 310.050 ;
        RECT 380.250 308.850 381.750 309.750 ;
        RECT 382.950 307.950 385.050 310.050 ;
        RECT 377.400 307.050 378.450 307.950 ;
        RECT 376.950 304.950 379.050 307.050 ;
        RECT 379.950 304.950 382.050 307.050 ;
        RECT 382.950 305.850 385.050 306.750 ;
        RECT 358.950 274.950 361.050 277.050 ;
        RECT 355.950 271.950 358.050 274.050 ;
        RECT 356.400 271.050 357.450 271.950 ;
        RECT 346.950 269.250 348.750 270.150 ;
        RECT 349.950 268.950 352.050 271.050 ;
        RECT 355.950 268.950 358.050 271.050 ;
        RECT 346.950 265.950 349.050 268.050 ;
        RECT 350.250 266.850 352.050 267.750 ;
        RECT 352.950 266.250 355.050 267.150 ;
        RECT 355.950 266.850 358.050 267.750 ;
        RECT 347.400 244.050 348.450 265.950 ;
        RECT 359.400 265.050 360.450 274.950 ;
        RECT 380.400 271.050 381.450 304.950 ;
        RECT 386.400 274.050 387.450 334.950 ;
        RECT 419.400 313.050 420.450 374.400 ;
        RECT 424.950 373.950 427.050 376.050 ;
        RECT 439.950 344.250 442.050 345.150 ;
        RECT 446.400 343.050 447.450 382.950 ;
        RECT 482.400 382.050 483.450 409.950 ;
        RECT 457.950 379.950 460.050 382.050 ;
        RECT 461.250 380.850 462.750 381.750 ;
        RECT 463.950 379.950 466.050 382.050 ;
        RECT 467.250 380.850 469.050 381.750 ;
        RECT 481.950 379.950 484.050 382.050 ;
        RECT 457.950 377.850 460.050 378.750 ;
        RECT 464.400 376.050 465.450 379.950 ;
        RECT 463.950 373.950 466.050 376.050 ;
        RECT 487.950 344.250 490.050 345.150 ;
        RECT 439.950 340.950 442.050 343.050 ;
        RECT 443.250 341.250 444.750 342.150 ;
        RECT 445.950 340.950 448.050 343.050 ;
        RECT 449.250 341.250 451.050 342.150 ;
        RECT 454.950 340.950 457.050 343.050 ;
        RECT 478.950 341.250 480.750 342.150 ;
        RECT 481.950 340.950 484.050 343.050 ;
        RECT 485.250 341.250 486.750 342.150 ;
        RECT 487.950 340.950 490.050 343.050 ;
        RECT 442.950 337.950 445.050 340.050 ;
        RECT 446.250 338.850 447.750 339.750 ;
        RECT 448.950 337.950 451.050 340.050 ;
        RECT 449.400 337.050 450.450 337.950 ;
        RECT 448.950 334.950 451.050 337.050 ;
        RECT 418.950 310.950 421.050 313.050 ;
        RECT 422.250 311.250 423.750 312.150 ;
        RECT 424.950 310.950 427.050 313.050 ;
        RECT 415.950 307.950 418.050 310.050 ;
        RECT 419.250 308.850 420.750 309.750 ;
        RECT 421.950 307.950 424.050 310.050 ;
        RECT 425.250 308.850 427.050 309.750 ;
        RECT 415.950 305.850 418.050 306.750 ;
        RECT 418.950 304.950 421.050 307.050 ;
        RECT 449.400 306.450 450.450 334.950 ;
        RECT 455.400 310.050 456.450 340.950 ;
        RECT 478.950 337.950 481.050 340.050 ;
        RECT 482.250 338.850 483.750 339.750 ;
        RECT 484.950 337.950 487.050 340.050 ;
        RECT 479.400 337.050 480.450 337.950 ;
        RECT 478.950 334.950 481.050 337.050 ;
        RECT 479.400 313.050 480.450 334.950 ;
        RECT 478.950 310.950 481.050 313.050 ;
        RECT 451.950 308.250 453.750 309.150 ;
        RECT 454.950 307.950 457.050 310.050 ;
        RECT 458.250 308.250 460.050 309.150 ;
        RECT 451.950 306.450 454.050 307.050 ;
        RECT 449.400 305.400 454.050 306.450 ;
        RECT 455.250 305.850 456.750 306.750 ;
        RECT 385.950 271.950 388.050 274.050 ;
        RECT 389.250 272.250 390.750 273.150 ;
        RECT 391.950 271.950 394.050 274.050 ;
        RECT 379.950 268.950 382.050 271.050 ;
        RECT 385.950 269.850 387.750 270.750 ;
        RECT 388.950 268.950 391.050 271.050 ;
        RECT 392.250 269.850 394.050 270.750 ;
        RECT 349.950 262.950 352.050 265.050 ;
        RECT 352.950 262.950 355.050 265.050 ;
        RECT 358.950 262.950 361.050 265.050 ;
        RECT 346.950 241.950 349.050 244.050 ;
        RECT 346.950 239.250 349.050 240.150 ;
        RECT 343.950 235.950 346.050 238.050 ;
        RECT 346.950 235.950 349.050 238.050 ;
        RECT 350.400 235.050 351.450 262.950 ;
        RECT 358.950 245.400 361.050 247.500 ;
        RECT 379.950 245.400 382.050 247.500 ;
        RECT 349.950 232.950 352.050 235.050 ;
        RECT 359.400 228.600 360.600 245.400 ;
        RECT 364.950 241.950 367.050 244.050 ;
        RECT 370.950 241.950 373.050 244.050 ;
        RECT 365.400 241.050 366.450 241.950 ;
        RECT 371.400 241.050 372.450 241.950 ;
        RECT 364.950 238.950 367.050 241.050 ;
        RECT 370.950 240.450 373.050 241.050 ;
        RECT 368.400 239.400 373.050 240.450 ;
        RECT 368.400 238.050 369.450 239.400 ;
        RECT 370.950 238.950 373.050 239.400 ;
        RECT 364.950 236.850 367.050 237.750 ;
        RECT 367.950 235.950 370.050 238.050 ;
        RECT 370.950 236.850 373.050 237.750 ;
        RECT 367.950 232.950 370.050 235.050 ;
        RECT 380.250 233.400 381.450 245.400 ;
        RECT 385.950 244.950 388.050 247.050 ;
        RECT 382.950 242.250 385.050 243.150 ;
        RECT 382.950 240.450 385.050 241.050 ;
        RECT 386.400 240.450 387.450 244.950 ;
        RECT 382.950 239.400 387.450 240.450 ;
        RECT 382.950 238.950 385.050 239.400 ;
        RECT 409.950 238.950 412.050 241.050 ;
        RECT 358.950 226.500 361.050 228.600 ;
        RECT 337.950 197.250 340.050 198.150 ;
        RECT 343.950 197.250 346.050 198.150 ;
        RECT 343.950 193.950 346.050 196.050 ;
        RECT 307.950 190.950 310.050 193.050 ;
        RECT 316.950 190.950 319.050 193.050 ;
        RECT 344.400 190.050 345.450 193.950 ;
        RECT 304.950 187.950 307.050 190.050 ;
        RECT 343.950 187.950 346.050 190.050 ;
        RECT 364.950 172.950 367.050 175.050 ;
        RECT 322.950 169.950 325.050 172.050 ;
        RECT 323.400 169.050 324.450 169.950 ;
        RECT 283.950 166.950 286.050 169.050 ;
        RECT 289.950 166.950 292.050 169.050 ;
        RECT 301.950 166.950 304.050 169.050 ;
        RECT 322.950 166.950 325.050 169.050 ;
        RECT 325.950 166.950 328.050 169.050 ;
        RECT 328.950 166.950 331.050 169.050 ;
        RECT 349.950 166.950 352.050 169.050 ;
        RECT 283.950 164.850 286.050 165.750 ;
        RECT 289.950 164.850 292.050 165.750 ;
        RECT 322.950 164.850 325.050 165.750 ;
        RECT 277.950 134.400 280.050 136.500 ;
        RECT 298.950 135.300 301.050 137.400 ;
        RECT 268.950 127.950 271.050 130.050 ;
        RECT 262.950 125.250 265.050 126.150 ;
        RECT 268.950 125.250 271.050 126.150 ;
        RECT 262.950 121.950 265.050 124.050 ;
        RECT 266.250 122.250 267.750 123.150 ;
        RECT 268.950 121.950 271.050 124.050 ;
        RECT 262.950 118.950 265.050 121.050 ;
        RECT 265.950 118.950 268.050 121.050 ;
        RECT 263.400 97.050 264.450 118.950 ;
        RECT 269.400 100.050 270.450 121.950 ;
        RECT 278.400 117.600 279.600 134.400 ;
        RECT 299.250 131.700 300.450 135.300 ;
        RECT 286.950 127.950 289.050 130.050 ;
        RECT 298.950 129.600 301.050 131.700 ;
        RECT 283.950 125.250 286.050 126.150 ;
        RECT 283.950 121.950 286.050 124.050 ;
        RECT 287.400 123.450 288.450 127.950 ;
        RECT 289.950 125.250 292.050 126.150 ;
        RECT 289.950 123.450 292.050 124.050 ;
        RECT 287.400 122.400 292.050 123.450 ;
        RECT 289.950 121.950 292.050 122.400 ;
        RECT 277.950 115.500 280.050 117.600 ;
        RECT 284.400 115.050 285.450 121.950 ;
        RECT 299.250 117.600 300.450 129.600 ;
        RECT 301.950 121.950 304.050 124.050 ;
        RECT 326.400 121.050 327.450 166.950 ;
        RECT 328.950 164.850 331.050 165.750 ;
        RECT 334.950 125.250 337.050 126.150 ;
        RECT 340.950 125.250 343.050 126.150 ;
        RECT 334.950 121.950 337.050 124.050 ;
        RECT 338.250 122.250 339.750 123.150 ;
        RECT 340.950 121.950 343.050 124.050 ;
        RECT 341.400 121.050 342.450 121.950 ;
        RECT 301.950 119.850 304.050 120.750 ;
        RECT 325.950 118.950 328.050 121.050 ;
        RECT 337.950 118.950 340.050 121.050 ;
        RECT 340.950 118.950 343.050 121.050 ;
        RECT 298.950 115.500 301.050 117.600 ;
        RECT 283.950 112.950 286.050 115.050 ;
        RECT 298.950 100.950 301.050 103.050 ;
        RECT 299.400 100.050 300.450 100.950 ;
        RECT 268.950 97.950 271.050 100.050 ;
        RECT 295.950 97.950 298.050 100.050 ;
        RECT 298.950 97.950 301.050 100.050 ;
        RECT 301.950 97.950 304.050 100.050 ;
        RECT 262.950 94.950 265.050 97.050 ;
        RECT 266.250 95.250 267.750 96.150 ;
        RECT 268.950 94.950 271.050 97.050 ;
        RECT 271.950 94.950 274.050 97.050 ;
        RECT 259.950 91.950 262.050 94.050 ;
        RECT 263.250 92.850 264.750 93.750 ;
        RECT 265.950 91.950 268.050 94.050 ;
        RECT 269.250 92.850 271.050 93.750 ;
        RECT 259.950 89.850 262.050 90.750 ;
        RECT 265.950 88.950 268.050 91.050 ;
        RECT 266.400 55.050 267.450 88.950 ;
        RECT 265.950 52.950 268.050 55.050 ;
        RECT 262.950 50.250 265.050 51.150 ;
        RECT 265.950 50.850 268.050 51.750 ;
        RECT 262.950 46.950 265.050 49.050 ;
        RECT 263.400 46.050 264.450 46.950 ;
        RECT 262.950 43.950 265.050 46.050 ;
        RECT 272.400 34.050 273.450 94.950 ;
        RECT 289.950 55.950 292.050 58.050 ;
        RECT 290.400 46.050 291.450 55.950 ;
        RECT 296.400 55.050 297.450 97.950 ;
        RECT 302.400 97.050 303.450 97.950 ;
        RECT 298.950 95.850 300.750 96.750 ;
        RECT 301.950 94.950 304.050 97.050 ;
        RECT 307.950 95.250 310.050 96.150 ;
        RECT 301.950 92.850 304.050 93.750 ;
        RECT 307.950 91.950 310.050 94.050 ;
        RECT 308.400 91.050 309.450 91.950 ;
        RECT 307.950 88.950 310.050 91.050 ;
        RECT 298.950 55.950 301.050 58.050 ;
        RECT 304.950 57.450 307.050 58.050 ;
        RECT 302.250 56.250 303.750 57.150 ;
        RECT 304.950 56.400 309.450 57.450 ;
        RECT 304.950 55.950 307.050 56.400 ;
        RECT 295.950 52.950 298.050 55.050 ;
        RECT 298.950 53.850 300.750 54.750 ;
        RECT 301.950 52.950 304.050 55.050 ;
        RECT 305.250 53.850 307.050 54.750 ;
        RECT 308.400 49.050 309.450 56.400 ;
        RECT 326.400 55.050 327.450 118.950 ;
        RECT 338.400 103.050 339.450 118.950 ;
        RECT 334.950 100.950 337.050 103.050 ;
        RECT 337.950 100.950 340.050 103.050 ;
        RECT 335.400 93.450 336.450 100.950 ;
        RECT 340.950 97.950 343.050 100.050 ;
        RECT 346.950 97.950 349.050 100.050 ;
        RECT 347.400 97.050 348.450 97.950 ;
        RECT 337.950 95.250 340.050 96.150 ;
        RECT 340.950 95.850 343.050 96.750 ;
        RECT 343.950 95.250 345.750 96.150 ;
        RECT 346.950 94.950 349.050 97.050 ;
        RECT 350.400 94.050 351.450 166.950 ;
        RECT 365.400 166.050 366.450 172.950 ;
        RECT 368.400 169.050 369.450 232.950 ;
        RECT 379.950 231.300 382.050 233.400 ;
        RECT 403.950 232.950 406.050 235.050 ;
        RECT 380.250 227.700 381.450 231.300 ;
        RECT 379.950 225.600 382.050 227.700 ;
        RECT 373.950 199.950 376.050 202.050 ;
        RECT 374.400 169.050 375.450 199.950 ;
        RECT 376.950 197.250 379.050 198.150 ;
        RECT 382.950 197.250 385.050 198.150 ;
        RECT 382.950 193.950 385.050 196.050 ;
        RECT 383.400 175.050 384.450 193.950 ;
        RECT 382.950 172.950 385.050 175.050 ;
        RECT 379.950 169.950 382.050 172.050 ;
        RECT 367.950 166.950 370.050 169.050 ;
        RECT 371.250 167.250 372.750 168.150 ;
        RECT 373.950 166.950 376.050 169.050 ;
        RECT 376.950 166.950 379.050 169.050 ;
        RECT 364.950 165.450 367.050 166.050 ;
        RECT 362.400 164.400 367.050 165.450 ;
        RECT 368.250 164.850 369.750 165.750 ;
        RECT 362.400 127.050 363.450 164.400 ;
        RECT 364.950 163.950 367.050 164.400 ;
        RECT 370.950 163.950 373.050 166.050 ;
        RECT 374.250 164.850 376.050 165.750 ;
        RECT 364.950 161.850 367.050 162.750 ;
        RECT 377.400 133.050 378.450 166.950 ;
        RECT 380.400 166.050 381.450 169.950 ;
        RECT 379.950 163.950 382.050 166.050 ;
        RECT 370.950 130.950 373.050 133.050 ;
        RECT 376.950 130.950 379.050 133.050 ;
        RECT 361.950 124.950 364.050 127.050 ;
        RECT 362.400 112.050 363.450 124.950 ;
        RECT 371.400 123.450 372.450 130.950 ;
        RECT 373.950 128.250 376.050 129.150 ;
        RECT 380.400 127.050 381.450 163.950 ;
        RECT 373.950 124.950 376.050 127.050 ;
        RECT 377.250 125.250 378.750 126.150 ;
        RECT 379.950 124.950 382.050 127.050 ;
        RECT 383.250 125.250 385.050 126.150 ;
        RECT 404.400 124.050 405.450 232.950 ;
        RECT 410.400 172.050 411.450 238.950 ;
        RECT 419.400 238.050 420.450 304.950 ;
        RECT 439.950 279.300 442.050 281.400 ;
        RECT 436.950 274.950 439.050 277.050 ;
        RECT 440.550 275.700 441.750 279.300 ;
        RECT 449.400 277.050 450.450 305.400 ;
        RECT 451.950 304.950 454.050 305.400 ;
        RECT 457.950 304.950 460.050 307.050 ;
        RECT 427.950 271.950 430.050 274.050 ;
        RECT 428.400 271.050 429.450 271.950 ;
        RECT 427.950 268.950 430.050 271.050 ;
        RECT 437.400 268.050 438.450 274.950 ;
        RECT 439.950 273.600 442.050 275.700 ;
        RECT 448.950 274.950 451.050 277.050 ;
        RECT 427.950 266.850 430.050 267.750 ;
        RECT 430.950 266.250 433.050 267.150 ;
        RECT 436.950 265.950 439.050 268.050 ;
        RECT 430.950 262.950 433.050 265.050 ;
        RECT 436.950 263.850 439.050 264.750 ;
        RECT 431.400 247.050 432.450 262.950 ;
        RECT 440.550 261.600 441.750 273.600 ;
        RECT 448.950 269.250 451.050 270.150 ;
        RECT 454.950 269.250 457.050 270.150 ;
        RECT 448.950 265.950 451.050 268.050 ;
        RECT 454.950 265.950 457.050 268.050 ;
        RECT 439.950 259.500 442.050 261.600 ;
        RECT 430.950 244.950 433.050 247.050 ;
        RECT 433.950 245.400 436.050 247.500 ;
        RECT 415.950 236.250 417.750 237.150 ;
        RECT 418.950 235.950 421.050 238.050 ;
        RECT 422.250 236.250 424.050 237.150 ;
        RECT 415.950 232.950 418.050 235.050 ;
        RECT 419.250 233.850 420.750 234.750 ;
        RECT 421.950 232.950 424.050 235.050 ;
        RECT 416.400 232.050 417.450 232.950 ;
        RECT 415.950 229.950 418.050 232.050 ;
        RECT 434.400 228.600 435.600 245.400 ;
        RECT 449.400 244.050 450.450 265.950 ;
        RECT 458.400 262.050 459.450 304.950 ;
        RECT 460.950 278.400 463.050 280.500 ;
        RECT 457.950 259.950 460.050 262.050 ;
        RECT 461.400 261.600 462.600 278.400 ;
        RECT 479.400 265.050 480.450 310.950 ;
        RECT 478.950 262.950 481.050 265.050 ;
        RECT 460.950 259.500 463.050 261.600 ;
        RECT 478.950 259.950 481.050 262.050 ;
        RECT 454.950 245.400 457.050 247.500 ;
        RECT 445.950 241.950 448.050 244.050 ;
        RECT 448.950 241.950 451.050 244.050 ;
        RECT 446.400 241.050 447.450 241.950 ;
        RECT 439.950 238.950 442.050 241.050 ;
        RECT 445.950 238.950 448.050 241.050 ;
        RECT 439.950 236.850 442.050 237.750 ;
        RECT 445.950 236.850 448.050 237.750 ;
        RECT 455.250 233.400 456.450 245.400 ;
        RECT 457.950 242.250 460.050 243.150 ;
        RECT 457.950 238.950 460.050 241.050 ;
        RECT 458.400 235.050 459.450 238.950 ;
        RECT 454.950 231.300 457.050 233.400 ;
        RECT 457.950 232.950 460.050 235.050 ;
        RECT 433.950 226.500 436.050 228.600 ;
        RECT 455.250 227.700 456.450 231.300 ;
        RECT 454.950 225.600 457.050 227.700 ;
        RECT 479.400 199.050 480.450 259.950 ;
        RECT 488.400 253.050 489.450 340.950 ;
        RECT 491.400 319.050 492.450 454.950 ;
        RECT 494.400 412.050 495.450 458.400 ;
        RECT 506.400 457.050 507.450 479.400 ;
        RECT 499.950 454.950 502.050 457.050 ;
        RECT 505.950 454.950 508.050 457.050 ;
        RECT 499.950 452.850 502.050 453.750 ;
        RECT 505.950 452.850 508.050 453.750 ;
        RECT 509.400 451.050 510.450 479.400 ;
        RECT 511.950 478.950 514.050 481.050 ;
        RECT 514.950 479.850 517.050 480.750 ;
        RECT 511.950 475.950 514.050 478.050 ;
        RECT 518.550 477.600 519.750 489.600 ;
        RECT 524.400 483.450 525.450 526.950 ;
        RECT 529.950 524.850 532.050 525.750 ;
        RECT 535.950 524.850 538.050 525.750 ;
        RECT 539.400 523.050 540.450 560.400 ;
        RECT 541.950 559.950 544.050 560.400 ;
        RECT 545.250 560.250 546.750 561.150 ;
        RECT 547.950 559.950 550.050 562.050 ;
        RECT 541.950 557.850 543.750 558.750 ;
        RECT 544.950 556.950 547.050 559.050 ;
        RECT 548.250 557.850 550.050 558.750 ;
        RECT 545.400 553.050 546.450 556.950 ;
        RECT 544.950 550.950 547.050 553.050 ;
        RECT 541.950 533.400 544.050 535.500 ;
        RECT 538.950 520.950 541.050 523.050 ;
        RECT 542.400 516.600 543.600 533.400 ;
        RECT 565.950 523.950 568.050 526.050 ;
        RECT 566.400 523.050 567.450 523.950 ;
        RECT 565.950 520.950 568.050 523.050 ;
        RECT 541.950 514.500 544.050 516.600 ;
        RECT 538.950 494.400 541.050 496.500 ;
        RECT 526.950 485.250 529.050 486.150 ;
        RECT 532.950 485.250 535.050 486.150 ;
        RECT 526.950 483.450 529.050 484.050 ;
        RECT 524.400 482.400 529.050 483.450 ;
        RECT 526.950 481.950 529.050 482.400 ;
        RECT 532.950 481.950 535.050 484.050 ;
        RECT 539.400 477.600 540.600 494.400 ;
        RECT 550.950 481.950 553.050 484.050 ;
        RECT 508.950 448.950 511.050 451.050 ;
        RECT 493.950 409.950 496.050 412.050 ;
        RECT 509.400 409.050 510.450 448.950 ;
        RECT 508.950 406.950 511.050 409.050 ;
        RECT 499.950 397.950 502.050 400.050 ;
        RECT 500.400 388.050 501.450 397.950 ;
        RECT 499.950 385.950 502.050 388.050 ;
        RECT 496.950 383.250 499.050 384.150 ;
        RECT 499.950 383.850 502.050 384.750 ;
        RECT 505.950 384.450 508.050 385.050 ;
        RECT 502.950 383.250 504.750 384.150 ;
        RECT 505.950 383.400 510.450 384.450 ;
        RECT 505.950 382.950 508.050 383.400 ;
        RECT 496.950 381.450 499.050 382.050 ;
        RECT 494.400 380.400 499.050 381.450 ;
        RECT 490.950 316.950 493.050 319.050 ;
        RECT 491.400 313.050 492.450 316.950 ;
        RECT 490.950 310.950 493.050 313.050 ;
        RECT 490.950 308.850 493.050 309.750 ;
        RECT 494.400 259.050 495.450 380.400 ;
        RECT 496.950 379.950 499.050 380.400 ;
        RECT 502.950 379.950 505.050 382.050 ;
        RECT 506.250 380.850 508.050 381.750 ;
        RECT 496.950 373.950 499.050 376.050 ;
        RECT 497.400 313.050 498.450 373.950 ;
        RECT 509.400 343.050 510.450 383.400 ;
        RECT 512.400 376.050 513.450 475.950 ;
        RECT 517.950 475.500 520.050 477.600 ;
        RECT 538.950 475.500 541.050 477.600 ;
        RECT 544.950 457.950 547.050 460.050 ;
        RECT 545.400 457.050 546.450 457.950 ;
        RECT 551.400 457.050 552.450 481.950 ;
        RECT 544.950 454.950 547.050 457.050 ;
        RECT 548.250 455.250 549.750 456.150 ;
        RECT 550.950 454.950 553.050 457.050 ;
        RECT 566.400 454.050 567.450 520.950 ;
        RECT 541.950 451.950 544.050 454.050 ;
        RECT 545.250 452.850 546.750 453.750 ;
        RECT 547.950 451.950 550.050 454.050 ;
        RECT 551.250 452.850 553.050 453.750 ;
        RECT 565.950 451.950 568.050 454.050 ;
        RECT 548.400 451.050 549.450 451.950 ;
        RECT 541.950 449.850 544.050 450.750 ;
        RECT 547.950 448.950 550.050 451.050 ;
        RECT 569.400 448.050 570.450 598.950 ;
        RECT 574.950 596.850 577.050 597.750 ;
        RECT 580.950 596.850 583.050 597.750 ;
        RECT 593.400 588.600 594.600 605.400 ;
        RECT 598.950 604.950 601.050 607.050 ;
        RECT 599.400 601.050 600.450 604.950 ;
        RECT 598.950 598.950 601.050 601.050 ;
        RECT 604.950 600.450 607.050 601.050 ;
        RECT 602.400 599.400 607.050 600.450 ;
        RECT 598.950 596.850 601.050 597.750 ;
        RECT 592.950 586.500 595.050 588.600 ;
        RECT 574.950 565.950 577.050 568.050 ;
        RECT 571.950 556.950 574.050 559.050 ;
        RECT 572.400 475.050 573.450 556.950 ;
        RECT 575.400 487.050 576.450 565.950 ;
        RECT 580.950 557.250 582.750 558.150 ;
        RECT 583.950 556.950 586.050 559.050 ;
        RECT 589.950 558.450 592.050 559.050 ;
        RECT 589.950 557.400 594.450 558.450 ;
        RECT 589.950 556.950 592.050 557.400 ;
        RECT 593.400 556.050 594.450 557.400 ;
        RECT 580.950 553.950 583.050 556.050 ;
        RECT 584.250 554.850 586.050 555.750 ;
        RECT 586.950 554.250 589.050 555.150 ;
        RECT 589.950 554.850 592.050 555.750 ;
        RECT 592.950 553.950 595.050 556.050 ;
        RECT 581.400 532.050 582.450 553.950 ;
        RECT 586.950 550.950 589.050 553.050 ;
        RECT 589.950 550.950 592.050 553.050 ;
        RECT 580.950 529.950 583.050 532.050 ;
        RECT 580.950 524.250 582.750 525.150 ;
        RECT 583.950 523.950 586.050 526.050 ;
        RECT 587.250 524.250 589.050 525.150 ;
        RECT 580.950 520.950 583.050 523.050 ;
        RECT 584.250 521.850 585.750 522.750 ;
        RECT 586.950 520.950 589.050 523.050 ;
        RECT 590.400 492.450 591.450 550.950 ;
        RECT 595.950 533.400 598.050 535.500 ;
        RECT 592.950 530.250 595.050 531.150 ;
        RECT 592.950 526.950 595.050 529.050 ;
        RECT 593.400 523.050 594.450 526.950 ;
        RECT 592.950 520.950 595.050 523.050 ;
        RECT 596.550 521.400 597.750 533.400 ;
        RECT 602.400 529.050 603.450 599.400 ;
        RECT 604.950 598.950 607.050 599.400 ;
        RECT 604.950 596.850 607.050 597.750 ;
        RECT 611.400 562.050 612.450 673.950 ;
        RECT 613.950 670.950 616.050 673.050 ;
        RECT 620.400 672.450 621.450 700.950 ;
        RECT 664.950 697.950 667.050 700.050 ;
        RECT 665.400 697.050 666.450 697.950 ;
        RECT 689.400 697.050 690.450 704.400 ;
        RECT 691.950 703.950 694.050 704.400 ;
        RECT 695.250 704.250 696.750 705.150 ;
        RECT 691.950 701.850 693.750 702.750 ;
        RECT 694.950 700.950 697.050 703.050 ;
        RECT 698.250 701.850 700.050 702.750 ;
        RECT 733.950 701.250 736.050 702.150 ;
        RECT 739.950 700.950 742.050 703.050 ;
        RECT 748.950 700.950 751.050 703.050 ;
        RECT 658.950 694.950 661.050 697.050 ;
        RECT 664.950 694.950 667.050 697.050 ;
        RECT 688.950 694.950 691.050 697.050 ;
        RECT 617.400 671.400 621.450 672.450 ;
        RECT 614.400 634.050 615.450 670.950 ;
        RECT 617.400 670.050 618.450 671.400 ;
        RECT 622.950 670.950 625.050 673.050 ;
        RECT 623.400 670.050 624.450 670.950 ;
        RECT 616.950 667.950 619.050 670.050 ;
        RECT 619.950 668.250 621.750 669.150 ;
        RECT 622.950 667.950 625.050 670.050 ;
        RECT 626.250 668.250 628.050 669.150 ;
        RECT 628.950 667.950 631.050 670.050 ;
        RECT 617.400 666.450 618.450 667.950 ;
        RECT 619.950 666.450 622.050 667.050 ;
        RECT 617.400 665.400 622.050 666.450 ;
        RECT 623.250 665.850 624.750 666.750 ;
        RECT 625.950 666.450 628.050 667.050 ;
        RECT 629.400 666.450 630.450 667.950 ;
        RECT 659.400 667.050 660.450 694.950 ;
        RECT 664.950 670.950 667.050 673.050 ;
        RECT 670.950 670.950 673.050 673.050 ;
        RECT 665.400 670.050 666.450 670.950 ;
        RECT 661.950 668.250 663.750 669.150 ;
        RECT 664.950 667.950 667.050 670.050 ;
        RECT 668.250 668.250 670.050 669.150 ;
        RECT 619.950 664.950 622.050 665.400 ;
        RECT 625.950 665.400 630.450 666.450 ;
        RECT 625.950 664.950 628.050 665.400 ;
        RECT 658.950 664.950 661.050 667.050 ;
        RECT 661.950 664.950 664.050 667.050 ;
        RECT 665.250 665.850 666.750 666.750 ;
        RECT 667.950 664.950 670.050 667.050 ;
        RECT 662.400 664.050 663.450 664.950 ;
        RECT 649.950 661.950 652.050 664.050 ;
        RECT 661.950 661.950 664.050 664.050 ;
        RECT 613.950 631.950 616.050 634.050 ;
        RECT 619.950 631.950 622.050 634.050 ;
        RECT 613.950 629.250 616.050 630.150 ;
        RECT 619.950 629.850 622.050 630.750 ;
        RECT 622.950 629.250 625.050 630.150 ;
        RECT 650.400 628.050 651.450 661.950 ;
        RECT 664.950 632.250 667.050 633.150 ;
        RECT 652.950 628.950 655.050 631.050 ;
        RECT 655.950 629.250 657.750 630.150 ;
        RECT 658.950 628.950 661.050 631.050 ;
        RECT 662.250 629.250 663.750 630.150 ;
        RECT 664.950 628.950 667.050 631.050 ;
        RECT 613.950 625.950 616.050 628.050 ;
        RECT 622.950 625.950 625.050 628.050 ;
        RECT 649.950 625.950 652.050 628.050 ;
        RECT 614.400 625.050 615.450 625.950 ;
        RECT 613.950 622.950 616.050 625.050 ;
        RECT 613.950 605.400 616.050 607.500 ;
        RECT 614.250 593.400 615.450 605.400 ;
        RECT 616.950 602.250 619.050 603.150 ;
        RECT 619.950 601.950 622.050 604.050 ;
        RECT 616.950 598.950 619.050 601.050 ;
        RECT 613.950 591.300 616.050 593.400 ;
        RECT 614.250 587.700 615.450 591.300 ;
        RECT 613.950 585.600 616.050 587.700 ;
        RECT 620.400 573.450 621.450 601.950 ;
        RECT 617.400 572.400 621.450 573.450 ;
        RECT 610.950 559.950 613.050 562.050 ;
        RECT 617.400 555.450 618.450 572.400 ;
        RECT 623.400 559.050 624.450 625.950 ;
        RECT 650.400 589.050 651.450 625.950 ;
        RECT 653.400 624.450 654.450 628.950 ;
        RECT 655.950 625.950 658.050 628.050 ;
        RECT 659.250 626.850 660.750 627.750 ;
        RECT 661.950 625.950 664.050 628.050 ;
        RECT 653.400 623.400 657.450 624.450 ;
        RECT 656.400 598.050 657.450 623.400 ;
        RECT 662.400 607.050 663.450 625.950 ;
        RECT 661.950 604.950 664.050 607.050 ;
        RECT 668.400 601.050 669.450 664.950 ;
        RECT 671.400 631.050 672.450 670.950 ;
        RECT 695.400 667.050 696.450 700.950 ;
        RECT 730.950 698.250 732.750 699.150 ;
        RECT 739.950 698.850 742.050 699.750 ;
        RECT 727.950 696.450 730.050 697.050 ;
        RECT 730.950 696.450 733.050 697.050 ;
        RECT 727.950 695.400 733.050 696.450 ;
        RECT 727.950 694.950 730.050 695.400 ;
        RECT 730.950 694.950 733.050 695.400 ;
        RECT 697.950 673.950 700.050 676.050 ;
        RECT 697.950 671.850 699.750 672.750 ;
        RECT 706.950 671.250 709.050 672.150 ;
        RECT 700.950 668.850 703.050 669.750 ;
        RECT 706.950 667.950 709.050 670.050 ;
        RECT 709.950 667.950 712.050 670.050 ;
        RECT 694.950 664.950 697.050 667.050 ;
        RECT 670.950 628.950 673.050 631.050 ;
        RECT 688.950 628.950 691.050 631.050 ;
        RECT 697.950 628.950 700.050 631.050 ;
        RECT 667.950 598.950 670.050 601.050 ;
        RECT 652.950 596.250 654.750 597.150 ;
        RECT 655.950 595.950 658.050 598.050 ;
        RECT 659.250 596.250 661.050 597.150 ;
        RECT 652.950 592.950 655.050 595.050 ;
        RECT 656.250 593.850 657.750 594.750 ;
        RECT 658.950 592.950 661.050 595.050 ;
        RECT 670.950 592.950 673.050 595.050 ;
        RECT 689.400 594.450 690.450 628.950 ;
        RECT 697.950 626.850 700.050 627.750 ;
        RECT 700.950 626.250 703.050 627.150 ;
        RECT 700.950 622.950 703.050 625.050 ;
        RECT 691.950 596.250 693.750 597.150 ;
        RECT 694.950 595.950 697.050 598.050 ;
        RECT 698.250 596.250 700.050 597.150 ;
        RECT 691.950 594.450 694.050 595.050 ;
        RECT 689.400 593.400 694.050 594.450 ;
        RECT 695.250 593.850 696.750 594.750 ;
        RECT 691.950 592.950 694.050 593.400 ;
        RECT 697.950 592.950 700.050 595.050 ;
        RECT 649.950 586.950 652.050 589.050 ;
        RECT 628.950 560.250 631.050 561.150 ;
        RECT 649.950 559.950 652.050 562.050 ;
        RECT 661.950 561.450 664.050 562.050 ;
        RECT 659.400 560.400 664.050 561.450 ;
        RECT 619.950 557.250 621.750 558.150 ;
        RECT 622.950 556.950 625.050 559.050 ;
        RECT 626.250 557.250 627.750 558.150 ;
        RECT 628.950 556.950 631.050 559.050 ;
        RECT 619.950 555.450 622.050 556.050 ;
        RECT 617.400 554.400 622.050 555.450 ;
        RECT 623.250 554.850 624.750 555.750 ;
        RECT 619.950 553.950 622.050 554.400 ;
        RECT 625.950 553.950 628.050 556.050 ;
        RECT 616.950 533.400 619.050 535.500 ;
        RECT 601.950 526.950 604.050 529.050 ;
        RECT 604.950 526.950 607.050 529.050 ;
        RECT 610.950 528.450 613.050 529.050 ;
        RECT 610.950 527.400 615.450 528.450 ;
        RECT 610.950 526.950 613.050 527.400 ;
        RECT 595.950 519.300 598.050 521.400 ;
        RECT 596.550 515.700 597.750 519.300 ;
        RECT 595.950 513.600 598.050 515.700 ;
        RECT 595.950 495.300 598.050 497.400 ;
        RECT 590.400 491.400 594.450 492.450 ;
        RECT 596.550 491.700 597.750 495.300 ;
        RECT 580.950 487.950 583.050 490.050 ;
        RECT 589.950 487.950 592.050 490.050 ;
        RECT 581.400 487.050 582.450 487.950 ;
        RECT 574.950 484.950 577.050 487.050 ;
        RECT 580.950 484.950 583.050 487.050 ;
        RECT 584.250 485.250 586.050 486.150 ;
        RECT 574.950 482.850 577.050 483.750 ;
        RECT 577.950 482.250 580.050 483.150 ;
        RECT 580.950 482.850 582.750 483.750 ;
        RECT 583.950 481.950 586.050 484.050 ;
        RECT 577.950 478.950 580.050 481.050 ;
        RECT 571.950 472.950 574.050 475.050 ;
        RECT 544.950 445.950 547.050 448.050 ;
        RECT 568.950 445.950 571.050 448.050 ;
        RECT 520.950 413.250 523.050 414.150 ;
        RECT 526.950 413.250 529.050 414.150 ;
        RECT 532.950 412.950 535.050 415.050 ;
        RECT 520.950 409.950 523.050 412.050 ;
        RECT 524.250 410.250 525.750 411.150 ;
        RECT 526.950 409.950 529.050 412.050 ;
        RECT 523.950 406.950 526.050 409.050 ;
        RECT 524.400 400.050 525.450 406.950 ;
        RECT 523.950 397.950 526.050 400.050 ;
        RECT 527.400 391.050 528.450 409.950 ;
        RECT 526.950 388.950 529.050 391.050 ;
        RECT 533.400 382.050 534.450 412.950 ;
        RECT 545.400 385.050 546.450 445.950 ;
        RECT 562.950 415.950 565.050 418.050 ;
        RECT 563.400 415.050 564.450 415.950 ;
        RECT 556.950 413.250 559.050 414.150 ;
        RECT 562.950 412.950 565.050 415.050 ;
        RECT 553.950 410.250 555.750 411.150 ;
        RECT 556.950 409.950 559.050 412.050 ;
        RECT 562.950 410.850 565.050 411.750 ;
        RECT 553.950 406.950 556.050 409.050 ;
        RECT 554.400 391.050 555.450 406.950 ;
        RECT 550.950 388.950 553.050 391.050 ;
        RECT 553.950 388.950 556.050 391.050 ;
        RECT 551.400 385.050 552.450 388.950 ;
        RECT 572.400 388.050 573.450 472.950 ;
        RECT 556.950 385.950 559.050 388.050 ;
        RECT 571.950 385.950 574.050 388.050 ;
        RECT 544.950 382.950 547.050 385.050 ;
        RECT 548.250 383.250 549.750 384.150 ;
        RECT 550.950 382.950 553.050 385.050 ;
        RECT 532.950 379.950 535.050 382.050 ;
        RECT 541.950 379.950 544.050 382.050 ;
        RECT 545.250 380.850 546.750 381.750 ;
        RECT 547.950 379.950 550.050 382.050 ;
        RECT 551.250 380.850 553.050 381.750 ;
        RECT 511.950 373.950 514.050 376.050 ;
        RECT 508.950 340.950 511.050 343.050 ;
        RECT 520.950 341.250 523.050 342.150 ;
        RECT 526.950 341.250 529.050 342.150 ;
        RECT 520.950 337.950 523.050 340.050 ;
        RECT 533.400 313.050 534.450 379.950 ;
        RECT 541.950 377.850 544.050 378.750 ;
        RECT 548.400 360.450 549.450 379.950 ;
        RECT 545.400 359.400 549.450 360.450 ;
        RECT 538.950 351.300 541.050 353.400 ;
        RECT 539.550 347.700 540.750 351.300 ;
        RECT 538.950 345.600 541.050 347.700 ;
        RECT 535.950 337.950 538.050 340.050 ;
        RECT 535.950 335.850 538.050 336.750 ;
        RECT 539.550 333.600 540.750 345.600 ;
        RECT 538.950 331.500 541.050 333.600 ;
        RECT 496.950 310.950 499.050 313.050 ;
        RECT 532.950 310.950 535.050 313.050 ;
        RECT 541.950 310.950 544.050 313.050 ;
        RECT 496.950 308.850 499.050 309.750 ;
        RECT 532.950 308.850 535.050 309.750 ;
        RECT 535.950 308.250 538.050 309.150 ;
        RECT 541.950 308.850 544.050 309.750 ;
        RECT 535.950 304.950 538.050 307.050 ;
        RECT 514.950 301.950 517.050 304.050 ;
        RECT 502.950 271.950 505.050 274.050 ;
        RECT 499.950 269.250 502.050 270.150 ;
        RECT 502.950 269.850 505.050 270.750 ;
        RECT 508.950 269.250 511.050 270.150 ;
        RECT 515.400 268.050 516.450 301.950 ;
        RECT 536.400 301.050 537.450 304.950 ;
        RECT 541.950 301.950 544.050 304.050 ;
        RECT 535.950 298.950 538.050 301.050 ;
        RECT 517.950 279.300 520.050 281.400 ;
        RECT 518.550 275.700 519.750 279.300 ;
        RECT 538.950 278.400 541.050 280.500 ;
        RECT 517.950 273.600 520.050 275.700 ;
        RECT 499.950 265.950 502.050 268.050 ;
        RECT 508.950 265.950 511.050 268.050 ;
        RECT 514.950 265.950 517.050 268.050 ;
        RECT 509.400 265.050 510.450 265.950 ;
        RECT 508.950 262.950 511.050 265.050 ;
        RECT 514.950 263.850 517.050 264.750 ;
        RECT 493.950 256.950 496.050 259.050 ;
        RECT 487.950 250.950 490.050 253.050 ;
        RECT 493.950 250.950 496.050 253.050 ;
        RECT 494.400 238.050 495.450 250.950 ;
        RECT 490.950 236.250 492.750 237.150 ;
        RECT 493.950 235.950 496.050 238.050 ;
        RECT 497.250 236.250 499.050 237.150 ;
        RECT 509.400 235.050 510.450 262.950 ;
        RECT 518.550 261.600 519.750 273.600 ;
        RECT 529.950 271.950 532.050 274.050 ;
        RECT 526.950 269.250 529.050 270.150 ;
        RECT 526.950 265.950 529.050 268.050 ;
        RECT 527.400 262.050 528.450 265.950 ;
        RECT 517.950 259.500 520.050 261.600 ;
        RECT 526.950 259.950 529.050 262.050 ;
        RECT 527.400 244.050 528.450 259.950 ;
        RECT 526.950 241.950 529.050 244.050 ;
        RECT 530.400 238.050 531.450 271.950 ;
        RECT 532.950 269.250 535.050 270.150 ;
        RECT 532.950 265.950 535.050 268.050 ;
        RECT 533.400 265.050 534.450 265.950 ;
        RECT 532.950 262.950 535.050 265.050 ;
        RECT 539.400 261.600 540.600 278.400 ;
        RECT 538.950 259.500 541.050 261.600 ;
        RECT 532.950 238.950 535.050 241.050 ;
        RECT 538.950 240.450 541.050 241.050 ;
        RECT 542.400 240.450 543.450 301.950 ;
        RECT 536.250 239.250 537.750 240.150 ;
        RECT 538.950 239.400 543.450 240.450 ;
        RECT 538.950 238.950 541.050 239.400 ;
        RECT 529.950 237.450 532.050 238.050 ;
        RECT 527.400 236.400 532.050 237.450 ;
        RECT 533.250 236.850 534.750 237.750 ;
        RECT 490.950 232.950 493.050 235.050 ;
        RECT 494.250 233.850 495.750 234.750 ;
        RECT 496.950 232.950 499.050 235.050 ;
        RECT 508.950 232.950 511.050 235.050 ;
        RECT 415.950 197.250 418.050 198.150 ;
        RECT 421.950 197.250 424.050 198.150 ;
        RECT 457.950 197.250 460.050 198.150 ;
        RECT 463.950 197.250 466.050 198.150 ;
        RECT 478.950 196.950 481.050 199.050 ;
        RECT 415.950 193.950 418.050 196.050 ;
        RECT 421.950 193.950 424.050 196.050 ;
        RECT 457.950 193.950 460.050 196.050 ;
        RECT 461.250 194.250 462.750 195.150 ;
        RECT 463.950 193.950 466.050 196.050 ;
        RECT 416.400 193.050 417.450 193.950 ;
        RECT 415.950 190.950 418.050 193.050 ;
        RECT 412.950 172.950 415.050 175.050 ;
        RECT 409.950 169.950 412.050 172.050 ;
        RECT 413.400 169.050 414.450 172.950 ;
        RECT 406.950 166.950 409.050 169.050 ;
        RECT 410.250 167.850 411.750 168.750 ;
        RECT 412.950 166.950 415.050 169.050 ;
        RECT 406.950 164.850 409.050 165.750 ;
        RECT 412.950 164.850 415.050 165.750 ;
        RECT 422.400 129.450 423.450 193.950 ;
        RECT 445.950 169.950 448.050 172.050 ;
        RECT 442.950 167.250 445.050 168.150 ;
        RECT 445.950 167.850 448.050 168.750 ;
        RECT 448.950 167.250 450.750 168.150 ;
        RECT 451.950 166.950 454.050 169.050 ;
        RECT 442.950 163.950 445.050 166.050 ;
        RECT 448.950 163.950 451.050 166.050 ;
        RECT 452.250 164.850 454.050 165.750 ;
        RECT 443.400 163.050 444.450 163.950 ;
        RECT 442.950 160.950 445.050 163.050 ;
        RECT 458.400 150.450 459.450 193.950 ;
        RECT 460.950 190.950 463.050 193.050 ;
        RECT 461.400 175.050 462.450 190.950 ;
        RECT 475.950 175.950 478.050 178.050 ;
        RECT 460.950 172.950 463.050 175.050 ;
        RECT 463.950 173.400 466.050 175.500 ;
        RECT 464.400 156.600 465.600 173.400 ;
        RECT 476.400 169.050 477.450 175.950 ;
        RECT 469.950 166.950 472.050 169.050 ;
        RECT 475.950 166.950 478.050 169.050 ;
        RECT 469.950 164.850 472.050 165.750 ;
        RECT 475.950 164.850 478.050 165.750 ;
        RECT 479.400 163.050 480.450 196.950 ;
        RECT 491.400 196.050 492.450 232.950 ;
        RECT 497.400 232.050 498.450 232.950 ;
        RECT 496.950 229.950 499.050 232.050 ;
        RECT 527.400 199.050 528.450 236.400 ;
        RECT 529.950 235.950 532.050 236.400 ;
        RECT 535.950 235.950 538.050 238.050 ;
        RECT 539.250 236.850 541.050 237.750 ;
        RECT 529.950 233.850 532.050 234.750 ;
        RECT 536.400 234.450 537.450 235.950 ;
        RECT 536.400 233.400 540.450 234.450 ;
        RECT 532.950 200.250 535.050 201.150 ;
        RECT 539.400 199.050 540.450 233.400 ;
        RECT 496.950 196.950 499.050 199.050 ;
        RECT 526.950 196.950 529.050 199.050 ;
        RECT 532.950 196.950 535.050 199.050 ;
        RECT 536.250 197.250 537.750 198.150 ;
        RECT 538.950 196.950 541.050 199.050 ;
        RECT 542.250 197.250 544.050 198.150 ;
        RECT 490.950 193.950 493.050 196.050 ;
        RECT 493.950 194.250 496.050 195.150 ;
        RECT 496.950 194.850 499.050 195.750 ;
        RECT 493.950 190.950 496.050 193.050 ;
        RECT 481.950 175.950 484.050 178.050 ;
        RECT 478.950 160.950 481.050 163.050 ;
        RECT 463.950 154.500 466.050 156.600 ;
        RECT 458.400 149.400 462.450 150.450 ;
        RECT 424.950 130.950 427.050 133.050 ;
        RECT 425.400 129.450 426.450 130.950 ;
        RECT 451.950 129.450 454.050 130.050 ;
        RECT 422.400 128.400 426.450 129.450 ;
        RECT 412.950 125.250 414.750 126.150 ;
        RECT 415.950 124.950 418.050 127.050 ;
        RECT 421.950 124.950 424.050 127.050 ;
        RECT 376.950 123.450 379.050 124.050 ;
        RECT 371.400 122.400 379.050 123.450 ;
        RECT 380.250 122.850 381.750 123.750 ;
        RECT 376.950 121.950 379.050 122.400 ;
        RECT 382.950 121.950 385.050 124.050 ;
        RECT 403.950 121.950 406.050 124.050 ;
        RECT 412.950 121.950 415.050 124.050 ;
        RECT 416.250 122.850 418.050 123.750 ;
        RECT 418.950 122.250 421.050 123.150 ;
        RECT 421.950 122.850 424.050 123.750 ;
        RECT 383.400 118.050 384.450 121.950 ;
        RECT 382.950 115.950 385.050 118.050 ;
        RECT 361.950 109.950 364.050 112.050 ;
        RECT 337.950 93.450 340.050 94.050 ;
        RECT 335.400 92.400 340.050 93.450 ;
        RECT 337.950 91.950 340.050 92.400 ;
        RECT 343.950 91.950 346.050 94.050 ;
        RECT 347.250 92.850 349.050 93.750 ;
        RECT 349.950 91.950 352.050 94.050 ;
        RECT 343.950 56.250 346.050 57.150 ;
        RECT 325.950 52.950 328.050 55.050 ;
        RECT 334.950 53.250 336.750 54.150 ;
        RECT 337.950 52.950 340.050 55.050 ;
        RECT 341.250 53.250 342.750 54.150 ;
        RECT 343.950 52.950 346.050 55.050 ;
        RECT 344.400 52.050 345.450 52.950 ;
        RECT 334.950 49.950 337.050 52.050 ;
        RECT 338.250 50.850 339.750 51.750 ;
        RECT 340.950 49.950 343.050 52.050 ;
        RECT 343.950 49.950 346.050 52.050 ;
        RECT 307.950 46.950 310.050 49.050 ;
        RECT 289.950 43.950 292.050 46.050 ;
        RECT 271.950 31.950 274.050 34.050 ;
        RECT 262.950 29.400 265.050 31.500 ;
        RECT 335.400 31.050 336.450 49.950 ;
        RECT 253.950 25.950 256.050 28.050 ;
        RECT 254.400 25.050 255.450 25.950 ;
        RECT 247.950 22.950 250.050 25.050 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 247.950 20.850 250.050 21.750 ;
        RECT 253.950 20.850 256.050 21.750 ;
        RECT 263.250 17.400 264.450 29.400 ;
        RECT 268.950 28.950 271.050 31.050 ;
        RECT 334.950 28.950 337.050 31.050 ;
        RECT 265.950 26.250 268.050 27.150 ;
        RECT 265.950 24.450 268.050 25.050 ;
        RECT 269.400 24.450 270.450 28.950 ;
        RECT 307.950 25.950 310.050 28.050 ;
        RECT 313.950 25.950 316.050 28.050 ;
        RECT 316.950 25.950 319.050 28.050 ;
        RECT 341.400 27.450 342.450 49.950 ;
        RECT 338.400 26.400 342.450 27.450 ;
        RECT 265.950 23.400 270.450 24.450 ;
        RECT 265.950 22.950 268.050 23.400 ;
        RECT 301.950 22.950 304.050 25.050 ;
        RECT 305.250 23.250 307.050 24.150 ;
        RECT 307.950 23.850 310.050 24.750 ;
        RECT 310.950 23.250 313.050 24.150 ;
        RECT 301.950 20.850 303.750 21.750 ;
        RECT 304.950 19.950 307.050 22.050 ;
        RECT 310.950 19.950 313.050 22.050 ;
        RECT 314.400 19.050 315.450 25.950 ;
        RECT 317.400 22.050 318.450 25.950 ;
        RECT 338.400 25.050 339.450 26.400 ;
        RECT 343.950 25.950 346.050 28.050 ;
        RECT 346.950 25.950 349.050 28.050 ;
        RECT 347.400 25.050 348.450 25.950 ;
        RECT 350.400 25.050 351.450 91.950 ;
        RECT 362.400 52.050 363.450 109.950 ;
        RECT 413.400 100.050 414.450 121.950 ;
        RECT 425.400 121.050 426.450 128.400 ;
        RECT 449.400 128.400 454.050 129.450 ;
        RECT 418.950 118.950 421.050 121.050 ;
        RECT 424.950 118.950 427.050 121.050 ;
        RECT 449.400 118.050 450.450 128.400 ;
        RECT 451.950 127.950 454.050 128.400 ;
        RECT 455.250 128.250 456.750 129.150 ;
        RECT 457.950 127.950 460.050 130.050 ;
        RECT 451.950 125.850 453.750 126.750 ;
        RECT 454.950 124.950 457.050 127.050 ;
        RECT 458.250 125.850 460.050 126.750 ;
        RECT 430.950 115.950 433.050 118.050 ;
        RECT 448.950 115.950 451.050 118.050 ;
        RECT 424.950 112.950 427.050 115.050 ;
        RECT 421.950 100.950 424.050 103.050 ;
        RECT 382.950 97.950 385.050 100.050 ;
        RECT 412.950 97.950 415.050 100.050 ;
        RECT 422.400 97.050 423.450 100.950 ;
        RECT 425.400 100.050 426.450 112.950 ;
        RECT 424.950 97.950 427.050 100.050 ;
        RECT 379.950 95.250 382.050 96.150 ;
        RECT 382.950 95.850 385.050 96.750 ;
        RECT 385.950 95.250 387.750 96.150 ;
        RECT 388.950 94.950 391.050 97.050 ;
        RECT 418.950 94.950 421.050 97.050 ;
        RECT 421.950 94.950 424.050 97.050 ;
        RECT 425.250 95.850 426.750 96.750 ;
        RECT 427.950 94.950 430.050 97.050 ;
        RECT 379.950 91.950 382.050 94.050 ;
        RECT 385.950 91.950 388.050 94.050 ;
        RECT 389.250 92.850 391.050 93.750 ;
        RECT 391.950 91.950 394.050 94.050 ;
        RECT 380.400 91.050 381.450 91.950 ;
        RECT 379.950 88.950 382.050 91.050 ;
        RECT 379.950 85.950 382.050 88.050 ;
        RECT 380.400 55.050 381.450 85.950 ;
        RECT 385.950 56.250 388.050 57.150 ;
        RECT 392.400 55.050 393.450 91.950 ;
        RECT 376.950 53.250 378.750 54.150 ;
        RECT 379.950 52.950 382.050 55.050 ;
        RECT 385.950 54.450 388.050 55.050 ;
        RECT 383.250 53.250 384.750 54.150 ;
        RECT 385.950 53.400 390.450 54.450 ;
        RECT 385.950 52.950 388.050 53.400 ;
        RECT 361.950 49.950 364.050 52.050 ;
        RECT 376.950 49.950 379.050 52.050 ;
        RECT 380.250 50.850 381.750 51.750 ;
        RECT 382.950 49.950 385.050 52.050 ;
        RECT 385.950 49.950 388.050 52.050 ;
        RECT 362.400 25.050 363.450 49.950 ;
        RECT 377.400 46.050 378.450 49.950 ;
        RECT 376.950 43.950 379.050 46.050 ;
        RECT 379.950 28.950 382.050 31.050 ;
        RECT 380.400 25.050 381.450 28.950 ;
        RECT 386.400 25.050 387.450 49.950 ;
        RECT 389.400 25.050 390.450 53.400 ;
        RECT 391.950 52.950 394.050 55.050 ;
        RECT 419.400 52.050 420.450 94.950 ;
        RECT 421.950 92.850 424.050 93.750 ;
        RECT 427.950 92.850 430.050 93.750 ;
        RECT 427.950 57.450 430.050 58.050 ;
        RECT 431.400 57.450 432.450 115.950 ;
        RECT 461.400 88.050 462.450 149.400 ;
        RECT 466.950 121.950 469.050 124.050 ;
        RECT 463.950 109.950 466.050 112.050 ;
        RECT 464.400 94.050 465.450 109.950 ;
        RECT 467.400 97.050 468.450 121.950 ;
        RECT 482.400 109.050 483.450 175.950 ;
        RECT 484.950 173.400 487.050 175.500 ;
        RECT 485.250 161.400 486.450 173.400 ;
        RECT 487.950 170.250 490.050 171.150 ;
        RECT 487.950 168.450 490.050 169.050 ;
        RECT 494.400 168.450 495.450 190.950 ;
        RECT 527.400 190.050 528.450 196.950 ;
        RECT 535.950 193.950 538.050 196.050 ;
        RECT 539.250 194.850 540.750 195.750 ;
        RECT 541.950 193.950 544.050 196.050 ;
        RECT 536.400 193.050 537.450 193.950 ;
        RECT 535.950 190.950 538.050 193.050 ;
        RECT 526.950 187.950 529.050 190.050 ;
        RECT 502.950 178.950 505.050 181.050 ;
        RECT 487.950 167.400 495.450 168.450 ;
        RECT 487.950 166.950 490.050 167.400 ;
        RECT 484.950 159.300 487.050 161.400 ;
        RECT 485.250 155.700 486.450 159.300 ;
        RECT 484.950 153.600 487.050 155.700 ;
        RECT 490.950 127.950 493.050 130.050 ;
        RECT 491.400 127.050 492.450 127.950 ;
        RECT 490.950 124.950 493.050 127.050 ;
        RECT 496.950 125.250 499.050 126.150 ;
        RECT 490.950 122.850 493.050 123.750 ;
        RECT 496.950 121.950 499.050 124.050 ;
        RECT 500.250 122.250 502.050 123.150 ;
        RECT 497.400 111.450 498.450 121.950 ;
        RECT 499.950 120.450 502.050 121.050 ;
        RECT 503.400 120.450 504.450 178.950 ;
        RECT 517.950 168.450 520.050 169.050 ;
        RECT 515.400 167.400 520.050 168.450 ;
        RECT 515.400 124.050 516.450 167.400 ;
        RECT 517.950 166.950 520.050 167.400 ;
        RECT 521.250 167.250 522.750 168.150 ;
        RECT 523.950 166.950 526.050 169.050 ;
        RECT 527.400 166.050 528.450 187.950 ;
        RECT 545.400 181.050 546.450 359.400 ;
        RECT 547.950 341.250 550.050 342.150 ;
        RECT 553.950 341.250 556.050 342.150 ;
        RECT 547.950 337.950 550.050 340.050 ;
        RECT 553.950 339.450 556.050 340.050 ;
        RECT 557.400 339.450 558.450 385.950 ;
        RECT 559.950 350.400 562.050 352.500 ;
        RECT 553.950 338.400 558.450 339.450 ;
        RECT 553.950 337.950 556.050 338.400 ;
        RECT 548.400 262.050 549.450 337.950 ;
        RECT 560.400 333.600 561.600 350.400 ;
        RECT 559.950 331.500 562.050 333.600 ;
        RECT 578.400 310.050 579.450 478.950 ;
        RECT 584.400 463.050 585.450 481.950 ;
        RECT 590.400 478.050 591.450 487.950 ;
        RECT 593.400 484.050 594.450 491.400 ;
        RECT 595.950 489.600 598.050 491.700 ;
        RECT 592.950 481.950 595.050 484.050 ;
        RECT 592.950 479.850 595.050 480.750 ;
        RECT 589.950 475.950 592.050 478.050 ;
        RECT 596.550 477.600 597.750 489.600 ;
        RECT 602.400 483.450 603.450 526.950 ;
        RECT 604.950 524.850 607.050 525.750 ;
        RECT 610.950 524.850 613.050 525.750 ;
        RECT 604.950 485.250 607.050 486.150 ;
        RECT 610.950 485.250 613.050 486.150 ;
        RECT 614.400 484.050 615.450 527.400 ;
        RECT 617.400 516.600 618.600 533.400 ;
        RECT 616.950 514.500 619.050 516.600 ;
        RECT 616.950 494.400 619.050 496.500 ;
        RECT 604.950 483.450 607.050 484.050 ;
        RECT 602.400 482.400 607.050 483.450 ;
        RECT 604.950 481.950 607.050 482.400 ;
        RECT 610.950 481.950 613.050 484.050 ;
        RECT 613.950 481.950 616.050 484.050 ;
        RECT 611.400 478.050 612.450 481.950 ;
        RECT 595.950 475.500 598.050 477.600 ;
        RECT 610.950 475.950 613.050 478.050 ;
        RECT 617.400 477.600 618.600 494.400 ;
        RECT 616.950 475.500 619.050 477.600 ;
        RECT 622.950 475.950 625.050 478.050 ;
        RECT 583.950 460.950 586.050 463.050 ;
        RECT 595.950 460.950 598.050 463.050 ;
        RECT 601.950 460.950 604.050 463.050 ;
        RECT 586.950 457.950 589.050 460.050 ;
        RECT 587.400 457.050 588.450 457.950 ;
        RECT 586.950 454.950 589.050 457.050 ;
        RECT 590.250 455.250 591.750 456.150 ;
        RECT 592.950 454.950 595.050 457.050 ;
        RECT 583.950 451.950 586.050 454.050 ;
        RECT 587.250 452.850 588.750 453.750 ;
        RECT 589.950 451.950 592.050 454.050 ;
        RECT 593.250 452.850 595.050 453.750 ;
        RECT 583.950 449.850 586.050 450.750 ;
        RECT 596.400 414.450 597.450 460.950 ;
        RECT 602.400 454.050 603.450 460.950 ;
        RECT 619.950 457.950 622.050 460.050 ;
        RECT 620.400 454.050 621.450 457.950 ;
        RECT 623.400 457.050 624.450 475.950 ;
        RECT 629.400 463.050 630.450 556.950 ;
        RECT 646.950 523.950 649.050 526.050 ;
        RECT 647.400 493.050 648.450 523.950 ;
        RECT 650.400 523.050 651.450 559.950 ;
        RECT 659.400 553.050 660.450 560.400 ;
        RECT 661.950 559.950 664.050 560.400 ;
        RECT 665.250 560.250 666.750 561.150 ;
        RECT 667.950 559.950 670.050 562.050 ;
        RECT 671.400 559.050 672.450 592.950 ;
        RECT 701.400 562.050 702.450 622.950 ;
        RECT 703.950 592.950 706.050 595.050 ;
        RECT 700.950 559.950 703.050 562.050 ;
        RECT 704.400 559.050 705.450 592.950 ;
        RECT 661.950 557.850 663.750 558.750 ;
        RECT 664.950 556.950 667.050 559.050 ;
        RECT 668.250 557.850 670.050 558.750 ;
        RECT 670.950 556.950 673.050 559.050 ;
        RECT 703.950 556.950 706.050 559.050 ;
        RECT 703.950 554.850 706.050 555.750 ;
        RECT 706.950 554.250 709.050 555.150 ;
        RECT 658.950 550.950 661.050 553.050 ;
        RECT 706.950 550.950 709.050 553.050 ;
        RECT 710.400 532.050 711.450 667.950 ;
        RECT 728.400 625.050 729.450 694.950 ;
        RECT 739.950 668.250 741.750 669.150 ;
        RECT 742.950 667.950 745.050 670.050 ;
        RECT 746.250 668.250 748.050 669.150 ;
        RECT 739.950 664.950 742.050 667.050 ;
        RECT 743.250 665.850 744.750 666.750 ;
        RECT 745.950 666.450 748.050 667.050 ;
        RECT 749.400 666.450 750.450 700.950 ;
        RECT 745.950 665.400 750.450 666.450 ;
        RECT 745.950 664.950 748.050 665.400 ;
        RECT 733.950 630.450 736.050 631.050 ;
        RECT 731.400 629.400 736.050 630.450 ;
        RECT 727.950 622.950 730.050 625.050 ;
        RECT 718.950 601.950 721.050 604.050 ;
        RECT 727.950 601.950 730.050 604.050 ;
        RECT 719.400 532.050 720.450 601.950 ;
        RECT 731.400 601.050 732.450 629.400 ;
        RECT 733.950 628.950 736.050 629.400 ;
        RECT 733.950 626.850 736.050 627.750 ;
        RECT 736.950 626.250 739.050 627.150 ;
        RECT 724.950 600.450 727.050 601.050 ;
        RECT 722.400 599.400 727.050 600.450 ;
        RECT 728.250 599.850 729.750 600.750 ;
        RECT 722.400 595.050 723.450 599.400 ;
        RECT 724.950 598.950 727.050 599.400 ;
        RECT 730.950 598.950 733.050 601.050 ;
        RECT 724.950 596.850 727.050 597.750 ;
        RECT 730.950 596.850 733.050 597.750 ;
        RECT 721.950 592.950 724.050 595.050 ;
        RECT 736.950 557.250 739.050 558.150 ;
        RECT 742.950 557.250 745.050 558.150 ;
        RECT 736.950 553.950 739.050 556.050 ;
        RECT 740.250 554.250 741.750 555.150 ;
        RECT 737.400 553.050 738.450 553.950 ;
        RECT 736.950 550.950 739.050 553.050 ;
        RECT 739.950 550.950 742.050 553.050 ;
        RECT 652.950 531.450 655.050 532.050 ;
        RECT 652.950 530.400 657.450 531.450 ;
        RECT 652.950 529.950 655.050 530.400 ;
        RECT 656.400 526.050 657.450 530.400 ;
        RECT 661.950 529.950 664.050 532.050 ;
        RECT 691.950 529.950 694.050 532.050 ;
        RECT 709.950 529.950 712.050 532.050 ;
        RECT 718.950 529.950 721.050 532.050 ;
        RECT 733.950 529.950 736.050 532.050 ;
        RECT 736.950 529.950 739.050 532.050 ;
        RECT 652.950 524.250 654.750 525.150 ;
        RECT 655.950 523.950 658.050 526.050 ;
        RECT 659.250 524.250 661.050 525.150 ;
        RECT 662.400 523.050 663.450 529.950 ;
        RECT 691.950 527.850 694.050 528.750 ;
        RECT 694.950 527.250 697.050 528.150 ;
        RECT 730.950 527.250 733.050 528.150 ;
        RECT 733.950 527.850 736.050 528.750 ;
        RECT 694.950 523.950 697.050 526.050 ;
        RECT 730.950 523.950 733.050 526.050 ;
        RECT 649.950 520.950 652.050 523.050 ;
        RECT 652.950 520.950 655.050 523.050 ;
        RECT 656.250 521.850 657.750 522.750 ;
        RECT 658.950 520.950 661.050 523.050 ;
        RECT 661.950 520.950 664.050 523.050 ;
        RECT 649.950 517.950 652.050 520.050 ;
        RECT 646.950 490.950 649.050 493.050 ;
        RECT 650.400 487.050 651.450 517.950 ;
        RECT 659.400 514.050 660.450 520.950 ;
        RECT 658.950 511.950 661.050 514.050 ;
        RECT 655.950 490.950 658.050 493.050 ;
        RECT 656.400 487.050 657.450 490.950 ;
        RECT 649.950 484.950 652.050 487.050 ;
        RECT 652.950 485.250 654.750 486.150 ;
        RECT 655.950 484.950 658.050 487.050 ;
        RECT 659.250 485.250 660.750 486.150 ;
        RECT 661.950 484.950 664.050 487.050 ;
        RECT 665.250 485.250 667.050 486.150 ;
        RECT 685.950 484.950 688.050 487.050 ;
        RECT 652.950 481.950 655.050 484.050 ;
        RECT 656.250 482.850 657.750 483.750 ;
        RECT 658.950 481.950 661.050 484.050 ;
        RECT 662.250 482.850 663.750 483.750 ;
        RECT 664.950 481.950 667.050 484.050 ;
        RECT 628.950 460.950 631.050 463.050 ;
        RECT 629.400 460.050 630.450 460.950 ;
        RECT 628.950 457.950 631.050 460.050 ;
        RECT 637.950 457.950 640.050 460.050 ;
        RECT 622.950 454.950 625.050 457.050 ;
        RECT 626.250 455.250 628.050 456.150 ;
        RECT 628.950 455.850 631.050 456.750 ;
        RECT 631.950 455.250 634.050 456.150 ;
        RECT 601.950 451.950 604.050 454.050 ;
        RECT 619.950 451.950 622.050 454.050 ;
        RECT 622.950 452.850 624.750 453.750 ;
        RECT 625.950 451.950 628.050 454.050 ;
        RECT 631.950 451.950 634.050 454.050 ;
        RECT 638.400 418.050 639.450 457.950 ;
        RECT 598.950 416.250 601.050 417.150 ;
        RECT 604.950 415.950 607.050 418.050 ;
        RECT 637.950 415.950 640.050 418.050 ;
        RECT 641.250 416.250 642.750 417.150 ;
        RECT 643.950 415.950 646.050 418.050 ;
        RECT 605.400 415.050 606.450 415.950 ;
        RECT 598.950 414.450 601.050 415.050 ;
        RECT 596.400 413.400 601.050 414.450 ;
        RECT 598.950 412.950 601.050 413.400 ;
        RECT 602.250 413.250 603.750 414.150 ;
        RECT 604.950 412.950 607.050 415.050 ;
        RECT 608.250 413.250 610.050 414.150 ;
        RECT 637.950 413.850 639.750 414.750 ;
        RECT 640.950 412.950 643.050 415.050 ;
        RECT 644.250 413.850 646.050 414.750 ;
        RECT 601.950 409.950 604.050 412.050 ;
        RECT 605.250 410.850 606.750 411.750 ;
        RECT 607.950 409.950 610.050 412.050 ;
        RECT 610.950 409.950 613.050 412.050 ;
        RECT 595.950 388.950 598.050 391.050 ;
        RECT 583.950 385.950 586.050 388.050 ;
        RECT 586.950 385.950 589.050 388.050 ;
        RECT 584.400 385.050 585.450 385.950 ;
        RECT 583.950 382.950 586.050 385.050 ;
        RECT 587.250 383.850 588.750 384.750 ;
        RECT 589.950 384.450 592.050 385.050 ;
        RECT 589.950 383.400 594.450 384.450 ;
        RECT 589.950 382.950 592.050 383.400 ;
        RECT 583.950 380.850 586.050 381.750 ;
        RECT 589.950 380.850 592.050 381.750 ;
        RECT 589.950 376.950 592.050 379.050 ;
        RECT 590.400 343.050 591.450 376.950 ;
        RECT 593.400 376.050 594.450 383.400 ;
        RECT 592.950 373.950 595.050 376.050 ;
        RECT 589.950 340.950 592.050 343.050 ;
        RECT 586.950 310.950 589.050 313.050 ;
        RECT 574.950 308.250 576.750 309.150 ;
        RECT 577.950 307.950 580.050 310.050 ;
        RECT 581.250 308.250 583.050 309.150 ;
        RECT 587.400 307.050 588.450 310.950 ;
        RECT 574.950 304.950 577.050 307.050 ;
        RECT 578.250 305.850 579.750 306.750 ;
        RECT 580.950 304.950 583.050 307.050 ;
        RECT 586.950 304.950 589.050 307.050 ;
        RECT 581.400 301.050 582.450 304.950 ;
        RECT 580.950 298.950 583.050 301.050 ;
        RECT 553.950 279.300 556.050 281.400 ;
        RECT 554.550 275.700 555.750 279.300 ;
        RECT 574.950 278.400 577.050 280.500 ;
        RECT 553.950 273.600 556.050 275.700 ;
        RECT 550.950 265.950 553.050 268.050 ;
        RECT 550.950 263.850 553.050 264.750 ;
        RECT 547.950 259.950 550.050 262.050 ;
        RECT 554.550 261.600 555.750 273.600 ;
        RECT 562.950 269.250 565.050 270.150 ;
        RECT 568.950 269.250 571.050 270.150 ;
        RECT 556.950 265.950 559.050 268.050 ;
        RECT 562.950 265.950 565.050 268.050 ;
        RECT 568.950 265.950 571.050 268.050 ;
        RECT 553.950 259.500 556.050 261.600 ;
        RECT 557.400 256.050 558.450 265.950 ;
        RECT 563.400 262.050 564.450 265.950 ;
        RECT 562.950 259.950 565.050 262.050 ;
        RECT 556.950 253.950 559.050 256.050 ;
        RECT 547.950 244.950 550.050 247.050 ;
        RECT 548.400 202.050 549.450 244.950 ;
        RECT 553.950 241.950 556.050 244.050 ;
        RECT 550.950 207.300 553.050 209.400 ;
        RECT 551.550 203.700 552.750 207.300 ;
        RECT 547.950 199.950 550.050 202.050 ;
        RECT 550.950 201.600 553.050 203.700 ;
        RECT 548.400 196.050 549.450 199.950 ;
        RECT 547.950 193.950 550.050 196.050 ;
        RECT 547.950 191.850 550.050 192.750 ;
        RECT 551.550 189.600 552.750 201.600 ;
        RECT 554.400 199.050 555.450 241.950 ;
        RECT 557.400 199.050 558.450 253.950 ;
        RECT 569.400 250.050 570.450 265.950 ;
        RECT 571.950 262.950 574.050 265.050 ;
        RECT 568.950 247.950 571.050 250.050 ;
        RECT 572.400 241.050 573.450 262.950 ;
        RECT 575.400 261.600 576.600 278.400 ;
        RECT 574.950 259.500 577.050 261.600 ;
        RECT 581.400 259.050 582.450 298.950 ;
        RECT 580.950 256.950 583.050 259.050 ;
        RECT 583.950 250.950 586.050 253.050 ;
        RECT 577.950 241.950 580.050 244.050 ;
        RECT 571.950 238.950 574.050 241.050 ;
        RECT 575.250 239.250 577.050 240.150 ;
        RECT 577.950 239.850 580.050 240.750 ;
        RECT 580.950 239.250 583.050 240.150 ;
        RECT 571.950 236.850 573.750 237.750 ;
        RECT 574.950 235.950 577.050 238.050 ;
        RECT 580.950 237.450 583.050 238.050 ;
        RECT 584.400 237.450 585.450 250.950 ;
        RECT 580.950 236.400 585.450 237.450 ;
        RECT 580.950 235.950 583.050 236.400 ;
        RECT 571.950 206.400 574.050 208.500 ;
        RECT 568.950 199.950 571.050 202.050 ;
        RECT 553.950 196.950 556.050 199.050 ;
        RECT 556.950 196.950 559.050 199.050 ;
        RECT 559.950 197.250 562.050 198.150 ;
        RECT 565.950 197.250 568.050 198.150 ;
        RECT 550.950 187.500 553.050 189.600 ;
        RECT 544.950 178.950 547.050 181.050 ;
        RECT 517.950 164.850 519.750 165.750 ;
        RECT 520.950 163.950 523.050 166.050 ;
        RECT 524.250 164.850 525.750 165.750 ;
        RECT 526.950 163.950 529.050 166.050 ;
        RECT 529.950 163.950 532.050 166.050 ;
        RECT 521.400 163.050 522.450 163.950 ;
        RECT 520.950 160.950 523.050 163.050 ;
        RECT 526.950 161.850 529.050 162.750 ;
        RECT 530.400 126.450 531.450 163.950 ;
        RECT 554.400 133.050 555.450 196.950 ;
        RECT 559.950 193.950 562.050 196.050 ;
        RECT 565.950 193.950 568.050 196.050 ;
        RECT 560.400 178.050 561.450 193.950 ;
        RECT 566.400 190.050 567.450 193.950 ;
        RECT 565.950 187.950 568.050 190.050 ;
        RECT 559.950 175.950 562.050 178.050 ;
        RECT 569.400 169.050 570.450 199.950 ;
        RECT 572.400 189.600 573.600 206.400 ;
        RECT 571.950 187.500 574.050 189.600 ;
        RECT 562.950 166.950 565.050 169.050 ;
        RECT 566.250 167.250 567.750 168.150 ;
        RECT 568.950 166.950 571.050 169.050 ;
        RECT 559.950 163.950 562.050 166.050 ;
        RECT 563.250 164.850 564.750 165.750 ;
        RECT 565.950 163.950 568.050 166.050 ;
        RECT 569.250 164.850 571.050 165.750 ;
        RECT 559.950 161.850 562.050 162.750 ;
        RECT 566.400 133.050 567.450 163.950 ;
        RECT 587.400 160.050 588.450 304.950 ;
        RECT 593.400 271.050 594.450 373.950 ;
        RECT 592.950 268.950 595.050 271.050 ;
        RECT 586.950 157.950 589.050 160.050 ;
        RECT 538.950 130.950 541.050 133.050 ;
        RECT 553.950 130.950 556.050 133.050 ;
        RECT 565.950 130.950 568.050 133.050 ;
        RECT 532.950 128.250 535.050 129.150 ;
        RECT 539.400 127.050 540.450 130.950 ;
        RECT 532.950 126.450 535.050 127.050 ;
        RECT 530.400 125.400 535.050 126.450 ;
        RECT 532.950 124.950 535.050 125.400 ;
        RECT 536.250 125.250 537.750 126.150 ;
        RECT 538.950 124.950 541.050 127.050 ;
        RECT 542.250 125.250 544.050 126.150 ;
        RECT 566.400 124.050 567.450 130.950 ;
        RECT 568.950 124.950 571.050 127.050 ;
        RECT 571.950 125.250 573.750 126.150 ;
        RECT 574.950 124.950 577.050 127.050 ;
        RECT 580.950 124.950 583.050 127.050 ;
        RECT 514.950 121.950 517.050 124.050 ;
        RECT 535.950 121.950 538.050 124.050 ;
        RECT 539.250 122.850 540.750 123.750 ;
        RECT 541.950 121.950 544.050 124.050 ;
        RECT 550.950 121.950 553.050 124.050 ;
        RECT 565.950 121.950 568.050 124.050 ;
        RECT 536.400 121.050 537.450 121.950 ;
        RECT 499.950 119.400 504.450 120.450 ;
        RECT 499.950 118.950 502.050 119.400 ;
        RECT 497.400 110.400 501.450 111.450 ;
        RECT 481.950 106.950 484.050 109.050 ;
        RECT 490.950 106.950 493.050 109.050 ;
        RECT 481.950 101.400 484.050 103.500 ;
        RECT 478.950 98.250 481.050 99.150 ;
        RECT 466.950 94.950 469.050 97.050 ;
        RECT 470.250 95.250 471.750 96.150 ;
        RECT 472.950 94.950 475.050 97.050 ;
        RECT 478.950 94.950 481.050 97.050 ;
        RECT 463.950 91.950 466.050 94.050 ;
        RECT 467.250 92.850 468.750 93.750 ;
        RECT 469.950 91.950 472.050 94.050 ;
        RECT 473.250 92.850 475.050 93.750 ;
        RECT 463.950 89.850 466.050 90.750 ;
        RECT 470.400 88.050 471.450 91.950 ;
        RECT 460.950 85.950 463.050 88.050 ;
        RECT 469.950 85.950 472.050 88.050 ;
        RECT 425.250 56.250 426.750 57.150 ;
        RECT 427.950 56.400 432.450 57.450 ;
        RECT 427.950 55.950 430.050 56.400 ;
        RECT 421.950 53.850 423.750 54.750 ;
        RECT 424.950 52.950 427.050 55.050 ;
        RECT 428.250 53.850 430.050 54.750 ;
        RECT 418.950 49.950 421.050 52.050 ;
        RECT 431.400 49.050 432.450 56.400 ;
        RECT 466.950 55.950 469.050 58.050 ;
        RECT 467.400 55.050 468.450 55.950 ;
        RECT 460.950 53.250 463.050 54.150 ;
        RECT 466.950 52.950 469.050 55.050 ;
        RECT 457.950 50.250 459.750 51.150 ;
        RECT 466.950 50.850 469.050 51.750 ;
        RECT 479.400 49.050 480.450 94.950 ;
        RECT 482.550 89.400 483.750 101.400 ;
        RECT 491.400 97.050 492.450 106.950 ;
        RECT 496.950 97.950 499.050 100.050 ;
        RECT 497.400 97.050 498.450 97.950 ;
        RECT 490.950 94.950 493.050 97.050 ;
        RECT 496.950 94.950 499.050 97.050 ;
        RECT 490.950 92.850 493.050 93.750 ;
        RECT 496.950 92.850 499.050 93.750 ;
        RECT 481.950 87.300 484.050 89.400 ;
        RECT 482.550 83.700 483.750 87.300 ;
        RECT 481.950 81.600 484.050 83.700 ;
        RECT 500.400 52.050 501.450 110.400 ;
        RECT 503.400 108.450 504.450 119.400 ;
        RECT 535.950 118.950 538.050 121.050 ;
        RECT 541.950 115.950 544.050 118.050 ;
        RECT 503.400 107.400 507.450 108.450 ;
        RECT 502.950 101.400 505.050 103.500 ;
        RECT 503.400 84.600 504.600 101.400 ;
        RECT 506.400 91.050 507.450 107.400 ;
        RECT 542.400 94.050 543.450 115.950 ;
        RECT 538.950 92.250 540.750 93.150 ;
        RECT 541.950 91.950 544.050 94.050 ;
        RECT 545.250 92.250 547.050 93.150 ;
        RECT 505.950 88.950 508.050 91.050 ;
        RECT 538.950 88.950 541.050 91.050 ;
        RECT 542.250 89.850 543.750 90.750 ;
        RECT 544.950 88.950 547.050 91.050 ;
        RECT 547.950 88.950 550.050 91.050 ;
        RECT 502.950 82.500 505.050 84.600 ;
        RECT 502.950 55.950 505.050 58.050 ;
        RECT 506.250 56.250 507.750 57.150 ;
        RECT 508.950 55.950 511.050 58.050 ;
        RECT 502.950 53.850 504.750 54.750 ;
        RECT 505.950 52.950 508.050 55.050 ;
        RECT 509.250 53.850 511.050 54.750 ;
        RECT 506.400 52.050 507.450 52.950 ;
        RECT 539.400 52.050 540.450 88.950 ;
        RECT 548.400 58.050 549.450 88.950 ;
        RECT 551.400 88.050 552.450 121.950 ;
        RECT 569.400 121.050 570.450 124.950 ;
        RECT 571.950 121.950 574.050 124.050 ;
        RECT 575.250 122.850 577.050 123.750 ;
        RECT 577.950 122.250 580.050 123.150 ;
        RECT 580.950 122.850 583.050 123.750 ;
        RECT 568.950 118.950 571.050 121.050 ;
        RECT 568.950 106.950 571.050 109.050 ;
        RECT 556.950 101.400 559.050 103.500 ;
        RECT 550.950 85.950 553.050 88.050 ;
        RECT 557.400 84.600 558.600 101.400 ;
        RECT 569.400 97.050 570.450 106.950 ;
        RECT 572.400 97.050 573.450 121.950 ;
        RECT 577.950 118.950 580.050 121.050 ;
        RECT 577.950 101.400 580.050 103.500 ;
        RECT 562.950 94.950 565.050 97.050 ;
        RECT 568.950 94.950 571.050 97.050 ;
        RECT 571.950 94.950 574.050 97.050 ;
        RECT 562.950 92.850 565.050 93.750 ;
        RECT 568.950 92.850 571.050 93.750 ;
        RECT 578.250 89.400 579.450 101.400 ;
        RECT 580.950 98.250 583.050 99.150 ;
        RECT 580.950 94.950 583.050 97.050 ;
        RECT 577.950 87.300 580.050 89.400 ;
        RECT 581.400 88.050 582.450 94.950 ;
        RECT 596.400 91.050 597.450 388.950 ;
        RECT 608.400 382.050 609.450 409.950 ;
        RECT 607.950 379.950 610.050 382.050 ;
        RECT 598.950 344.250 601.050 345.150 ;
        RECT 598.950 340.950 601.050 343.050 ;
        RECT 602.250 341.250 603.750 342.150 ;
        RECT 604.950 340.950 607.050 343.050 ;
        RECT 608.250 341.250 610.050 342.150 ;
        RECT 601.950 337.950 604.050 340.050 ;
        RECT 605.250 338.850 606.750 339.750 ;
        RECT 607.950 337.950 610.050 340.050 ;
        RECT 602.400 274.050 603.450 337.950 ;
        RECT 608.400 337.050 609.450 337.950 ;
        RECT 607.950 334.950 610.050 337.050 ;
        RECT 611.400 306.450 612.450 409.950 ;
        RECT 619.950 385.950 622.050 388.050 ;
        RECT 619.950 383.850 622.050 384.750 ;
        RECT 622.950 383.250 625.050 384.150 ;
        RECT 653.400 382.050 654.450 481.950 ;
        RECT 670.950 457.950 673.050 460.050 ;
        RECT 661.950 452.250 663.750 453.150 ;
        RECT 664.950 451.950 667.050 454.050 ;
        RECT 668.250 452.250 670.050 453.150 ;
        RECT 661.950 448.950 664.050 451.050 ;
        RECT 665.250 449.850 666.750 450.750 ;
        RECT 667.950 448.950 670.050 451.050 ;
        RECT 662.400 435.450 663.450 448.950 ;
        RECT 659.400 434.400 663.450 435.450 ;
        RECT 659.400 415.050 660.450 434.400 ;
        RECT 661.950 415.950 664.050 418.050 ;
        RECT 662.400 415.050 663.450 415.950 ;
        RECT 658.950 412.950 661.050 415.050 ;
        RECT 661.950 412.950 664.050 415.050 ;
        RECT 662.400 385.050 663.450 412.950 ;
        RECT 671.400 409.050 672.450 457.950 ;
        RECT 679.950 454.950 682.050 457.050 ;
        RECT 680.400 415.050 681.450 454.950 ;
        RECT 673.950 412.950 676.050 415.050 ;
        RECT 679.950 412.950 682.050 415.050 ;
        RECT 683.250 413.250 685.050 414.150 ;
        RECT 673.950 410.850 676.050 411.750 ;
        RECT 676.950 410.250 679.050 411.150 ;
        RECT 679.950 410.850 681.750 411.750 ;
        RECT 682.950 411.450 685.050 412.050 ;
        RECT 686.400 411.450 687.450 484.950 ;
        RECT 695.400 481.050 696.450 523.950 ;
        RECT 712.950 511.950 715.050 514.050 ;
        RECT 703.950 487.950 706.050 490.050 ;
        RECT 704.400 487.050 705.450 487.950 ;
        RECT 697.950 484.950 700.050 487.050 ;
        RECT 703.950 484.950 706.050 487.050 ;
        RECT 707.250 485.250 709.050 486.150 ;
        RECT 697.950 482.850 700.050 483.750 ;
        RECT 700.950 482.250 703.050 483.150 ;
        RECT 703.950 482.850 705.750 483.750 ;
        RECT 706.950 481.950 709.050 484.050 ;
        RECT 709.950 481.950 712.050 484.050 ;
        RECT 694.950 478.950 697.050 481.050 ;
        RECT 700.950 478.950 703.050 481.050 ;
        RECT 706.950 457.950 709.050 460.050 ;
        RECT 710.400 457.050 711.450 481.950 ;
        RECT 713.400 481.050 714.450 511.950 ;
        RECT 731.400 490.050 732.450 523.950 ;
        RECT 733.950 490.950 736.050 493.050 ;
        RECT 730.950 487.950 733.050 490.050 ;
        RECT 727.950 484.950 730.050 487.050 ;
        RECT 712.950 478.950 715.050 481.050 ;
        RECT 728.400 463.050 729.450 484.950 ;
        RECT 734.400 484.050 735.450 490.950 ;
        RECT 733.950 481.950 736.050 484.050 ;
        RECT 727.950 460.950 730.050 463.050 ;
        RECT 712.950 457.950 715.050 460.050 ;
        RECT 703.950 454.950 706.050 457.050 ;
        RECT 707.250 455.850 708.750 456.750 ;
        RECT 709.950 454.950 712.050 457.050 ;
        RECT 703.950 452.850 706.050 453.750 ;
        RECT 709.950 452.850 712.050 453.750 ;
        RECT 713.400 451.050 714.450 457.950 ;
        RECT 712.950 448.950 715.050 451.050 ;
        RECT 709.950 412.950 712.050 415.050 ;
        RECT 715.950 414.450 718.050 415.050 ;
        RECT 713.400 413.400 718.050 414.450 ;
        RECT 682.950 410.400 687.450 411.450 ;
        RECT 682.950 409.950 685.050 410.400 ;
        RECT 670.950 406.950 673.050 409.050 ;
        RECT 676.950 406.950 679.050 409.050 ;
        RECT 703.950 406.950 706.050 409.050 ;
        RECT 670.950 385.950 673.050 388.050 ;
        RECT 697.950 385.950 700.050 388.050 ;
        RECT 658.950 382.950 661.050 385.050 ;
        RECT 661.950 382.950 664.050 385.050 ;
        RECT 667.950 384.450 670.050 385.050 ;
        RECT 671.400 384.450 672.450 385.950 ;
        RECT 665.250 383.250 666.750 384.150 ;
        RECT 667.950 383.400 672.450 384.450 ;
        RECT 697.950 383.850 700.050 384.750 ;
        RECT 667.950 382.950 670.050 383.400 ;
        RECT 659.400 382.050 660.450 382.950 ;
        RECT 622.950 379.950 625.050 382.050 ;
        RECT 652.950 379.950 655.050 382.050 ;
        RECT 658.950 379.950 661.050 382.050 ;
        RECT 662.250 380.850 663.750 381.750 ;
        RECT 664.950 379.950 667.050 382.050 ;
        RECT 668.250 380.850 670.050 381.750 ;
        RECT 665.400 379.050 666.450 379.950 ;
        RECT 658.950 377.850 661.050 378.750 ;
        RECT 664.950 376.950 667.050 379.050 ;
        RECT 652.950 343.950 655.050 346.050 ;
        RECT 640.950 341.250 643.050 342.150 ;
        RECT 646.950 341.250 649.050 342.150 ;
        RECT 640.950 337.950 643.050 340.050 ;
        RECT 644.250 338.250 645.750 339.150 ;
        RECT 646.950 337.950 649.050 340.050 ;
        RECT 641.400 337.050 642.450 337.950 ;
        RECT 640.950 334.950 643.050 337.050 ;
        RECT 643.950 334.950 646.050 337.050 ;
        RECT 619.950 315.450 622.050 316.050 ;
        RECT 617.400 314.400 622.050 315.450 ;
        RECT 617.400 310.050 618.450 314.400 ;
        RECT 619.950 313.950 622.050 314.400 ;
        RECT 622.950 313.950 625.050 316.050 ;
        RECT 613.950 308.250 615.750 309.150 ;
        RECT 616.950 307.950 619.050 310.050 ;
        RECT 620.250 308.250 622.050 309.150 ;
        RECT 613.950 306.450 616.050 307.050 ;
        RECT 611.400 305.400 616.050 306.450 ;
        RECT 617.250 305.850 618.750 306.750 ;
        RECT 619.950 306.450 622.050 307.050 ;
        RECT 623.400 306.450 624.450 313.950 ;
        RECT 641.400 310.050 642.450 334.950 ;
        RECT 644.400 316.050 645.450 334.950 ;
        RECT 653.400 316.050 654.450 343.950 ;
        RECT 671.400 343.050 672.450 383.400 ;
        RECT 700.950 383.250 703.050 384.150 ;
        RECT 700.950 381.450 703.050 382.050 ;
        RECT 704.400 381.450 705.450 406.950 ;
        RECT 710.400 382.050 711.450 412.950 ;
        RECT 713.400 412.050 714.450 413.400 ;
        RECT 715.950 412.950 718.050 413.400 ;
        RECT 721.950 412.950 724.050 415.050 ;
        RECT 725.250 413.250 727.050 414.150 ;
        RECT 712.950 409.950 715.050 412.050 ;
        RECT 715.950 410.850 718.050 411.750 ;
        RECT 718.950 410.250 721.050 411.150 ;
        RECT 721.950 410.850 723.750 411.750 ;
        RECT 724.950 411.450 727.050 412.050 ;
        RECT 728.400 411.450 729.450 460.950 ;
        RECT 734.400 454.050 735.450 481.950 ;
        RECT 737.400 459.450 738.450 529.950 ;
        RECT 740.400 493.050 741.450 550.950 ;
        RECT 739.950 490.950 742.050 493.050 ;
        RECT 748.950 488.250 751.050 489.150 ;
        RECT 739.950 485.250 741.750 486.150 ;
        RECT 742.950 484.950 745.050 487.050 ;
        RECT 746.250 485.250 747.750 486.150 ;
        RECT 748.950 484.950 751.050 487.050 ;
        RECT 739.950 481.950 742.050 484.050 ;
        RECT 743.250 482.850 744.750 483.750 ;
        RECT 745.950 481.950 748.050 484.050 ;
        RECT 746.400 481.050 747.450 481.950 ;
        RECT 745.950 478.950 748.050 481.050 ;
        RECT 748.950 460.950 751.050 463.050 ;
        RECT 737.400 458.400 741.450 459.450 ;
        RECT 737.400 457.050 738.450 458.400 ;
        RECT 740.400 457.050 741.450 458.400 ;
        RECT 745.950 457.950 748.050 460.050 ;
        RECT 746.400 457.050 747.450 457.950 ;
        RECT 736.950 454.950 739.050 457.050 ;
        RECT 739.950 454.950 742.050 457.050 ;
        RECT 743.250 455.250 744.750 456.150 ;
        RECT 745.950 454.950 748.050 457.050 ;
        RECT 749.400 454.050 750.450 460.950 ;
        RECT 733.950 451.950 736.050 454.050 ;
        RECT 739.950 452.850 741.750 453.750 ;
        RECT 742.950 451.950 745.050 454.050 ;
        RECT 746.250 452.850 747.750 453.750 ;
        RECT 748.950 451.950 751.050 454.050 ;
        RECT 748.950 449.850 751.050 450.750 ;
        RECT 724.950 410.400 729.450 411.450 ;
        RECT 724.950 409.950 727.050 410.400 ;
        RECT 718.950 406.950 721.050 409.050 ;
        RECT 730.950 387.450 733.050 388.050 ;
        RECT 728.400 386.400 733.050 387.450 ;
        RECT 728.400 385.050 729.450 386.400 ;
        RECT 730.950 385.950 733.050 386.400 ;
        RECT 727.950 382.950 730.050 385.050 ;
        RECT 730.950 383.850 733.050 384.750 ;
        RECT 733.950 383.250 736.050 384.150 ;
        RECT 700.950 380.400 705.450 381.450 ;
        RECT 700.950 379.950 703.050 380.400 ;
        RECT 709.950 379.950 712.050 382.050 ;
        RECT 676.950 346.950 679.050 349.050 ;
        RECT 709.950 346.950 712.050 349.050 ;
        RECT 677.400 346.050 678.450 346.950 ;
        RECT 676.950 343.950 679.050 346.050 ;
        RECT 680.250 344.250 681.750 345.150 ;
        RECT 682.950 343.950 685.050 346.050 ;
        RECT 670.950 340.950 673.050 343.050 ;
        RECT 676.950 341.850 678.750 342.750 ;
        RECT 679.950 340.950 682.050 343.050 ;
        RECT 683.250 341.850 685.050 342.750 ;
        RECT 710.400 342.450 711.450 346.950 ;
        RECT 712.950 342.450 715.050 343.050 ;
        RECT 710.400 341.400 715.050 342.450 ;
        RECT 694.950 337.950 697.050 340.050 ;
        RECT 695.400 316.050 696.450 337.950 ;
        RECT 643.950 313.950 646.050 316.050 ;
        RECT 652.950 313.950 655.050 316.050 ;
        RECT 694.950 313.950 697.050 316.050 ;
        RECT 649.950 311.250 652.050 312.150 ;
        RECT 652.950 311.850 655.050 312.750 ;
        RECT 658.950 312.450 661.050 313.050 ;
        RECT 691.950 312.450 694.050 313.050 ;
        RECT 655.950 311.250 657.750 312.150 ;
        RECT 658.950 311.400 663.450 312.450 ;
        RECT 658.950 310.950 661.050 311.400 ;
        RECT 640.950 307.950 643.050 310.050 ;
        RECT 649.950 307.950 652.050 310.050 ;
        RECT 655.950 307.950 658.050 310.050 ;
        RECT 659.250 308.850 661.050 309.750 ;
        RECT 650.400 307.050 651.450 307.950 ;
        RECT 613.950 304.950 616.050 305.400 ;
        RECT 619.950 305.400 624.450 306.450 ;
        RECT 619.950 304.950 622.050 305.400 ;
        RECT 649.950 304.950 652.050 307.050 ;
        RECT 619.950 301.950 622.050 304.050 ;
        RECT 601.950 271.950 604.050 274.050 ;
        RECT 610.950 271.950 613.050 274.050 ;
        RECT 616.950 273.450 619.050 274.050 ;
        RECT 620.400 273.450 621.450 301.950 ;
        RECT 614.250 272.250 615.750 273.150 ;
        RECT 616.950 272.400 621.450 273.450 ;
        RECT 616.950 271.950 619.050 272.400 ;
        RECT 662.400 271.050 663.450 311.400 ;
        RECT 689.400 311.400 694.050 312.450 ;
        RECT 695.250 311.850 696.750 312.750 ;
        RECT 689.400 304.050 690.450 311.400 ;
        RECT 691.950 310.950 694.050 311.400 ;
        RECT 691.950 308.850 694.050 309.750 ;
        RECT 697.950 308.850 700.050 309.750 ;
        RECT 688.950 301.950 691.050 304.050 ;
        RECT 610.950 269.850 612.750 270.750 ;
        RECT 613.950 268.950 616.050 271.050 ;
        RECT 617.250 269.850 619.050 270.750 ;
        RECT 637.950 268.950 640.050 271.050 ;
        RECT 652.950 269.250 654.750 270.150 ;
        RECT 655.950 268.950 658.050 271.050 ;
        RECT 661.950 270.450 664.050 271.050 ;
        RECT 661.950 269.400 666.450 270.450 ;
        RECT 661.950 268.950 664.050 269.400 ;
        RECT 614.400 253.050 615.450 268.950 ;
        RECT 613.950 250.950 616.050 253.050 ;
        RECT 613.950 247.950 616.050 250.050 ;
        RECT 614.400 241.050 615.450 247.950 ;
        RECT 619.950 241.950 622.050 244.050 ;
        RECT 613.950 238.950 616.050 241.050 ;
        RECT 617.250 239.250 619.050 240.150 ;
        RECT 619.950 239.850 622.050 240.750 ;
        RECT 622.950 239.250 625.050 240.150 ;
        RECT 613.950 236.850 615.750 237.750 ;
        RECT 616.950 235.950 619.050 238.050 ;
        RECT 622.950 235.950 625.050 238.050 ;
        RECT 610.950 198.450 613.050 199.050 ;
        RECT 610.950 197.400 615.450 198.450 ;
        RECT 610.950 196.950 613.050 197.400 ;
        RECT 607.950 194.250 610.050 195.150 ;
        RECT 610.950 194.850 613.050 195.750 ;
        RECT 607.950 190.950 610.050 193.050 ;
        RECT 601.950 187.950 604.050 190.050 ;
        RECT 602.400 169.050 603.450 187.950 ;
        RECT 614.400 175.050 615.450 197.400 ;
        RECT 617.400 196.050 618.450 235.950 ;
        RECT 616.950 193.950 619.050 196.050 ;
        RECT 622.950 190.950 625.050 193.050 ;
        RECT 613.950 172.950 616.050 175.050 ;
        RECT 607.950 169.950 610.050 172.050 ;
        RECT 601.950 166.950 604.050 169.050 ;
        RECT 605.250 167.250 607.050 168.150 ;
        RECT 607.950 167.850 610.050 168.750 ;
        RECT 610.950 167.250 613.050 168.150 ;
        RECT 601.950 164.850 603.750 165.750 ;
        RECT 604.950 163.950 607.050 166.050 ;
        RECT 610.950 163.950 613.050 166.050 ;
        RECT 610.950 157.950 613.050 160.050 ;
        RECT 611.400 130.050 612.450 157.950 ;
        RECT 616.950 131.250 619.050 132.150 ;
        RECT 610.950 127.950 613.050 130.050 ;
        RECT 614.250 128.250 615.750 129.150 ;
        RECT 616.950 127.950 619.050 130.050 ;
        RECT 620.250 128.250 622.050 129.150 ;
        RECT 610.950 125.850 612.750 126.750 ;
        RECT 613.950 124.950 616.050 127.050 ;
        RECT 614.400 124.050 615.450 124.950 ;
        RECT 613.950 121.950 616.050 124.050 ;
        RECT 607.950 115.950 610.050 118.050 ;
        RECT 604.950 94.950 607.050 97.050 ;
        RECT 595.950 88.950 598.050 91.050 ;
        RECT 556.950 82.500 559.050 84.600 ;
        RECT 578.250 83.700 579.450 87.300 ;
        RECT 580.950 85.950 583.050 88.050 ;
        RECT 577.950 81.600 580.050 83.700 ;
        RECT 541.950 56.250 544.050 57.150 ;
        RECT 547.950 55.950 550.050 58.050 ;
        RECT 548.400 55.050 549.450 55.950 ;
        RECT 541.950 52.950 544.050 55.050 ;
        RECT 545.250 53.250 546.750 54.150 ;
        RECT 547.950 52.950 550.050 55.050 ;
        RECT 551.250 53.250 553.050 54.150 ;
        RECT 583.950 53.250 586.050 54.150 ;
        RECT 589.950 52.950 592.050 55.050 ;
        RECT 499.950 49.950 502.050 52.050 ;
        RECT 505.950 49.950 508.050 52.050 ;
        RECT 538.950 49.950 541.050 52.050 ;
        RECT 430.950 46.950 433.050 49.050 ;
        RECT 457.950 46.950 460.050 49.050 ;
        RECT 478.950 46.950 481.050 49.050 ;
        RECT 481.950 46.950 484.050 49.050 ;
        RECT 424.950 31.950 427.050 34.050 ;
        RECT 460.950 31.950 463.050 34.050 ;
        RECT 425.400 25.050 426.450 31.950 ;
        RECT 427.950 25.950 430.050 28.050 ;
        RECT 337.950 22.950 340.050 25.050 ;
        RECT 340.950 22.950 343.050 25.050 ;
        RECT 344.250 23.850 345.750 24.750 ;
        RECT 346.950 22.950 349.050 25.050 ;
        RECT 349.950 22.950 352.050 25.050 ;
        RECT 361.950 22.950 364.050 25.050 ;
        RECT 379.950 22.950 382.050 25.050 ;
        RECT 383.250 23.250 384.750 24.150 ;
        RECT 385.950 22.950 388.050 25.050 ;
        RECT 388.950 22.950 391.050 25.050 ;
        RECT 424.950 22.950 427.050 25.050 ;
        RECT 428.250 23.850 429.750 24.750 ;
        RECT 430.950 22.950 433.050 25.050 ;
        RECT 350.400 22.050 351.450 22.950 ;
        RECT 389.400 22.050 390.450 22.950 ;
        RECT 316.950 19.950 319.050 22.050 ;
        RECT 340.950 20.850 343.050 21.750 ;
        RECT 346.950 20.850 349.050 21.750 ;
        RECT 349.950 19.950 352.050 22.050 ;
        RECT 379.950 20.850 381.750 21.750 ;
        RECT 382.950 19.950 385.050 22.050 ;
        RECT 386.250 20.850 387.750 21.750 ;
        RECT 388.950 19.950 391.050 22.050 ;
        RECT 424.950 20.850 427.050 21.750 ;
        RECT 430.950 20.850 433.050 21.750 ;
        RECT 262.950 15.300 265.050 17.400 ;
        RECT 313.950 16.950 316.050 19.050 ;
        RECT 388.950 17.850 391.050 18.750 ;
        RECT 461.400 18.450 462.450 31.950 ;
        RECT 482.400 25.050 483.450 46.950 ;
        RECT 508.950 28.950 511.050 31.050 ;
        RECT 505.950 25.950 508.050 28.050 ;
        RECT 509.400 25.050 510.450 28.950 ;
        RECT 535.950 25.950 538.050 28.050 ;
        RECT 542.400 27.450 543.450 52.950 ;
        RECT 544.950 49.950 547.050 52.050 ;
        RECT 548.250 50.850 549.750 51.750 ;
        RECT 550.950 49.950 553.050 52.050 ;
        RECT 580.950 50.250 582.750 51.150 ;
        RECT 583.950 49.950 586.050 52.050 ;
        RECT 589.950 50.850 592.050 51.750 ;
        RECT 545.400 34.050 546.450 49.950 ;
        RECT 605.400 49.050 606.450 94.950 ;
        RECT 580.950 46.950 583.050 49.050 ;
        RECT 604.950 46.950 607.050 49.050 ;
        RECT 544.950 31.950 547.050 34.050 ;
        RECT 608.400 28.050 609.450 115.950 ;
        RECT 617.400 103.050 618.450 127.950 ;
        RECT 619.950 124.950 622.050 127.050 ;
        RECT 620.400 118.050 621.450 124.950 ;
        RECT 623.400 124.050 624.450 190.950 ;
        RECT 638.400 163.050 639.450 268.950 ;
        RECT 652.950 265.950 655.050 268.050 ;
        RECT 656.250 266.850 658.050 267.750 ;
        RECT 658.950 266.250 661.050 267.150 ;
        RECT 661.950 266.850 664.050 267.750 ;
        RECT 653.400 244.050 654.450 265.950 ;
        RECT 658.950 262.950 661.050 265.050 ;
        RECT 659.400 262.050 660.450 262.950 ;
        RECT 658.950 259.950 661.050 262.050 ;
        RECT 661.950 259.950 664.050 262.050 ;
        RECT 652.950 241.950 655.050 244.050 ;
        RECT 662.400 241.050 663.450 259.950 ;
        RECT 665.400 244.050 666.450 269.400 ;
        RECT 691.950 269.250 694.050 270.150 ;
        RECT 697.950 269.250 700.050 270.150 ;
        RECT 691.950 265.950 694.050 268.050 ;
        RECT 695.250 266.250 696.750 267.150 ;
        RECT 692.400 261.450 693.450 265.950 ;
        RECT 694.950 262.950 697.050 265.050 ;
        RECT 697.950 262.950 700.050 265.050 ;
        RECT 692.400 260.400 696.450 261.450 ;
        RECT 679.950 256.950 682.050 259.050 ;
        RECT 664.950 241.950 667.050 244.050 ;
        RECT 655.950 239.250 658.050 240.150 ;
        RECT 661.950 238.950 664.050 241.050 ;
        RECT 665.250 239.850 667.050 240.750 ;
        RECT 655.950 235.950 658.050 238.050 ;
        RECT 661.950 236.850 664.050 237.750 ;
        RECT 649.950 199.950 652.050 202.050 ;
        RECT 640.950 197.250 643.050 198.150 ;
        RECT 646.950 197.250 649.050 198.150 ;
        RECT 640.950 193.950 643.050 196.050 ;
        RECT 646.950 195.450 649.050 196.050 ;
        RECT 650.400 195.450 651.450 199.950 ;
        RECT 644.250 194.250 645.750 195.150 ;
        RECT 646.950 194.400 651.450 195.450 ;
        RECT 680.400 195.450 681.450 256.950 ;
        RECT 695.400 247.050 696.450 260.400 ;
        RECT 694.950 244.950 697.050 247.050 ;
        RECT 695.400 241.050 696.450 244.950 ;
        RECT 685.950 238.950 688.050 241.050 ;
        RECT 694.950 238.950 697.050 241.050 ;
        RECT 686.400 202.050 687.450 238.950 ;
        RECT 694.950 236.850 697.050 237.750 ;
        RECT 691.950 202.950 694.050 205.050 ;
        RECT 685.950 199.950 688.050 202.050 ;
        RECT 686.400 199.050 687.450 199.950 ;
        RECT 692.400 199.050 693.450 202.950 ;
        RECT 682.950 197.250 684.750 198.150 ;
        RECT 685.950 196.950 688.050 199.050 ;
        RECT 691.950 196.950 694.050 199.050 ;
        RECT 698.400 196.050 699.450 262.950 ;
        RECT 710.400 262.050 711.450 341.400 ;
        RECT 712.950 340.950 715.050 341.400 ;
        RECT 718.950 340.950 721.050 343.050 ;
        RECT 722.250 341.250 724.050 342.150 ;
        RECT 728.400 340.050 729.450 382.950 ;
        RECT 733.950 379.950 736.050 382.050 ;
        RECT 730.950 340.950 733.050 343.050 ;
        RECT 757.950 342.450 760.050 343.050 ;
        RECT 755.400 341.400 760.050 342.450 ;
        RECT 712.950 338.850 715.050 339.750 ;
        RECT 715.950 338.250 718.050 339.150 ;
        RECT 718.950 338.850 720.750 339.750 ;
        RECT 721.950 337.950 724.050 340.050 ;
        RECT 727.950 337.950 730.050 340.050 ;
        RECT 715.950 334.950 718.050 337.050 ;
        RECT 727.950 312.450 730.050 313.050 ;
        RECT 725.400 311.400 730.050 312.450 ;
        RECT 725.400 304.050 726.450 311.400 ;
        RECT 727.950 310.950 730.050 311.400 ;
        RECT 727.950 308.850 730.050 309.750 ;
        RECT 731.400 306.450 732.450 340.950 ;
        RECT 736.950 334.950 739.050 337.050 ;
        RECT 737.400 313.050 738.450 334.950 ;
        RECT 736.950 310.950 739.050 313.050 ;
        RECT 733.950 308.250 736.050 309.150 ;
        RECT 736.950 308.850 739.050 309.750 ;
        RECT 728.400 305.400 732.450 306.450 ;
        RECT 724.950 301.950 727.050 304.050 ;
        RECT 728.400 267.450 729.450 305.400 ;
        RECT 730.950 269.250 733.050 270.150 ;
        RECT 736.950 269.250 739.050 270.150 ;
        RECT 730.950 267.450 733.050 268.050 ;
        RECT 728.400 266.400 733.050 267.450 ;
        RECT 736.950 267.450 739.050 268.050 ;
        RECT 730.950 265.950 733.050 266.400 ;
        RECT 734.250 266.250 735.750 267.150 ;
        RECT 736.950 266.400 741.450 267.450 ;
        RECT 736.950 265.950 739.050 266.400 ;
        RECT 709.950 259.950 712.050 262.050 ;
        RECT 703.950 238.950 706.050 241.050 ;
        RECT 724.950 238.950 727.050 241.050 ;
        RECT 700.950 236.250 703.050 237.150 ;
        RECT 703.950 236.850 706.050 237.750 ;
        RECT 725.400 199.050 726.450 238.950 ;
        RECT 731.400 202.050 732.450 265.950 ;
        RECT 733.950 262.950 736.050 265.050 ;
        RECT 734.400 262.050 735.450 262.950 ;
        RECT 733.950 259.950 736.050 262.050 ;
        RECT 740.400 244.050 741.450 266.400 ;
        RECT 739.950 241.950 742.050 244.050 ;
        RECT 736.950 238.950 739.050 241.050 ;
        RECT 740.250 239.850 741.750 240.750 ;
        RECT 736.950 236.850 739.050 237.750 ;
        RECT 742.950 236.850 745.050 237.750 ;
        RECT 755.400 205.050 756.450 341.400 ;
        RECT 757.950 340.950 760.050 341.400 ;
        RECT 757.950 338.850 760.050 339.750 ;
        RECT 760.950 338.250 763.050 339.150 ;
        RECT 760.950 334.950 763.050 337.050 ;
        RECT 761.400 265.050 762.450 334.950 ;
        RECT 760.950 262.950 763.050 265.050 ;
        RECT 754.950 202.950 757.050 205.050 ;
        RECT 730.950 199.950 733.050 202.050 ;
        RECT 721.950 197.250 724.050 198.150 ;
        RECT 724.950 196.950 727.050 199.050 ;
        RECT 727.950 197.850 730.050 198.750 ;
        RECT 730.950 197.250 733.050 198.150 ;
        RECT 682.950 195.450 685.050 196.050 ;
        RECT 680.400 194.400 685.050 195.450 ;
        RECT 686.250 194.850 688.050 195.750 ;
        RECT 646.950 193.950 649.050 194.400 ;
        RECT 682.950 193.950 685.050 194.400 ;
        RECT 688.950 194.250 691.050 195.150 ;
        RECT 691.950 194.850 694.050 195.750 ;
        RECT 697.950 193.950 700.050 196.050 ;
        RECT 721.950 195.450 724.050 196.050 ;
        RECT 725.400 195.450 726.450 196.950 ;
        RECT 721.950 194.400 726.450 195.450 ;
        RECT 721.950 193.950 724.050 194.400 ;
        RECT 730.950 193.950 733.050 196.050 ;
        RECT 643.950 190.950 646.050 193.050 ;
        RECT 688.950 190.950 691.050 193.050 ;
        RECT 721.950 190.950 724.050 193.050 ;
        RECT 733.950 190.950 736.050 193.050 ;
        RECT 649.950 172.950 652.050 175.050 ;
        RECT 685.950 172.950 688.050 175.050 ;
        RECT 650.400 172.050 651.450 172.950 ;
        RECT 643.950 169.950 646.050 172.050 ;
        RECT 649.950 169.950 652.050 172.050 ;
        RECT 682.950 171.450 685.050 172.050 ;
        RECT 680.400 170.400 685.050 171.450 ;
        RECT 644.400 169.050 645.450 169.950 ;
        RECT 643.950 166.950 646.050 169.050 ;
        RECT 647.250 167.250 649.050 168.150 ;
        RECT 649.950 167.850 652.050 168.750 ;
        RECT 652.950 167.250 655.050 168.150 ;
        RECT 680.400 166.050 681.450 170.400 ;
        RECT 682.950 169.950 685.050 170.400 ;
        RECT 686.400 169.050 687.450 172.950 ;
        RECT 682.950 167.850 684.750 168.750 ;
        RECT 685.950 166.950 688.050 169.050 ;
        RECT 691.950 167.250 694.050 168.150 ;
        RECT 643.950 164.850 645.750 165.750 ;
        RECT 646.950 163.950 649.050 166.050 ;
        RECT 652.950 163.950 655.050 166.050 ;
        RECT 679.950 163.950 682.050 166.050 ;
        RECT 685.950 164.850 688.050 165.750 ;
        RECT 691.950 163.950 694.050 166.050 ;
        RECT 647.400 163.050 648.450 163.950 ;
        RECT 637.950 160.950 640.050 163.050 ;
        RECT 646.950 160.950 649.050 163.050 ;
        RECT 649.950 130.950 652.050 133.050 ;
        RECT 650.400 130.050 651.450 130.950 ;
        RECT 649.950 127.950 652.050 130.050 ;
        RECT 653.250 128.250 654.750 129.150 ;
        RECT 655.950 127.950 658.050 130.050 ;
        RECT 664.950 127.950 667.050 130.050 ;
        RECT 649.950 125.850 651.750 126.750 ;
        RECT 652.950 124.950 655.050 127.050 ;
        RECT 656.250 125.850 658.050 126.750 ;
        RECT 622.950 121.950 625.050 124.050 ;
        RECT 655.950 121.950 658.050 124.050 ;
        RECT 619.950 115.950 622.050 118.050 ;
        RECT 616.950 100.950 619.050 103.050 ;
        RECT 652.950 100.950 655.050 103.050 ;
        RECT 616.950 97.950 619.050 100.050 ;
        RECT 613.950 96.450 616.050 97.050 ;
        RECT 611.400 95.400 616.050 96.450 ;
        RECT 617.250 95.850 618.750 96.750 ;
        RECT 611.400 52.050 612.450 95.400 ;
        RECT 613.950 94.950 616.050 95.400 ;
        RECT 619.950 94.950 622.050 97.050 ;
        RECT 653.400 94.050 654.450 100.950 ;
        RECT 613.950 92.850 616.050 93.750 ;
        RECT 619.950 92.850 622.050 93.750 ;
        RECT 652.950 91.950 655.050 94.050 ;
        RECT 656.400 91.050 657.450 121.950 ;
        RECT 658.950 97.950 661.050 100.050 ;
        RECT 659.400 94.050 660.450 97.950 ;
        RECT 665.400 94.050 666.450 127.950 ;
        RECT 680.400 127.050 681.450 163.950 ;
        RECT 692.400 163.050 693.450 163.950 ;
        RECT 691.950 160.950 694.050 163.050 ;
        RECT 694.950 130.950 697.050 133.050 ;
        RECT 695.400 130.050 696.450 130.950 ;
        RECT 688.950 127.950 691.050 130.050 ;
        RECT 694.950 129.450 697.050 130.050 ;
        RECT 692.250 128.250 693.750 129.150 ;
        RECT 694.950 128.400 699.450 129.450 ;
        RECT 694.950 127.950 697.050 128.400 ;
        RECT 679.950 124.950 682.050 127.050 ;
        RECT 688.950 125.850 690.750 126.750 ;
        RECT 691.950 124.950 694.050 127.050 ;
        RECT 695.250 125.850 697.050 126.750 ;
        RECT 698.400 123.450 699.450 128.400 ;
        RECT 695.400 122.400 699.450 123.450 ;
        RECT 658.950 91.950 661.050 94.050 ;
        RECT 662.250 92.250 664.050 93.150 ;
        RECT 664.950 91.950 667.050 94.050 ;
        RECT 652.950 89.850 654.750 90.750 ;
        RECT 655.950 88.950 658.050 91.050 ;
        RECT 659.250 89.850 660.750 90.750 ;
        RECT 661.950 88.950 664.050 91.050 ;
        RECT 655.950 86.850 658.050 87.750 ;
        RECT 658.950 55.950 661.050 58.050 ;
        RECT 664.950 56.250 667.050 57.150 ;
        RECT 659.400 55.050 660.450 55.950 ;
        RECT 695.400 55.050 696.450 122.400 ;
        RECT 703.950 100.950 706.050 103.050 ;
        RECT 709.950 100.950 712.050 103.050 ;
        RECT 700.950 97.950 703.050 100.050 ;
        RECT 697.950 95.250 700.050 96.150 ;
        RECT 697.950 91.950 700.050 94.050 ;
        RECT 701.400 58.050 702.450 97.950 ;
        RECT 704.400 97.050 705.450 100.950 ;
        RECT 706.950 97.950 709.050 100.050 ;
        RECT 703.950 94.950 706.050 97.050 ;
        RECT 707.250 95.850 709.050 96.750 ;
        RECT 703.950 92.850 706.050 93.750 ;
        RECT 700.950 57.450 703.050 58.050 ;
        RECT 698.400 56.400 703.050 57.450 ;
        RECT 706.950 57.450 709.050 58.050 ;
        RECT 710.400 57.450 711.450 100.950 ;
        RECT 722.400 97.050 723.450 190.950 ;
        RECT 734.400 169.050 735.450 190.950 ;
        RECT 724.950 168.450 727.050 169.050 ;
        RECT 724.950 167.400 729.450 168.450 ;
        RECT 724.950 166.950 727.050 167.400 ;
        RECT 724.950 164.850 727.050 165.750 ;
        RECT 728.400 130.050 729.450 167.400 ;
        RECT 733.950 166.950 736.050 169.050 ;
        RECT 730.950 164.250 733.050 165.150 ;
        RECT 733.950 164.850 736.050 165.750 ;
        RECT 727.950 129.450 730.050 130.050 ;
        RECT 725.400 128.400 730.050 129.450 ;
        RECT 721.950 94.950 724.050 97.050 ;
        RECT 725.400 88.050 726.450 128.400 ;
        RECT 727.950 127.950 730.050 128.400 ;
        RECT 731.250 128.250 732.750 129.150 ;
        RECT 727.950 125.850 729.750 126.750 ;
        RECT 730.950 124.950 733.050 127.050 ;
        RECT 734.250 125.850 736.050 126.750 ;
        RECT 739.950 100.950 742.050 103.050 ;
        RECT 740.400 100.050 741.450 100.950 ;
        RECT 739.950 97.950 742.050 100.050 ;
        RECT 736.950 94.950 739.050 97.050 ;
        RECT 740.250 95.850 741.750 96.750 ;
        RECT 742.950 96.450 745.050 97.050 ;
        RECT 742.950 95.400 747.450 96.450 ;
        RECT 742.950 94.950 745.050 95.400 ;
        RECT 736.950 92.850 739.050 93.750 ;
        RECT 742.950 92.850 745.050 93.750 ;
        RECT 724.950 85.950 727.050 88.050 ;
        RECT 622.950 52.950 625.050 55.050 ;
        RECT 655.950 53.250 657.750 54.150 ;
        RECT 658.950 52.950 661.050 55.050 ;
        RECT 662.250 53.250 663.750 54.150 ;
        RECT 664.950 52.950 667.050 55.050 ;
        RECT 694.950 52.950 697.050 55.050 ;
        RECT 698.400 52.050 699.450 56.400 ;
        RECT 700.950 55.950 703.050 56.400 ;
        RECT 704.250 56.250 705.750 57.150 ;
        RECT 706.950 56.400 711.450 57.450 ;
        RECT 706.950 55.950 709.050 56.400 ;
        RECT 700.950 53.850 702.750 54.750 ;
        RECT 703.950 52.950 706.050 55.050 ;
        RECT 707.250 53.850 709.050 54.750 ;
        RECT 725.400 52.050 726.450 85.950 ;
        RECT 736.950 53.250 739.050 54.150 ;
        RECT 742.950 53.250 745.050 54.150 ;
        RECT 610.950 49.950 613.050 52.050 ;
        RECT 622.950 50.850 625.050 51.750 ;
        RECT 625.950 50.250 628.050 51.150 ;
        RECT 655.950 49.950 658.050 52.050 ;
        RECT 659.250 50.850 660.750 51.750 ;
        RECT 661.950 49.950 664.050 52.050 ;
        RECT 697.950 49.950 700.050 52.050 ;
        RECT 724.950 49.950 727.050 52.050 ;
        RECT 733.950 51.450 736.050 52.050 ;
        RECT 736.950 51.450 739.050 52.050 ;
        RECT 733.950 50.400 739.050 51.450 ;
        RECT 733.950 49.950 736.050 50.400 ;
        RECT 736.950 49.950 739.050 50.400 ;
        RECT 740.250 50.250 741.750 51.150 ;
        RECT 746.400 49.050 747.450 95.400 ;
        RECT 622.950 46.950 625.050 49.050 ;
        RECT 625.950 46.950 628.050 49.050 ;
        RECT 739.950 46.950 742.050 49.050 ;
        RECT 745.950 46.950 748.050 49.050 ;
        RECT 539.400 26.400 543.450 27.450 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 506.250 23.850 507.750 24.750 ;
        RECT 508.950 24.450 511.050 25.050 ;
        RECT 508.950 23.400 513.450 24.450 ;
        RECT 508.950 22.950 511.050 23.400 ;
        RECT 463.950 20.250 465.750 21.150 ;
        RECT 466.950 19.950 469.050 22.050 ;
        RECT 470.250 20.250 472.050 21.150 ;
        RECT 482.400 19.050 483.450 22.950 ;
        RECT 502.950 20.850 505.050 21.750 ;
        RECT 508.950 20.850 511.050 21.750 ;
        RECT 512.400 19.050 513.450 23.400 ;
        RECT 536.400 22.050 537.450 25.950 ;
        RECT 539.400 25.050 540.450 26.400 ;
        RECT 544.950 25.950 547.050 28.050 ;
        RECT 607.950 25.950 610.050 28.050 ;
        RECT 545.400 25.050 546.450 25.950 ;
        RECT 538.950 22.950 541.050 25.050 ;
        RECT 542.250 23.250 543.750 24.150 ;
        RECT 544.950 22.950 547.050 25.050 ;
        RECT 623.400 22.050 624.450 46.950 ;
        RECT 626.400 28.050 627.450 46.950 ;
        RECT 625.950 25.950 628.050 28.050 ;
        RECT 637.950 25.950 640.050 28.050 ;
        RECT 730.950 25.950 733.050 28.050 ;
        RECT 535.950 19.950 538.050 22.050 ;
        RECT 538.950 20.850 540.750 21.750 ;
        RECT 541.950 19.950 544.050 22.050 ;
        RECT 545.250 20.850 546.750 21.750 ;
        RECT 547.950 19.950 550.050 22.050 ;
        RECT 583.950 20.250 585.750 21.150 ;
        RECT 586.950 19.950 589.050 22.050 ;
        RECT 590.250 20.250 592.050 21.150 ;
        RECT 616.950 19.950 619.050 22.050 ;
        RECT 619.950 20.250 621.750 21.150 ;
        RECT 622.950 19.950 625.050 22.050 ;
        RECT 626.250 20.250 628.050 21.150 ;
        RECT 628.950 19.950 631.050 22.050 ;
        RECT 463.950 18.450 466.050 19.050 ;
        RECT 461.400 17.400 466.050 18.450 ;
        RECT 467.250 17.850 468.750 18.750 ;
        RECT 463.950 16.950 466.050 17.400 ;
        RECT 469.950 16.950 472.050 19.050 ;
        RECT 481.950 16.950 484.050 19.050 ;
        RECT 511.950 16.950 514.050 19.050 ;
        RECT 547.950 17.850 550.050 18.750 ;
        RECT 587.250 17.850 588.750 18.750 ;
        RECT 589.950 16.950 592.050 19.050 ;
        RECT 617.400 18.450 618.450 19.950 ;
        RECT 619.950 18.450 622.050 19.050 ;
        RECT 617.400 17.400 622.050 18.450 ;
        RECT 623.250 17.850 624.750 18.750 ;
        RECT 625.950 18.450 628.050 19.050 ;
        RECT 629.400 18.450 630.450 19.950 ;
        RECT 638.400 19.050 639.450 25.950 ;
        RECT 658.950 23.850 661.050 24.750 ;
        RECT 661.950 23.250 664.050 24.150 ;
        RECT 730.950 23.850 733.050 24.750 ;
        RECT 733.950 23.250 736.050 24.150 ;
        RECT 661.950 19.950 664.050 22.050 ;
        RECT 694.950 20.250 696.750 21.150 ;
        RECT 697.950 19.950 700.050 22.050 ;
        RECT 701.250 20.250 703.050 21.150 ;
        RECT 733.950 19.950 736.050 22.050 ;
        RECT 662.400 19.050 663.450 19.950 ;
        RECT 734.400 19.050 735.450 19.950 ;
        RECT 619.950 16.950 622.050 17.400 ;
        RECT 625.950 17.400 630.450 18.450 ;
        RECT 625.950 16.950 628.050 17.400 ;
        RECT 637.950 16.950 640.050 19.050 ;
        RECT 661.950 16.950 664.050 19.050 ;
        RECT 694.950 16.950 697.050 19.050 ;
        RECT 698.250 17.850 699.750 18.750 ;
        RECT 700.950 16.950 703.050 19.050 ;
        RECT 733.950 16.950 736.050 19.050 ;
        RECT 205.950 9.600 208.050 11.700 ;
        RECT 226.950 10.500 229.050 12.600 ;
        RECT 241.950 10.500 244.050 12.600 ;
        RECT 263.250 11.700 264.450 15.300 ;
        RECT 262.950 9.600 265.050 11.700 ;
      LAYER metal3 ;
        RECT 112.950 705.600 115.050 706.050 ;
        RECT 151.950 705.600 154.050 706.050 ;
        RECT 112.950 704.400 154.050 705.600 ;
        RECT 112.950 703.950 115.050 704.400 ;
        RECT 151.950 703.950 154.050 704.400 ;
        RECT 610.950 705.600 613.050 706.050 ;
        RECT 616.950 705.600 619.050 706.050 ;
        RECT 610.950 704.400 619.050 705.600 ;
        RECT 610.950 703.950 613.050 704.400 ;
        RECT 616.950 703.950 619.050 704.400 ;
        RECT 64.950 702.600 67.050 703.050 ;
        RECT 76.950 702.600 79.050 703.050 ;
        RECT 64.950 701.400 79.050 702.600 ;
        RECT 64.950 700.950 67.050 701.400 ;
        RECT 76.950 700.950 79.050 701.400 ;
        RECT 187.950 702.600 190.050 703.050 ;
        RECT 199.950 702.600 202.050 703.050 ;
        RECT 229.950 702.600 232.050 703.050 ;
        RECT 187.950 701.400 198.600 702.600 ;
        RECT 187.950 700.950 190.050 701.400 ;
        RECT 73.950 699.600 76.050 700.050 ;
        RECT 142.950 699.600 145.050 700.050 ;
        RECT 73.950 698.400 145.050 699.600 ;
        RECT 73.950 697.950 76.050 698.400 ;
        RECT 142.950 697.950 145.050 698.400 ;
        RECT 148.950 699.600 151.050 700.050 ;
        RECT 197.400 699.600 198.600 701.400 ;
        RECT 199.950 701.400 232.050 702.600 ;
        RECT 199.950 700.950 202.050 701.400 ;
        RECT 229.950 700.950 232.050 701.400 ;
        RECT 262.950 702.600 265.050 703.050 ;
        RECT 268.950 702.600 271.050 703.050 ;
        RECT 262.950 701.400 271.050 702.600 ;
        RECT 262.950 700.950 265.050 701.400 ;
        RECT 268.950 700.950 271.050 701.400 ;
        RECT 505.950 702.600 508.050 703.050 ;
        RECT 535.950 702.600 538.050 703.050 ;
        RECT 541.950 702.600 544.050 703.050 ;
        RECT 505.950 701.400 544.050 702.600 ;
        RECT 505.950 700.950 508.050 701.400 ;
        RECT 535.950 700.950 538.050 701.400 ;
        RECT 541.950 700.950 544.050 701.400 ;
        RECT 547.950 700.950 550.050 703.050 ;
        RECT 739.950 702.600 742.050 703.050 ;
        RECT 748.950 702.600 751.050 703.050 ;
        RECT 739.950 701.400 751.050 702.600 ;
        RECT 739.950 700.950 742.050 701.400 ;
        RECT 748.950 700.950 751.050 701.400 ;
        RECT 214.950 699.600 217.050 700.050 ;
        RECT 148.950 698.400 195.600 699.600 ;
        RECT 197.400 698.400 217.050 699.600 ;
        RECT 148.950 697.950 151.050 698.400 ;
        RECT 194.400 697.050 195.600 698.400 ;
        RECT 214.950 697.950 217.050 698.400 ;
        RECT 265.950 699.600 268.050 700.050 ;
        RECT 343.950 699.600 346.050 700.050 ;
        RECT 385.950 699.600 388.050 700.050 ;
        RECT 265.950 698.400 388.050 699.600 ;
        RECT 265.950 697.950 268.050 698.400 ;
        RECT 343.950 697.950 346.050 698.400 ;
        RECT 385.950 697.950 388.050 698.400 ;
        RECT 418.950 699.600 421.050 700.050 ;
        RECT 424.950 699.600 427.050 700.050 ;
        RECT 418.950 698.400 427.050 699.600 ;
        RECT 548.400 699.600 549.600 700.950 ;
        RECT 548.400 698.400 585.600 699.600 ;
        RECT 418.950 697.950 421.050 698.400 ;
        RECT 424.950 697.950 427.050 698.400 ;
        RECT 584.400 697.050 585.600 698.400 ;
        RECT 34.950 696.600 37.050 697.050 ;
        RECT 73.950 696.600 76.050 697.050 ;
        RECT 79.950 696.600 82.050 697.050 ;
        RECT 34.950 695.400 82.050 696.600 ;
        RECT 34.950 694.950 37.050 695.400 ;
        RECT 73.950 694.950 76.050 695.400 ;
        RECT 79.950 694.950 82.050 695.400 ;
        RECT 193.950 694.950 196.050 697.050 ;
        RECT 214.950 696.600 217.050 697.050 ;
        RECT 226.950 696.600 229.050 697.050 ;
        RECT 262.950 696.600 265.050 697.050 ;
        RECT 304.950 696.600 307.050 697.050 ;
        RECT 214.950 695.400 307.050 696.600 ;
        RECT 214.950 694.950 217.050 695.400 ;
        RECT 226.950 694.950 229.050 695.400 ;
        RECT 262.950 694.950 265.050 695.400 ;
        RECT 304.950 694.950 307.050 695.400 ;
        RECT 475.950 696.600 478.050 697.050 ;
        RECT 499.950 696.600 502.050 697.050 ;
        RECT 532.950 696.600 535.050 697.050 ;
        RECT 580.950 696.600 583.050 697.050 ;
        RECT 475.950 695.400 583.050 696.600 ;
        RECT 475.950 694.950 478.050 695.400 ;
        RECT 499.950 694.950 502.050 695.400 ;
        RECT 532.950 694.950 535.050 695.400 ;
        RECT 580.950 694.950 583.050 695.400 ;
        RECT 583.950 694.950 586.050 697.050 ;
        RECT 658.950 696.600 661.050 697.050 ;
        RECT 664.950 696.600 667.050 697.050 ;
        RECT 658.950 695.400 667.050 696.600 ;
        RECT 658.950 694.950 661.050 695.400 ;
        RECT 664.950 694.950 667.050 695.400 ;
        RECT 688.950 696.600 691.050 697.050 ;
        RECT 727.950 696.600 730.050 697.050 ;
        RECT 688.950 695.400 730.050 696.600 ;
        RECT 688.950 694.950 691.050 695.400 ;
        RECT 727.950 694.950 730.050 695.400 ;
        RECT 37.950 693.600 40.050 694.050 ;
        RECT 184.950 693.600 187.050 694.050 ;
        RECT 235.950 693.600 238.050 694.050 ;
        RECT 37.950 692.400 238.050 693.600 ;
        RECT 37.950 691.950 40.050 692.400 ;
        RECT 184.950 691.950 187.050 692.400 ;
        RECT 235.950 691.950 238.050 692.400 ;
        RECT 202.950 690.600 205.050 691.050 ;
        RECT 229.950 690.600 232.050 691.050 ;
        RECT 274.950 690.600 277.050 691.050 ;
        RECT 202.950 689.400 277.050 690.600 ;
        RECT 202.950 688.950 205.050 689.400 ;
        RECT 229.950 688.950 232.050 689.400 ;
        RECT 274.950 688.950 277.050 689.400 ;
        RECT 550.950 684.600 553.050 685.050 ;
        RECT 586.950 684.600 589.050 685.050 ;
        RECT 550.950 683.400 589.050 684.600 ;
        RECT 550.950 682.950 553.050 683.400 ;
        RECT 586.950 682.950 589.050 683.400 ;
        RECT 70.950 681.600 73.050 682.050 ;
        RECT 103.950 681.600 106.050 682.050 ;
        RECT 70.950 680.400 106.050 681.600 ;
        RECT 70.950 679.950 73.050 680.400 ;
        RECT 103.950 679.950 106.050 680.400 ;
        RECT 469.950 681.600 472.050 682.050 ;
        RECT 505.950 681.600 508.050 682.050 ;
        RECT 469.950 680.400 508.050 681.600 ;
        RECT 469.950 679.950 472.050 680.400 ;
        RECT 505.950 679.950 508.050 680.400 ;
        RECT 442.950 678.600 445.050 679.050 ;
        RECT 544.950 678.600 547.050 679.050 ;
        RECT 442.950 677.400 547.050 678.600 ;
        RECT 442.950 676.950 445.050 677.400 ;
        RECT 544.950 676.950 547.050 677.400 ;
        RECT 64.950 675.600 67.050 676.050 ;
        RECT 76.950 675.600 79.050 676.050 ;
        RECT 64.950 674.400 79.050 675.600 ;
        RECT 64.950 673.950 67.050 674.400 ;
        RECT 76.950 673.950 79.050 674.400 ;
        RECT 103.950 675.600 106.050 676.050 ;
        RECT 112.950 675.600 115.050 676.050 ;
        RECT 103.950 674.400 115.050 675.600 ;
        RECT 103.950 673.950 106.050 674.400 ;
        RECT 112.950 673.950 115.050 674.400 ;
        RECT 187.950 675.600 190.050 676.050 ;
        RECT 193.950 675.600 196.050 676.050 ;
        RECT 187.950 674.400 196.050 675.600 ;
        RECT 187.950 673.950 190.050 674.400 ;
        RECT 193.950 673.950 196.050 674.400 ;
        RECT 208.950 675.600 211.050 676.050 ;
        RECT 250.950 675.600 253.050 676.050 ;
        RECT 286.950 675.600 289.050 676.050 ;
        RECT 208.950 674.400 289.050 675.600 ;
        RECT 208.950 673.950 211.050 674.400 ;
        RECT 250.950 673.950 253.050 674.400 ;
        RECT 286.950 673.950 289.050 674.400 ;
        RECT 304.950 675.600 307.050 676.050 ;
        RECT 343.950 675.600 346.050 676.050 ;
        RECT 304.950 674.400 346.050 675.600 ;
        RECT 304.950 673.950 307.050 674.400 ;
        RECT 343.950 673.950 346.050 674.400 ;
        RECT 352.950 675.600 355.050 676.050 ;
        RECT 370.950 675.600 373.050 676.050 ;
        RECT 427.950 675.600 430.050 676.050 ;
        RECT 469.950 675.600 472.050 676.050 ;
        RECT 352.950 674.400 472.050 675.600 ;
        RECT 352.950 673.950 355.050 674.400 ;
        RECT 370.950 673.950 373.050 674.400 ;
        RECT 427.950 673.950 430.050 674.400 ;
        RECT 469.950 673.950 472.050 674.400 ;
        RECT 475.950 675.600 478.050 676.050 ;
        RECT 502.950 675.600 505.050 676.050 ;
        RECT 475.950 674.400 505.050 675.600 ;
        RECT 475.950 673.950 478.050 674.400 ;
        RECT 502.950 673.950 505.050 674.400 ;
        RECT 610.950 675.600 613.050 676.050 ;
        RECT 697.950 675.600 700.050 676.050 ;
        RECT 610.950 674.400 700.050 675.600 ;
        RECT 610.950 673.950 613.050 674.400 ;
        RECT 697.950 673.950 700.050 674.400 ;
        RECT 106.950 670.950 109.050 673.050 ;
        RECT 136.950 672.600 139.050 673.050 ;
        RECT 181.950 672.600 184.050 673.050 ;
        RECT 226.950 672.600 229.050 673.050 ;
        RECT 136.950 671.400 184.050 672.600 ;
        RECT 136.950 670.950 139.050 671.400 ;
        RECT 181.950 670.950 184.050 671.400 ;
        RECT 185.400 671.400 229.050 672.600 ;
        RECT 31.950 669.600 34.050 670.050 ;
        RECT 40.950 669.600 43.050 670.050 ;
        RECT 31.950 668.400 43.050 669.600 ;
        RECT 31.950 667.950 34.050 668.400 ;
        RECT 40.950 667.950 43.050 668.400 ;
        RECT 67.950 669.600 70.050 670.050 ;
        RECT 107.400 669.600 108.600 670.950 ;
        RECT 185.400 670.050 186.600 671.400 ;
        RECT 226.950 670.950 229.050 671.400 ;
        RECT 232.950 672.600 235.050 673.050 ;
        RECT 256.950 672.600 259.050 673.050 ;
        RECT 232.950 671.400 259.050 672.600 ;
        RECT 232.950 670.950 235.050 671.400 ;
        RECT 256.950 670.950 259.050 671.400 ;
        RECT 265.950 672.600 268.050 673.050 ;
        RECT 274.950 672.600 277.050 673.050 ;
        RECT 265.950 671.400 277.050 672.600 ;
        RECT 265.950 670.950 268.050 671.400 ;
        RECT 274.950 670.950 277.050 671.400 ;
        RECT 292.950 672.600 295.050 673.050 ;
        RECT 337.950 672.600 340.050 673.050 ;
        RECT 292.950 671.400 340.050 672.600 ;
        RECT 292.950 670.950 295.050 671.400 ;
        RECT 337.950 670.950 340.050 671.400 ;
        RECT 388.950 672.600 391.050 673.050 ;
        RECT 421.950 672.600 424.050 673.050 ;
        RECT 388.950 671.400 424.050 672.600 ;
        RECT 388.950 670.950 391.050 671.400 ;
        RECT 421.950 670.950 424.050 671.400 ;
        RECT 466.950 672.600 469.050 673.050 ;
        RECT 499.950 672.600 502.050 673.050 ;
        RECT 466.950 671.400 502.050 672.600 ;
        RECT 466.950 670.950 469.050 671.400 ;
        RECT 499.950 670.950 502.050 671.400 ;
        RECT 550.950 672.600 553.050 673.050 ;
        RECT 583.950 672.600 586.050 673.050 ;
        RECT 550.950 671.400 586.050 672.600 ;
        RECT 550.950 670.950 553.050 671.400 ;
        RECT 583.950 670.950 586.050 671.400 ;
        RECT 613.950 672.600 616.050 673.050 ;
        RECT 622.950 672.600 625.050 673.050 ;
        RECT 613.950 671.400 625.050 672.600 ;
        RECT 613.950 670.950 616.050 671.400 ;
        RECT 622.950 670.950 625.050 671.400 ;
        RECT 664.950 672.600 667.050 673.050 ;
        RECT 670.950 672.600 673.050 673.050 ;
        RECT 664.950 671.400 673.050 672.600 ;
        RECT 664.950 670.950 667.050 671.400 ;
        RECT 670.950 670.950 673.050 671.400 ;
        RECT 67.950 668.400 108.600 669.600 ;
        RECT 67.950 667.950 70.050 668.400 ;
        RECT 184.950 667.950 187.050 670.050 ;
        RECT 193.950 669.600 196.050 670.050 ;
        RECT 223.950 669.600 226.050 670.050 ;
        RECT 193.950 668.400 226.050 669.600 ;
        RECT 193.950 667.950 196.050 668.400 ;
        RECT 223.950 667.950 226.050 668.400 ;
        RECT 229.950 669.600 232.050 670.050 ;
        RECT 238.950 669.600 241.050 670.050 ;
        RECT 229.950 668.400 241.050 669.600 ;
        RECT 229.950 667.950 232.050 668.400 ;
        RECT 238.950 667.950 241.050 668.400 ;
        RECT 271.950 669.600 274.050 670.050 ;
        RECT 340.950 669.600 343.050 670.050 ;
        RECT 271.950 668.400 343.050 669.600 ;
        RECT 271.950 667.950 274.050 668.400 ;
        RECT 340.950 667.950 343.050 668.400 ;
        RECT 346.950 669.600 349.050 670.050 ;
        RECT 382.950 669.600 385.050 670.050 ;
        RECT 346.950 668.400 385.050 669.600 ;
        RECT 346.950 667.950 349.050 668.400 ;
        RECT 382.950 667.950 385.050 668.400 ;
        RECT 391.950 669.600 394.050 670.050 ;
        RECT 424.950 669.600 427.050 670.050 ;
        RECT 467.400 669.600 468.600 670.950 ;
        RECT 391.950 668.400 468.600 669.600 ;
        RECT 502.950 669.600 505.050 670.050 ;
        RECT 541.950 669.600 544.050 670.050 ;
        RECT 502.950 668.400 544.050 669.600 ;
        RECT 391.950 667.950 394.050 668.400 ;
        RECT 424.950 667.950 427.050 668.400 ;
        RECT 502.950 667.950 505.050 668.400 ;
        RECT 541.950 667.950 544.050 668.400 ;
        RECT 586.950 669.600 589.050 670.050 ;
        RECT 616.950 669.600 619.050 670.050 ;
        RECT 586.950 668.400 619.050 669.600 ;
        RECT 586.950 667.950 589.050 668.400 ;
        RECT 616.950 667.950 619.050 668.400 ;
        RECT 628.950 669.600 631.050 670.050 ;
        RECT 706.950 669.600 709.050 670.050 ;
        RECT 628.950 668.400 709.050 669.600 ;
        RECT 628.950 667.950 631.050 668.400 ;
        RECT 706.950 667.950 709.050 668.400 ;
        RECT 709.950 669.600 712.050 670.050 ;
        RECT 742.950 669.600 745.050 670.050 ;
        RECT 709.950 668.400 745.050 669.600 ;
        RECT 709.950 667.950 712.050 668.400 ;
        RECT 742.950 667.950 745.050 668.400 ;
        RECT 187.950 666.600 190.050 667.050 ;
        RECT 214.950 666.600 217.050 667.050 ;
        RECT 187.950 665.400 217.050 666.600 ;
        RECT 187.950 664.950 190.050 665.400 ;
        RECT 214.950 664.950 217.050 665.400 ;
        RECT 463.950 666.600 466.050 667.050 ;
        RECT 544.950 666.600 547.050 667.050 ;
        RECT 463.950 665.400 547.050 666.600 ;
        RECT 463.950 664.950 466.050 665.400 ;
        RECT 544.950 664.950 547.050 665.400 ;
        RECT 658.950 666.600 661.050 667.050 ;
        RECT 667.950 666.600 670.050 667.050 ;
        RECT 658.950 665.400 670.050 666.600 ;
        RECT 658.950 664.950 661.050 665.400 ;
        RECT 667.950 664.950 670.050 665.400 ;
        RECT 694.950 666.600 697.050 667.050 ;
        RECT 739.950 666.600 742.050 667.050 ;
        RECT 694.950 665.400 742.050 666.600 ;
        RECT 694.950 664.950 697.050 665.400 ;
        RECT 739.950 664.950 742.050 665.400 ;
        RECT 94.950 663.600 97.050 664.050 ;
        RECT 133.950 663.600 136.050 664.050 ;
        RECT 208.950 663.600 211.050 664.050 ;
        RECT 94.950 662.400 211.050 663.600 ;
        RECT 94.950 661.950 97.050 662.400 ;
        RECT 133.950 661.950 136.050 662.400 ;
        RECT 208.950 661.950 211.050 662.400 ;
        RECT 649.950 663.600 652.050 664.050 ;
        RECT 661.950 663.600 664.050 664.050 ;
        RECT 649.950 662.400 664.050 663.600 ;
        RECT 649.950 661.950 652.050 662.400 ;
        RECT 661.950 661.950 664.050 662.400 ;
        RECT 388.950 654.600 391.050 655.050 ;
        RECT 460.950 654.600 463.050 655.050 ;
        RECT 388.950 653.400 463.050 654.600 ;
        RECT 388.950 652.950 391.050 653.400 ;
        RECT 460.950 652.950 463.050 653.400 ;
        RECT 31.950 651.600 34.050 652.050 ;
        RECT 64.950 651.600 67.050 652.050 ;
        RECT 31.950 650.400 67.050 651.600 ;
        RECT 31.950 649.950 34.050 650.400 ;
        RECT 64.950 649.950 67.050 650.400 ;
        RECT 298.950 651.600 301.050 652.050 ;
        RECT 379.950 651.600 382.050 652.050 ;
        RECT 298.950 650.400 382.050 651.600 ;
        RECT 298.950 649.950 301.050 650.400 ;
        RECT 379.950 649.950 382.050 650.400 ;
        RECT 145.950 642.600 148.050 643.050 ;
        RECT 190.950 642.600 193.050 643.050 ;
        RECT 145.950 641.400 193.050 642.600 ;
        RECT 145.950 640.950 148.050 641.400 ;
        RECT 190.950 640.950 193.050 641.400 ;
        RECT 232.950 633.600 235.050 634.050 ;
        RECT 265.950 633.600 268.050 634.050 ;
        RECT 232.950 632.400 268.050 633.600 ;
        RECT 232.950 631.950 235.050 632.400 ;
        RECT 265.950 631.950 268.050 632.400 ;
        RECT 418.950 631.950 421.050 634.050 ;
        RECT 535.950 633.600 538.050 634.050 ;
        RECT 544.950 633.600 547.050 634.050 ;
        RECT 535.950 632.400 547.050 633.600 ;
        RECT 535.950 631.950 538.050 632.400 ;
        RECT 544.950 631.950 547.050 632.400 ;
        RECT 574.950 633.600 577.050 634.050 ;
        RECT 613.950 633.600 616.050 634.050 ;
        RECT 619.950 633.600 622.050 634.050 ;
        RECT 574.950 632.400 622.050 633.600 ;
        RECT 574.950 631.950 577.050 632.400 ;
        RECT 613.950 631.950 616.050 632.400 ;
        RECT 619.950 631.950 622.050 632.400 ;
        RECT 181.950 630.600 184.050 631.050 ;
        RECT 193.950 630.600 196.050 631.050 ;
        RECT 181.950 629.400 196.050 630.600 ;
        RECT 181.950 628.950 184.050 629.400 ;
        RECT 193.950 628.950 196.050 629.400 ;
        RECT 211.950 630.600 214.050 631.050 ;
        RECT 226.950 630.600 229.050 631.050 ;
        RECT 211.950 629.400 229.050 630.600 ;
        RECT 211.950 628.950 214.050 629.400 ;
        RECT 226.950 628.950 229.050 629.400 ;
        RECT 307.950 630.600 310.050 631.050 ;
        RECT 343.950 630.600 346.050 631.050 ;
        RECT 415.950 630.600 418.050 631.050 ;
        RECT 307.950 629.400 418.050 630.600 ;
        RECT 307.950 628.950 310.050 629.400 ;
        RECT 343.950 628.950 346.050 629.400 ;
        RECT 415.950 628.950 418.050 629.400 ;
        RECT 76.950 627.600 79.050 628.050 ;
        RECT 103.950 627.600 106.050 628.050 ;
        RECT 112.950 627.600 115.050 628.050 ;
        RECT 76.950 626.400 115.050 627.600 ;
        RECT 76.950 625.950 79.050 626.400 ;
        RECT 103.950 625.950 106.050 626.400 ;
        RECT 112.950 625.950 115.050 626.400 ;
        RECT 220.950 627.600 223.050 628.050 ;
        RECT 238.950 627.600 241.050 628.050 ;
        RECT 220.950 626.400 241.050 627.600 ;
        RECT 220.950 625.950 223.050 626.400 ;
        RECT 238.950 625.950 241.050 626.400 ;
        RECT 301.950 627.600 304.050 628.050 ;
        RECT 346.950 627.600 349.050 628.050 ;
        RECT 385.950 627.600 388.050 628.050 ;
        RECT 301.950 626.400 388.050 627.600 ;
        RECT 301.950 625.950 304.050 626.400 ;
        RECT 346.950 625.950 349.050 626.400 ;
        RECT 385.950 625.950 388.050 626.400 ;
        RECT 34.950 624.600 37.050 625.050 ;
        RECT 40.950 624.600 43.050 625.050 ;
        RECT 67.950 624.600 70.050 625.050 ;
        RECT 34.950 623.400 70.050 624.600 ;
        RECT 34.950 622.950 37.050 623.400 ;
        RECT 40.950 622.950 43.050 623.400 ;
        RECT 67.950 622.950 70.050 623.400 ;
        RECT 118.950 624.600 121.050 625.050 ;
        RECT 142.950 624.600 145.050 625.050 ;
        RECT 118.950 623.400 145.050 624.600 ;
        RECT 419.400 624.600 420.600 631.950 ;
        RECT 421.950 630.600 424.050 631.050 ;
        RECT 442.950 630.600 445.050 631.050 ;
        RECT 472.950 630.600 475.050 631.050 ;
        RECT 421.950 629.400 475.050 630.600 ;
        RECT 421.950 628.950 424.050 629.400 ;
        RECT 442.950 628.950 445.050 629.400 ;
        RECT 472.950 628.950 475.050 629.400 ;
        RECT 493.950 630.600 496.050 631.050 ;
        RECT 499.950 630.600 502.050 631.050 ;
        RECT 493.950 629.400 502.050 630.600 ;
        RECT 493.950 628.950 496.050 629.400 ;
        RECT 499.950 628.950 502.050 629.400 ;
        RECT 511.950 630.600 514.050 631.050 ;
        RECT 550.950 630.600 553.050 631.050 ;
        RECT 511.950 629.400 553.050 630.600 ;
        RECT 511.950 628.950 514.050 629.400 ;
        RECT 550.950 628.950 553.050 629.400 ;
        RECT 652.950 630.600 655.050 631.050 ;
        RECT 658.950 630.600 661.050 631.050 ;
        RECT 652.950 629.400 661.050 630.600 ;
        RECT 652.950 628.950 655.050 629.400 ;
        RECT 658.950 628.950 661.050 629.400 ;
        RECT 664.950 630.600 667.050 631.050 ;
        RECT 670.950 630.600 673.050 631.050 ;
        RECT 664.950 629.400 673.050 630.600 ;
        RECT 664.950 628.950 667.050 629.400 ;
        RECT 670.950 628.950 673.050 629.400 ;
        RECT 688.950 630.600 691.050 631.050 ;
        RECT 697.950 630.600 700.050 631.050 ;
        RECT 688.950 629.400 700.050 630.600 ;
        RECT 688.950 628.950 691.050 629.400 ;
        RECT 697.950 628.950 700.050 629.400 ;
        RECT 460.950 627.600 463.050 628.050 ;
        RECT 502.950 627.600 505.050 628.050 ;
        RECT 460.950 626.400 505.050 627.600 ;
        RECT 460.950 625.950 463.050 626.400 ;
        RECT 502.950 625.950 505.050 626.400 ;
        RECT 649.950 627.600 652.050 628.050 ;
        RECT 655.950 627.600 658.050 628.050 ;
        RECT 649.950 626.400 658.050 627.600 ;
        RECT 649.950 625.950 652.050 626.400 ;
        RECT 655.950 625.950 658.050 626.400 ;
        RECT 427.950 624.600 430.050 625.050 ;
        RECT 419.400 623.400 430.050 624.600 ;
        RECT 118.950 622.950 121.050 623.400 ;
        RECT 142.950 622.950 145.050 623.400 ;
        RECT 427.950 622.950 430.050 623.400 ;
        RECT 430.950 624.600 433.050 625.050 ;
        RECT 586.950 624.600 589.050 625.050 ;
        RECT 613.950 624.600 616.050 625.050 ;
        RECT 430.950 623.400 616.050 624.600 ;
        RECT 430.950 622.950 433.050 623.400 ;
        RECT 586.950 622.950 589.050 623.400 ;
        RECT 613.950 622.950 616.050 623.400 ;
        RECT 700.950 624.600 703.050 625.050 ;
        RECT 727.950 624.600 730.050 625.050 ;
        RECT 700.950 623.400 730.050 624.600 ;
        RECT 700.950 622.950 703.050 623.400 ;
        RECT 727.950 622.950 730.050 623.400 ;
        RECT 415.950 621.600 418.050 622.050 ;
        RECT 424.950 621.600 427.050 622.050 ;
        RECT 463.950 621.600 466.050 622.050 ;
        RECT 415.950 620.400 466.050 621.600 ;
        RECT 415.950 619.950 418.050 620.400 ;
        RECT 424.950 619.950 427.050 620.400 ;
        RECT 463.950 619.950 466.050 620.400 ;
        RECT 505.950 621.600 508.050 622.050 ;
        RECT 547.950 621.600 550.050 622.050 ;
        RECT 505.950 620.400 550.050 621.600 ;
        RECT 505.950 619.950 508.050 620.400 ;
        RECT 547.950 619.950 550.050 620.400 ;
        RECT 466.950 618.600 469.050 619.050 ;
        RECT 574.950 618.600 577.050 619.050 ;
        RECT 466.950 617.400 577.050 618.600 ;
        RECT 466.950 616.950 469.050 617.400 ;
        RECT 574.950 616.950 577.050 617.400 ;
        RECT 262.950 606.600 265.050 607.050 ;
        RECT 304.950 606.600 307.050 607.050 ;
        RECT 337.950 606.600 340.050 607.050 ;
        RECT 262.950 605.400 340.050 606.600 ;
        RECT 262.950 604.950 265.050 605.400 ;
        RECT 304.950 604.950 307.050 605.400 ;
        RECT 337.950 604.950 340.050 605.400 ;
        RECT 340.950 606.600 343.050 607.050 ;
        RECT 346.950 606.600 349.050 607.050 ;
        RECT 340.950 605.400 349.050 606.600 ;
        RECT 340.950 604.950 343.050 605.400 ;
        RECT 346.950 604.950 349.050 605.400 ;
        RECT 499.950 606.600 502.050 607.050 ;
        RECT 541.950 606.600 544.050 607.050 ;
        RECT 499.950 605.400 544.050 606.600 ;
        RECT 499.950 604.950 502.050 605.400 ;
        RECT 541.950 604.950 544.050 605.400 ;
        RECT 598.950 606.600 601.050 607.050 ;
        RECT 661.950 606.600 664.050 607.050 ;
        RECT 598.950 605.400 664.050 606.600 ;
        RECT 598.950 604.950 601.050 605.400 ;
        RECT 661.950 604.950 664.050 605.400 ;
        RECT 34.950 603.600 37.050 604.050 ;
        RECT 49.950 603.600 52.050 604.050 ;
        RECT 34.950 602.400 52.050 603.600 ;
        RECT 34.950 601.950 37.050 602.400 ;
        RECT 49.950 601.950 52.050 602.400 ;
        RECT 55.950 603.600 58.050 604.050 ;
        RECT 94.950 603.600 97.050 604.050 ;
        RECT 55.950 602.400 97.050 603.600 ;
        RECT 55.950 601.950 58.050 602.400 ;
        RECT 94.950 601.950 97.050 602.400 ;
        RECT 109.950 603.600 112.050 604.050 ;
        RECT 139.950 603.600 142.050 604.050 ;
        RECT 109.950 602.400 142.050 603.600 ;
        RECT 109.950 601.950 112.050 602.400 ;
        RECT 139.950 601.950 142.050 602.400 ;
        RECT 160.950 603.600 163.050 604.050 ;
        RECT 181.950 603.600 184.050 604.050 ;
        RECT 211.950 603.600 214.050 604.050 ;
        RECT 160.950 602.400 214.050 603.600 ;
        RECT 160.950 601.950 163.050 602.400 ;
        RECT 181.950 601.950 184.050 602.400 ;
        RECT 211.950 601.950 214.050 602.400 ;
        RECT 259.950 603.600 262.050 604.050 ;
        RECT 334.950 603.600 337.050 604.050 ;
        RECT 259.950 602.400 337.050 603.600 ;
        RECT 259.950 601.950 262.050 602.400 ;
        RECT 334.950 601.950 337.050 602.400 ;
        RECT 340.950 603.600 343.050 604.050 ;
        RECT 376.950 603.600 379.050 604.050 ;
        RECT 340.950 602.400 379.050 603.600 ;
        RECT 340.950 601.950 343.050 602.400 ;
        RECT 376.950 601.950 379.050 602.400 ;
        RECT 577.950 603.600 580.050 604.050 ;
        RECT 619.950 603.600 622.050 604.050 ;
        RECT 577.950 602.400 622.050 603.600 ;
        RECT 577.950 601.950 580.050 602.400 ;
        RECT 619.950 601.950 622.050 602.400 ;
        RECT 718.950 603.600 721.050 604.050 ;
        RECT 727.950 603.600 730.050 604.050 ;
        RECT 718.950 602.400 730.050 603.600 ;
        RECT 718.950 601.950 721.050 602.400 ;
        RECT 727.950 601.950 730.050 602.400 ;
        RECT 37.950 600.600 40.050 601.050 ;
        RECT 43.950 600.600 46.050 601.050 ;
        RECT 37.950 599.400 46.050 600.600 ;
        RECT 37.950 598.950 40.050 599.400 ;
        RECT 43.950 598.950 46.050 599.400 ;
        RECT 61.950 600.600 64.050 601.050 ;
        RECT 79.950 600.600 82.050 601.050 ;
        RECT 61.950 599.400 82.050 600.600 ;
        RECT 61.950 598.950 64.050 599.400 ;
        RECT 79.950 598.950 82.050 599.400 ;
        RECT 88.950 600.600 91.050 601.050 ;
        RECT 175.950 600.600 178.050 601.050 ;
        RECT 88.950 599.400 178.050 600.600 ;
        RECT 88.950 598.950 91.050 599.400 ;
        RECT 175.950 598.950 178.050 599.400 ;
        RECT 199.950 600.600 202.050 601.050 ;
        RECT 253.950 600.600 256.050 601.050 ;
        RECT 199.950 599.400 256.050 600.600 ;
        RECT 199.950 598.950 202.050 599.400 ;
        RECT 253.950 598.950 256.050 599.400 ;
        RECT 382.950 600.600 385.050 601.050 ;
        RECT 412.950 600.600 415.050 601.050 ;
        RECT 382.950 599.400 415.050 600.600 ;
        RECT 382.950 598.950 385.050 599.400 ;
        RECT 412.950 598.950 415.050 599.400 ;
        RECT 505.950 600.600 508.050 601.050 ;
        RECT 523.950 600.600 526.050 601.050 ;
        RECT 505.950 599.400 526.050 600.600 ;
        RECT 505.950 598.950 508.050 599.400 ;
        RECT 523.950 598.950 526.050 599.400 ;
        RECT 532.950 600.600 535.050 601.050 ;
        RECT 541.950 600.600 544.050 601.050 ;
        RECT 532.950 599.400 544.050 600.600 ;
        RECT 532.950 598.950 535.050 599.400 ;
        RECT 541.950 598.950 544.050 599.400 ;
        RECT 568.950 600.600 571.050 601.050 ;
        RECT 580.950 600.600 583.050 601.050 ;
        RECT 586.950 600.600 589.050 601.050 ;
        RECT 568.950 599.400 589.050 600.600 ;
        RECT 568.950 598.950 571.050 599.400 ;
        RECT 580.950 598.950 583.050 599.400 ;
        RECT 586.950 598.950 589.050 599.400 ;
        RECT 616.950 600.600 619.050 601.050 ;
        RECT 667.950 600.600 670.050 601.050 ;
        RECT 616.950 599.400 670.050 600.600 ;
        RECT 616.950 598.950 619.050 599.400 ;
        RECT 667.950 598.950 670.050 599.400 ;
        RECT 178.950 597.600 181.050 598.050 ;
        RECT 223.950 597.600 226.050 598.050 ;
        RECT 178.950 596.400 226.050 597.600 ;
        RECT 178.950 595.950 181.050 596.400 ;
        RECT 223.950 595.950 226.050 596.400 ;
        RECT 466.950 597.600 469.050 598.050 ;
        RECT 475.950 597.600 478.050 598.050 ;
        RECT 694.950 597.600 697.050 598.050 ;
        RECT 466.950 596.400 478.050 597.600 ;
        RECT 466.950 595.950 469.050 596.400 ;
        RECT 475.950 595.950 478.050 596.400 ;
        RECT 653.400 596.400 697.050 597.600 ;
        RECT 653.400 595.050 654.600 596.400 ;
        RECT 694.950 595.950 697.050 596.400 ;
        RECT 142.950 594.600 145.050 595.050 ;
        RECT 184.950 594.600 187.050 595.050 ;
        RECT 202.950 594.600 205.050 595.050 ;
        RECT 142.950 593.400 205.050 594.600 ;
        RECT 142.950 592.950 145.050 593.400 ;
        RECT 184.950 592.950 187.050 593.400 ;
        RECT 202.950 592.950 205.050 593.400 ;
        RECT 262.950 594.600 265.050 595.050 ;
        RECT 295.950 594.600 298.050 595.050 ;
        RECT 262.950 593.400 298.050 594.600 ;
        RECT 262.950 592.950 265.050 593.400 ;
        RECT 295.950 592.950 298.050 593.400 ;
        RECT 301.950 594.600 304.050 595.050 ;
        RECT 454.950 594.600 457.050 595.050 ;
        RECT 463.950 594.600 466.050 595.050 ;
        RECT 301.950 593.400 466.050 594.600 ;
        RECT 301.950 592.950 304.050 593.400 ;
        RECT 454.950 592.950 457.050 593.400 ;
        RECT 463.950 592.950 466.050 593.400 ;
        RECT 496.950 594.600 499.050 595.050 ;
        RECT 502.950 594.600 505.050 595.050 ;
        RECT 496.950 593.400 505.050 594.600 ;
        RECT 496.950 592.950 499.050 593.400 ;
        RECT 502.950 592.950 505.050 593.400 ;
        RECT 652.950 592.950 655.050 595.050 ;
        RECT 658.950 594.600 661.050 595.050 ;
        RECT 670.950 594.600 673.050 595.050 ;
        RECT 658.950 593.400 673.050 594.600 ;
        RECT 658.950 592.950 661.050 593.400 ;
        RECT 670.950 592.950 673.050 593.400 ;
        RECT 697.950 594.600 700.050 595.050 ;
        RECT 703.950 594.600 706.050 595.050 ;
        RECT 721.950 594.600 724.050 595.050 ;
        RECT 697.950 593.400 724.050 594.600 ;
        RECT 697.950 592.950 700.050 593.400 ;
        RECT 703.950 592.950 706.050 593.400 ;
        RECT 721.950 592.950 724.050 593.400 ;
        RECT 415.950 591.600 418.050 592.050 ;
        RECT 427.950 591.600 430.050 592.050 ;
        RECT 415.950 590.400 430.050 591.600 ;
        RECT 415.950 589.950 418.050 590.400 ;
        RECT 427.950 589.950 430.050 590.400 ;
        RECT 376.950 588.600 379.050 589.050 ;
        RECT 649.950 588.600 652.050 589.050 ;
        RECT 376.950 587.400 652.050 588.600 ;
        RECT 376.950 586.950 379.050 587.400 ;
        RECT 649.950 586.950 652.050 587.400 ;
        RECT 208.950 582.600 211.050 583.050 ;
        RECT 214.950 582.600 217.050 583.050 ;
        RECT 208.950 581.400 217.050 582.600 ;
        RECT 208.950 580.950 211.050 581.400 ;
        RECT 214.950 580.950 217.050 581.400 ;
        RECT 313.950 570.600 316.050 571.050 ;
        RECT 526.950 570.600 529.050 571.050 ;
        RECT 529.950 570.600 532.050 571.050 ;
        RECT 313.950 569.400 532.050 570.600 ;
        RECT 313.950 568.950 316.050 569.400 ;
        RECT 526.950 568.950 529.050 569.400 ;
        RECT 529.950 568.950 532.050 569.400 ;
        RECT 424.950 567.600 427.050 568.050 ;
        RECT 574.950 567.600 577.050 568.050 ;
        RECT 424.950 566.400 577.050 567.600 ;
        RECT 424.950 565.950 427.050 566.400 ;
        RECT 574.950 565.950 577.050 566.400 ;
        RECT 43.950 564.600 46.050 565.050 ;
        RECT 151.950 564.600 154.050 565.050 ;
        RECT 43.950 563.400 154.050 564.600 ;
        RECT 43.950 562.950 46.050 563.400 ;
        RECT 151.950 562.950 154.050 563.400 ;
        RECT 457.950 564.600 460.050 565.050 ;
        RECT 490.950 564.600 493.050 565.050 ;
        RECT 457.950 563.400 493.050 564.600 ;
        RECT 457.950 562.950 460.050 563.400 ;
        RECT 490.950 562.950 493.050 563.400 ;
        RECT 64.950 561.600 67.050 562.050 ;
        RECT 70.950 561.600 73.050 562.050 ;
        RECT 64.950 560.400 73.050 561.600 ;
        RECT 64.950 559.950 67.050 560.400 ;
        RECT 70.950 559.950 73.050 560.400 ;
        RECT 412.950 561.600 415.050 562.050 ;
        RECT 433.950 561.600 436.050 562.050 ;
        RECT 457.950 561.600 460.050 562.050 ;
        RECT 460.950 561.600 463.050 562.050 ;
        RECT 412.950 560.400 432.600 561.600 ;
        RECT 412.950 559.950 415.050 560.400 ;
        RECT 115.950 558.600 118.050 559.050 ;
        RECT 127.950 558.600 130.050 559.050 ;
        RECT 115.950 557.400 130.050 558.600 ;
        RECT 115.950 556.950 118.050 557.400 ;
        RECT 127.950 556.950 130.050 557.400 ;
        RECT 232.950 558.600 235.050 559.050 ;
        RECT 250.950 558.600 253.050 559.050 ;
        RECT 349.950 558.600 352.050 559.050 ;
        RECT 373.950 558.600 376.050 559.050 ;
        RECT 418.950 558.600 421.050 559.050 ;
        RECT 232.950 557.400 336.600 558.600 ;
        RECT 232.950 556.950 235.050 557.400 ;
        RECT 250.950 556.950 253.050 557.400 ;
        RECT 49.950 555.600 52.050 556.050 ;
        RECT 70.950 555.600 73.050 556.050 ;
        RECT 49.950 554.400 73.050 555.600 ;
        RECT 49.950 553.950 52.050 554.400 ;
        RECT 70.950 553.950 73.050 554.400 ;
        RECT 79.950 555.600 82.050 556.050 ;
        RECT 112.950 555.600 115.050 556.050 ;
        RECT 79.950 554.400 115.050 555.600 ;
        RECT 79.950 553.950 82.050 554.400 ;
        RECT 112.950 553.950 115.050 554.400 ;
        RECT 253.950 555.600 256.050 556.050 ;
        RECT 259.950 555.600 262.050 556.050 ;
        RECT 253.950 554.400 262.050 555.600 ;
        RECT 335.400 555.600 336.600 557.400 ;
        RECT 349.950 557.400 421.050 558.600 ;
        RECT 431.400 558.600 432.600 560.400 ;
        RECT 433.950 560.400 463.050 561.600 ;
        RECT 433.950 559.950 436.050 560.400 ;
        RECT 457.950 559.950 460.050 560.400 ;
        RECT 460.950 559.950 463.050 560.400 ;
        RECT 466.950 561.600 469.050 562.050 ;
        RECT 475.950 561.600 478.050 562.050 ;
        RECT 466.950 560.400 478.050 561.600 ;
        RECT 466.950 559.950 469.050 560.400 ;
        RECT 475.950 559.950 478.050 560.400 ;
        RECT 511.950 561.600 514.050 562.050 ;
        RECT 547.950 561.600 550.050 562.050 ;
        RECT 610.950 561.600 613.050 562.050 ;
        RECT 511.950 560.400 613.050 561.600 ;
        RECT 511.950 559.950 514.050 560.400 ;
        RECT 547.950 559.950 550.050 560.400 ;
        RECT 610.950 559.950 613.050 560.400 ;
        RECT 649.950 561.600 652.050 562.050 ;
        RECT 667.950 561.600 670.050 562.050 ;
        RECT 700.950 561.600 703.050 562.050 ;
        RECT 649.950 560.400 703.050 561.600 ;
        RECT 649.950 559.950 652.050 560.400 ;
        RECT 667.950 559.950 670.050 560.400 ;
        RECT 700.950 559.950 703.050 560.400 ;
        RECT 454.950 558.600 457.050 559.050 ;
        RECT 463.950 558.600 466.050 559.050 ;
        RECT 431.400 557.400 466.050 558.600 ;
        RECT 349.950 556.950 352.050 557.400 ;
        RECT 373.950 556.950 376.050 557.400 ;
        RECT 418.950 556.950 421.050 557.400 ;
        RECT 454.950 556.950 457.050 557.400 ;
        RECT 463.950 556.950 466.050 557.400 ;
        RECT 493.950 558.600 496.050 559.050 ;
        RECT 499.950 558.600 502.050 559.050 ;
        RECT 493.950 557.400 502.050 558.600 ;
        RECT 493.950 556.950 496.050 557.400 ;
        RECT 499.950 556.950 502.050 557.400 ;
        RECT 505.950 556.950 508.050 559.050 ;
        RECT 571.950 558.600 574.050 559.050 ;
        RECT 583.950 558.600 586.050 559.050 ;
        RECT 628.950 558.600 631.050 559.050 ;
        RECT 571.950 557.400 586.050 558.600 ;
        RECT 571.950 556.950 574.050 557.400 ;
        RECT 583.950 556.950 586.050 557.400 ;
        RECT 590.400 557.400 631.050 558.600 ;
        RECT 430.950 555.600 433.050 556.050 ;
        RECT 506.400 555.600 507.600 556.950 ;
        RECT 590.400 555.600 591.600 557.400 ;
        RECT 628.950 556.950 631.050 557.400 ;
        RECT 664.950 558.600 667.050 559.050 ;
        RECT 670.950 558.600 673.050 559.050 ;
        RECT 664.950 557.400 673.050 558.600 ;
        RECT 664.950 556.950 667.050 557.400 ;
        RECT 670.950 556.950 673.050 557.400 ;
        RECT 335.400 554.400 591.600 555.600 ;
        RECT 592.950 555.600 595.050 556.050 ;
        RECT 625.950 555.600 628.050 556.050 ;
        RECT 592.950 554.400 628.050 555.600 ;
        RECT 253.950 553.950 256.050 554.400 ;
        RECT 259.950 553.950 262.050 554.400 ;
        RECT 430.950 553.950 433.050 554.400 ;
        RECT 592.950 553.950 595.050 554.400 ;
        RECT 625.950 553.950 628.050 554.400 ;
        RECT 31.950 552.600 34.050 553.050 ;
        RECT 76.950 552.600 79.050 553.050 ;
        RECT 31.950 551.400 79.050 552.600 ;
        RECT 31.950 550.950 34.050 551.400 ;
        RECT 76.950 550.950 79.050 551.400 ;
        RECT 118.950 552.600 121.050 553.050 ;
        RECT 154.950 552.600 157.050 553.050 ;
        RECT 118.950 551.400 157.050 552.600 ;
        RECT 118.950 550.950 121.050 551.400 ;
        RECT 154.950 550.950 157.050 551.400 ;
        RECT 187.950 552.600 190.050 553.050 ;
        RECT 193.950 552.600 196.050 553.050 ;
        RECT 187.950 551.400 196.050 552.600 ;
        RECT 187.950 550.950 190.050 551.400 ;
        RECT 193.950 550.950 196.050 551.400 ;
        RECT 385.950 552.600 388.050 553.050 ;
        RECT 412.950 552.600 415.050 553.050 ;
        RECT 385.950 551.400 415.050 552.600 ;
        RECT 385.950 550.950 388.050 551.400 ;
        RECT 412.950 550.950 415.050 551.400 ;
        RECT 436.950 552.600 439.050 553.050 ;
        RECT 508.950 552.600 511.050 553.050 ;
        RECT 532.950 552.600 535.050 553.050 ;
        RECT 436.950 551.400 535.050 552.600 ;
        RECT 436.950 550.950 439.050 551.400 ;
        RECT 508.950 550.950 511.050 551.400 ;
        RECT 532.950 550.950 535.050 551.400 ;
        RECT 544.950 552.600 547.050 553.050 ;
        RECT 586.950 552.600 589.050 553.050 ;
        RECT 544.950 551.400 589.050 552.600 ;
        RECT 544.950 550.950 547.050 551.400 ;
        RECT 586.950 550.950 589.050 551.400 ;
        RECT 589.950 552.600 592.050 553.050 ;
        RECT 658.950 552.600 661.050 553.050 ;
        RECT 706.950 552.600 709.050 553.050 ;
        RECT 736.950 552.600 739.050 553.050 ;
        RECT 589.950 551.400 739.050 552.600 ;
        RECT 589.950 550.950 592.050 551.400 ;
        RECT 658.950 550.950 661.050 551.400 ;
        RECT 706.950 550.950 709.050 551.400 ;
        RECT 736.950 550.950 739.050 551.400 ;
        RECT 112.950 549.600 115.050 550.050 ;
        RECT 124.950 549.600 127.050 550.050 ;
        RECT 112.950 548.400 127.050 549.600 ;
        RECT 112.950 547.950 115.050 548.400 ;
        RECT 124.950 547.950 127.050 548.400 ;
        RECT 217.950 549.600 220.050 550.050 ;
        RECT 247.950 549.600 250.050 550.050 ;
        RECT 277.950 549.600 280.050 550.050 ;
        RECT 217.950 548.400 280.050 549.600 ;
        RECT 217.950 547.950 220.050 548.400 ;
        RECT 247.950 547.950 250.050 548.400 ;
        RECT 277.950 547.950 280.050 548.400 ;
        RECT 220.950 546.600 223.050 547.050 ;
        RECT 256.950 546.600 259.050 547.050 ;
        RECT 220.950 545.400 259.050 546.600 ;
        RECT 220.950 544.950 223.050 545.400 ;
        RECT 256.950 544.950 259.050 545.400 ;
        RECT 346.950 546.600 349.050 547.050 ;
        RECT 382.950 546.600 385.050 547.050 ;
        RECT 346.950 545.400 385.050 546.600 ;
        RECT 346.950 544.950 349.050 545.400 ;
        RECT 382.950 544.950 385.050 545.400 ;
        RECT 388.950 546.600 391.050 547.050 ;
        RECT 391.950 546.600 394.050 547.050 ;
        RECT 427.950 546.600 430.050 547.050 ;
        RECT 388.950 545.400 430.050 546.600 ;
        RECT 388.950 544.950 391.050 545.400 ;
        RECT 391.950 544.950 394.050 545.400 ;
        RECT 427.950 544.950 430.050 545.400 ;
        RECT 373.950 534.600 376.050 535.050 ;
        RECT 379.950 534.600 382.050 535.050 ;
        RECT 373.950 533.400 382.050 534.600 ;
        RECT 373.950 532.950 376.050 533.400 ;
        RECT 379.950 532.950 382.050 533.400 ;
        RECT 37.950 531.600 40.050 532.050 ;
        RECT 67.950 531.600 70.050 532.050 ;
        RECT 73.950 531.600 76.050 532.050 ;
        RECT 37.950 530.400 76.050 531.600 ;
        RECT 37.950 529.950 40.050 530.400 ;
        RECT 67.950 529.950 70.050 530.400 ;
        RECT 73.950 529.950 76.050 530.400 ;
        RECT 115.950 531.600 118.050 532.050 ;
        RECT 154.950 531.600 157.050 532.050 ;
        RECT 115.950 530.400 157.050 531.600 ;
        RECT 115.950 529.950 118.050 530.400 ;
        RECT 154.950 529.950 157.050 530.400 ;
        RECT 313.950 531.600 316.050 532.050 ;
        RECT 346.950 531.600 349.050 532.050 ;
        RECT 313.950 530.400 349.050 531.600 ;
        RECT 313.950 529.950 316.050 530.400 ;
        RECT 346.950 529.950 349.050 530.400 ;
        RECT 370.950 531.600 373.050 532.050 ;
        RECT 382.950 531.600 385.050 532.050 ;
        RECT 370.950 530.400 385.050 531.600 ;
        RECT 370.950 529.950 373.050 530.400 ;
        RECT 382.950 529.950 385.050 530.400 ;
        RECT 535.950 531.600 538.050 532.050 ;
        RECT 580.950 531.600 583.050 532.050 ;
        RECT 535.950 530.400 583.050 531.600 ;
        RECT 535.950 529.950 538.050 530.400 ;
        RECT 580.950 529.950 583.050 530.400 ;
        RECT 661.950 531.600 664.050 532.050 ;
        RECT 691.950 531.600 694.050 532.050 ;
        RECT 709.950 531.600 712.050 532.050 ;
        RECT 661.950 530.400 712.050 531.600 ;
        RECT 661.950 529.950 664.050 530.400 ;
        RECT 691.950 529.950 694.050 530.400 ;
        RECT 709.950 529.950 712.050 530.400 ;
        RECT 718.950 531.600 721.050 532.050 ;
        RECT 733.950 531.600 736.050 532.050 ;
        RECT 736.950 531.600 739.050 532.050 ;
        RECT 718.950 530.400 739.050 531.600 ;
        RECT 718.950 529.950 721.050 530.400 ;
        RECT 733.950 529.950 736.050 530.400 ;
        RECT 736.950 529.950 739.050 530.400 ;
        RECT 34.950 528.600 37.050 529.050 ;
        RECT 64.950 528.600 67.050 529.050 ;
        RECT 106.950 528.600 109.050 529.050 ;
        RECT 34.950 527.400 109.050 528.600 ;
        RECT 34.950 526.950 37.050 527.400 ;
        RECT 64.950 526.950 67.050 527.400 ;
        RECT 106.950 526.950 109.050 527.400 ;
        RECT 187.950 528.600 190.050 529.050 ;
        RECT 226.950 528.600 229.050 529.050 ;
        RECT 187.950 527.400 229.050 528.600 ;
        RECT 187.950 526.950 190.050 527.400 ;
        RECT 226.950 526.950 229.050 527.400 ;
        RECT 265.950 528.600 268.050 529.050 ;
        RECT 271.950 528.600 274.050 529.050 ;
        RECT 265.950 527.400 274.050 528.600 ;
        RECT 265.950 526.950 268.050 527.400 ;
        RECT 271.950 526.950 274.050 527.400 ;
        RECT 277.950 528.600 280.050 529.050 ;
        RECT 343.950 528.600 346.050 529.050 ;
        RECT 277.950 527.400 346.050 528.600 ;
        RECT 277.950 526.950 280.050 527.400 ;
        RECT 343.950 526.950 346.050 527.400 ;
        RECT 388.950 528.600 391.050 529.050 ;
        RECT 421.950 528.600 424.050 529.050 ;
        RECT 388.950 527.400 424.050 528.600 ;
        RECT 388.950 526.950 391.050 527.400 ;
        RECT 421.950 526.950 424.050 527.400 ;
        RECT 424.950 528.600 427.050 529.050 ;
        RECT 475.950 528.600 478.050 529.050 ;
        RECT 424.950 527.400 478.050 528.600 ;
        RECT 424.950 526.950 427.050 527.400 ;
        RECT 475.950 526.950 478.050 527.400 ;
        RECT 499.950 528.600 502.050 529.050 ;
        RECT 505.950 528.600 508.050 529.050 ;
        RECT 499.950 527.400 508.050 528.600 ;
        RECT 499.950 526.950 502.050 527.400 ;
        RECT 505.950 526.950 508.050 527.400 ;
        RECT 511.950 528.600 514.050 529.050 ;
        RECT 517.950 528.600 520.050 529.050 ;
        RECT 511.950 527.400 520.050 528.600 ;
        RECT 511.950 526.950 514.050 527.400 ;
        RECT 517.950 526.950 520.050 527.400 ;
        RECT 523.950 528.600 526.050 529.050 ;
        RECT 529.950 528.600 532.050 529.050 ;
        RECT 601.950 528.600 604.050 529.050 ;
        RECT 604.950 528.600 607.050 529.050 ;
        RECT 523.950 527.400 607.050 528.600 ;
        RECT 523.950 526.950 526.050 527.400 ;
        RECT 529.950 526.950 532.050 527.400 ;
        RECT 601.950 526.950 604.050 527.400 ;
        RECT 604.950 526.950 607.050 527.400 ;
        RECT 70.950 525.600 73.050 526.050 ;
        RECT 79.950 525.600 82.050 526.050 ;
        RECT 70.950 524.400 82.050 525.600 ;
        RECT 70.950 523.950 73.050 524.400 ;
        RECT 79.950 523.950 82.050 524.400 ;
        RECT 256.950 525.600 259.050 526.050 ;
        RECT 268.950 525.600 271.050 526.050 ;
        RECT 256.950 524.400 271.050 525.600 ;
        RECT 256.950 523.950 259.050 524.400 ;
        RECT 268.950 523.950 271.050 524.400 ;
        RECT 310.950 525.600 313.050 526.050 ;
        RECT 373.950 525.600 376.050 526.050 ;
        RECT 379.950 525.600 382.050 526.050 ;
        RECT 310.950 524.400 382.050 525.600 ;
        RECT 310.950 523.950 313.050 524.400 ;
        RECT 373.950 523.950 376.050 524.400 ;
        RECT 379.950 523.950 382.050 524.400 ;
        RECT 385.950 525.600 388.050 526.050 ;
        RECT 391.950 525.600 394.050 526.050 ;
        RECT 385.950 524.400 394.050 525.600 ;
        RECT 385.950 523.950 388.050 524.400 ;
        RECT 391.950 523.950 394.050 524.400 ;
        RECT 466.950 525.600 469.050 526.050 ;
        RECT 487.950 525.600 490.050 526.050 ;
        RECT 466.950 524.400 490.050 525.600 ;
        RECT 466.950 523.950 469.050 524.400 ;
        RECT 487.950 523.950 490.050 524.400 ;
        RECT 493.950 525.600 496.050 526.050 ;
        RECT 502.950 525.600 505.050 526.050 ;
        RECT 565.950 525.600 568.050 526.050 ;
        RECT 493.950 524.400 568.050 525.600 ;
        RECT 493.950 523.950 496.050 524.400 ;
        RECT 502.950 523.950 505.050 524.400 ;
        RECT 565.950 523.950 568.050 524.400 ;
        RECT 583.950 525.600 586.050 526.050 ;
        RECT 646.950 525.600 649.050 526.050 ;
        RECT 583.950 524.400 649.050 525.600 ;
        RECT 583.950 523.950 586.050 524.400 ;
        RECT 646.950 523.950 649.050 524.400 ;
        RECT 67.950 522.600 70.050 523.050 ;
        RECT 109.950 522.600 112.050 523.050 ;
        RECT 67.950 521.400 112.050 522.600 ;
        RECT 67.950 520.950 70.050 521.400 ;
        RECT 109.950 520.950 112.050 521.400 ;
        RECT 229.950 522.600 232.050 523.050 ;
        RECT 316.950 522.600 319.050 523.050 ;
        RECT 229.950 521.400 319.050 522.600 ;
        RECT 229.950 520.950 232.050 521.400 ;
        RECT 316.950 520.950 319.050 521.400 ;
        RECT 421.950 522.600 424.050 523.050 ;
        RECT 427.950 522.600 430.050 523.050 ;
        RECT 463.950 522.600 466.050 523.050 ;
        RECT 421.950 521.400 466.050 522.600 ;
        RECT 421.950 520.950 424.050 521.400 ;
        RECT 427.950 520.950 430.050 521.400 ;
        RECT 463.950 520.950 466.050 521.400 ;
        RECT 508.950 522.600 511.050 523.050 ;
        RECT 538.950 522.600 541.050 523.050 ;
        RECT 508.950 521.400 541.050 522.600 ;
        RECT 508.950 520.950 511.050 521.400 ;
        RECT 538.950 520.950 541.050 521.400 ;
        RECT 565.950 522.600 568.050 523.050 ;
        RECT 580.950 522.600 583.050 523.050 ;
        RECT 565.950 521.400 583.050 522.600 ;
        RECT 565.950 520.950 568.050 521.400 ;
        RECT 580.950 520.950 583.050 521.400 ;
        RECT 586.950 522.600 589.050 523.050 ;
        RECT 592.950 522.600 595.050 523.050 ;
        RECT 649.950 522.600 652.050 523.050 ;
        RECT 586.950 521.400 652.050 522.600 ;
        RECT 586.950 520.950 589.050 521.400 ;
        RECT 592.950 520.950 595.050 521.400 ;
        RECT 649.950 520.950 652.050 521.400 ;
        RECT 652.950 522.600 655.050 523.050 ;
        RECT 661.950 522.600 664.050 523.050 ;
        RECT 652.950 521.400 664.050 522.600 ;
        RECT 652.950 520.950 655.050 521.400 ;
        RECT 661.950 520.950 664.050 521.400 ;
        RECT 457.950 519.600 460.050 520.050 ;
        RECT 469.950 519.600 472.050 520.050 ;
        RECT 457.950 518.400 472.050 519.600 ;
        RECT 457.950 517.950 460.050 518.400 ;
        RECT 469.950 517.950 472.050 518.400 ;
        RECT 658.950 513.600 661.050 514.050 ;
        RECT 712.950 513.600 715.050 514.050 ;
        RECT 658.950 512.400 715.050 513.600 ;
        RECT 658.950 511.950 661.050 512.400 ;
        RECT 712.950 511.950 715.050 512.400 ;
        RECT 160.950 507.600 163.050 508.050 ;
        RECT 274.950 507.600 277.050 508.050 ;
        RECT 286.950 507.600 289.050 508.050 ;
        RECT 160.950 506.400 289.050 507.600 ;
        RECT 160.950 505.950 163.050 506.400 ;
        RECT 274.950 505.950 277.050 506.400 ;
        RECT 286.950 505.950 289.050 506.400 ;
        RECT 73.950 492.600 76.050 493.050 ;
        RECT 82.950 492.600 85.050 493.050 ;
        RECT 73.950 491.400 85.050 492.600 ;
        RECT 73.950 490.950 76.050 491.400 ;
        RECT 82.950 490.950 85.050 491.400 ;
        RECT 292.950 492.600 295.050 493.050 ;
        RECT 310.950 492.600 313.050 493.050 ;
        RECT 292.950 491.400 313.050 492.600 ;
        RECT 292.950 490.950 295.050 491.400 ;
        RECT 310.950 490.950 313.050 491.400 ;
        RECT 337.950 492.600 340.050 493.050 ;
        RECT 427.950 492.600 430.050 493.050 ;
        RECT 508.950 492.600 511.050 493.050 ;
        RECT 337.950 491.400 511.050 492.600 ;
        RECT 337.950 490.950 340.050 491.400 ;
        RECT 427.950 490.950 430.050 491.400 ;
        RECT 508.950 490.950 511.050 491.400 ;
        RECT 646.950 492.600 649.050 493.050 ;
        RECT 655.950 492.600 658.050 493.050 ;
        RECT 646.950 491.400 658.050 492.600 ;
        RECT 646.950 490.950 649.050 491.400 ;
        RECT 655.950 490.950 658.050 491.400 ;
        RECT 733.950 492.600 736.050 493.050 ;
        RECT 739.950 492.600 742.050 493.050 ;
        RECT 733.950 491.400 742.050 492.600 ;
        RECT 733.950 490.950 736.050 491.400 ;
        RECT 739.950 490.950 742.050 491.400 ;
        RECT 76.950 489.600 79.050 490.050 ;
        RECT 106.950 489.600 109.050 490.050 ;
        RECT 76.950 488.400 109.050 489.600 ;
        RECT 76.950 487.950 79.050 488.400 ;
        RECT 106.950 487.950 109.050 488.400 ;
        RECT 256.950 489.600 259.050 490.050 ;
        RECT 304.950 489.600 307.050 490.050 ;
        RECT 256.950 488.400 307.050 489.600 ;
        RECT 256.950 487.950 259.050 488.400 ;
        RECT 304.950 487.950 307.050 488.400 ;
        RECT 487.950 489.600 490.050 490.050 ;
        RECT 580.950 489.600 583.050 490.050 ;
        RECT 487.950 488.400 583.050 489.600 ;
        RECT 487.950 487.950 490.050 488.400 ;
        RECT 580.950 487.950 583.050 488.400 ;
        RECT 589.950 489.600 592.050 490.050 ;
        RECT 703.950 489.600 706.050 490.050 ;
        RECT 589.950 488.400 706.050 489.600 ;
        RECT 589.950 487.950 592.050 488.400 ;
        RECT 703.950 487.950 706.050 488.400 ;
        RECT 730.950 489.600 733.050 490.050 ;
        RECT 730.950 488.400 750.600 489.600 ;
        RECT 730.950 487.950 733.050 488.400 ;
        RECT 749.400 487.050 750.600 488.400 ;
        RECT 25.950 486.600 28.050 487.050 ;
        RECT 115.950 486.600 118.050 487.050 ;
        RECT 148.950 486.600 151.050 487.050 ;
        RECT 250.950 486.600 253.050 487.050 ;
        RECT 274.950 486.600 277.050 487.050 ;
        RECT 277.950 486.600 280.050 487.050 ;
        RECT 25.950 485.400 153.600 486.600 ;
        RECT 25.950 484.950 28.050 485.400 ;
        RECT 115.950 484.950 118.050 485.400 ;
        RECT 148.950 484.950 151.050 485.400 ;
        RECT 152.400 484.050 153.600 485.400 ;
        RECT 250.950 485.400 280.050 486.600 ;
        RECT 250.950 484.950 253.050 485.400 ;
        RECT 274.950 484.950 277.050 485.400 ;
        RECT 277.950 484.950 280.050 485.400 ;
        RECT 463.950 486.600 466.050 487.050 ;
        RECT 472.950 486.600 475.050 487.050 ;
        RECT 496.950 486.600 499.050 487.050 ;
        RECT 463.950 485.400 499.050 486.600 ;
        RECT 463.950 484.950 466.050 485.400 ;
        RECT 472.950 484.950 475.050 485.400 ;
        RECT 496.950 484.950 499.050 485.400 ;
        RECT 649.950 486.600 652.050 487.050 ;
        RECT 661.950 486.600 664.050 487.050 ;
        RECT 649.950 485.400 664.050 486.600 ;
        RECT 649.950 484.950 652.050 485.400 ;
        RECT 661.950 484.950 664.050 485.400 ;
        RECT 685.950 486.600 688.050 487.050 ;
        RECT 697.950 486.600 700.050 487.050 ;
        RECT 685.950 485.400 700.050 486.600 ;
        RECT 685.950 484.950 688.050 485.400 ;
        RECT 697.950 484.950 700.050 485.400 ;
        RECT 727.950 486.600 730.050 487.050 ;
        RECT 742.950 486.600 745.050 487.050 ;
        RECT 727.950 485.400 745.050 486.600 ;
        RECT 727.950 484.950 730.050 485.400 ;
        RECT 742.950 484.950 745.050 485.400 ;
        RECT 748.950 484.950 751.050 487.050 ;
        RECT 37.950 483.600 40.050 484.050 ;
        RECT 76.950 483.600 79.050 484.050 ;
        RECT 109.950 483.600 112.050 484.050 ;
        RECT 37.950 482.400 79.050 483.600 ;
        RECT 37.950 481.950 40.050 482.400 ;
        RECT 76.950 481.950 79.050 482.400 ;
        RECT 101.400 482.400 112.050 483.600 ;
        RECT 73.950 480.600 76.050 481.050 ;
        RECT 79.950 480.600 82.050 481.050 ;
        RECT 101.400 480.600 102.600 482.400 ;
        RECT 109.950 481.950 112.050 482.400 ;
        RECT 151.950 481.950 154.050 484.050 ;
        RECT 211.950 483.600 214.050 484.050 ;
        RECT 265.950 483.600 268.050 484.050 ;
        RECT 211.950 482.400 268.050 483.600 ;
        RECT 211.950 481.950 214.050 482.400 ;
        RECT 265.950 481.950 268.050 482.400 ;
        RECT 430.950 483.600 433.050 484.050 ;
        RECT 436.950 483.600 439.050 484.050 ;
        RECT 430.950 482.400 439.050 483.600 ;
        RECT 430.950 481.950 433.050 482.400 ;
        RECT 436.950 481.950 439.050 482.400 ;
        RECT 505.950 483.600 508.050 484.050 ;
        RECT 532.950 483.600 535.050 484.050 ;
        RECT 505.950 482.400 535.050 483.600 ;
        RECT 505.950 481.950 508.050 482.400 ;
        RECT 532.950 481.950 535.050 482.400 ;
        RECT 550.950 483.600 553.050 484.050 ;
        RECT 592.950 483.600 595.050 484.050 ;
        RECT 550.950 482.400 595.050 483.600 ;
        RECT 550.950 481.950 553.050 482.400 ;
        RECT 592.950 481.950 595.050 482.400 ;
        RECT 613.950 483.600 616.050 484.050 ;
        RECT 658.950 483.600 661.050 484.050 ;
        RECT 613.950 482.400 661.050 483.600 ;
        RECT 613.950 481.950 616.050 482.400 ;
        RECT 658.950 481.950 661.050 482.400 ;
        RECT 664.950 483.600 667.050 484.050 ;
        RECT 706.950 483.600 709.050 484.050 ;
        RECT 664.950 482.400 709.050 483.600 ;
        RECT 664.950 481.950 667.050 482.400 ;
        RECT 706.950 481.950 709.050 482.400 ;
        RECT 709.950 483.600 712.050 484.050 ;
        RECT 733.950 483.600 736.050 484.050 ;
        RECT 739.950 483.600 742.050 484.050 ;
        RECT 709.950 482.400 742.050 483.600 ;
        RECT 709.950 481.950 712.050 482.400 ;
        RECT 733.950 481.950 736.050 482.400 ;
        RECT 739.950 481.950 742.050 482.400 ;
        RECT 73.950 479.400 102.600 480.600 ;
        RECT 106.950 480.600 109.050 481.050 ;
        RECT 118.950 480.600 121.050 481.050 ;
        RECT 157.950 480.600 160.050 481.050 ;
        RECT 106.950 479.400 160.050 480.600 ;
        RECT 73.950 478.950 76.050 479.400 ;
        RECT 79.950 478.950 82.050 479.400 ;
        RECT 106.950 478.950 109.050 479.400 ;
        RECT 118.950 478.950 121.050 479.400 ;
        RECT 157.950 478.950 160.050 479.400 ;
        RECT 193.950 480.600 196.050 481.050 ;
        RECT 256.950 480.600 259.050 481.050 ;
        RECT 193.950 479.400 259.050 480.600 ;
        RECT 193.950 478.950 196.050 479.400 ;
        RECT 256.950 478.950 259.050 479.400 ;
        RECT 271.950 480.600 274.050 481.050 ;
        RECT 286.950 480.600 289.050 481.050 ;
        RECT 271.950 479.400 289.050 480.600 ;
        RECT 271.950 478.950 274.050 479.400 ;
        RECT 286.950 478.950 289.050 479.400 ;
        RECT 337.950 480.600 340.050 481.050 ;
        RECT 382.950 480.600 385.050 481.050 ;
        RECT 337.950 479.400 385.050 480.600 ;
        RECT 337.950 478.950 340.050 479.400 ;
        RECT 382.950 478.950 385.050 479.400 ;
        RECT 460.950 480.600 463.050 481.050 ;
        RECT 511.950 480.600 514.050 481.050 ;
        RECT 460.950 479.400 514.050 480.600 ;
        RECT 460.950 478.950 463.050 479.400 ;
        RECT 511.950 478.950 514.050 479.400 ;
        RECT 694.950 480.600 697.050 481.050 ;
        RECT 700.950 480.600 703.050 481.050 ;
        RECT 694.950 479.400 703.050 480.600 ;
        RECT 694.950 478.950 697.050 479.400 ;
        RECT 700.950 478.950 703.050 479.400 ;
        RECT 712.950 480.600 715.050 481.050 ;
        RECT 745.950 480.600 748.050 481.050 ;
        RECT 712.950 479.400 748.050 480.600 ;
        RECT 712.950 478.950 715.050 479.400 ;
        RECT 745.950 478.950 748.050 479.400 ;
        RECT 232.950 477.600 235.050 478.050 ;
        RECT 244.950 477.600 247.050 478.050 ;
        RECT 232.950 476.400 247.050 477.600 ;
        RECT 232.950 475.950 235.050 476.400 ;
        RECT 244.950 475.950 247.050 476.400 ;
        RECT 499.950 477.600 502.050 478.050 ;
        RECT 511.950 477.600 514.050 478.050 ;
        RECT 589.950 477.600 592.050 478.050 ;
        RECT 499.950 476.400 592.050 477.600 ;
        RECT 499.950 475.950 502.050 476.400 ;
        RECT 511.950 475.950 514.050 476.400 ;
        RECT 589.950 475.950 592.050 476.400 ;
        RECT 610.950 477.600 613.050 478.050 ;
        RECT 622.950 477.600 625.050 478.050 ;
        RECT 610.950 476.400 625.050 477.600 ;
        RECT 610.950 475.950 613.050 476.400 ;
        RECT 622.950 475.950 625.050 476.400 ;
        RECT 346.950 474.600 349.050 475.050 ;
        RECT 385.950 474.600 388.050 475.050 ;
        RECT 571.950 474.600 574.050 475.050 ;
        RECT 346.950 473.400 574.050 474.600 ;
        RECT 346.950 472.950 349.050 473.400 ;
        RECT 385.950 472.950 388.050 473.400 ;
        RECT 571.950 472.950 574.050 473.400 ;
        RECT 112.950 462.600 115.050 463.050 ;
        RECT 118.950 462.600 121.050 463.050 ;
        RECT 112.950 461.400 121.050 462.600 ;
        RECT 112.950 460.950 115.050 461.400 ;
        RECT 118.950 460.950 121.050 461.400 ;
        RECT 331.950 462.600 334.050 463.050 ;
        RECT 379.950 462.600 382.050 463.050 ;
        RECT 331.950 461.400 382.050 462.600 ;
        RECT 331.950 460.950 334.050 461.400 ;
        RECT 379.950 460.950 382.050 461.400 ;
        RECT 385.950 462.600 388.050 463.050 ;
        RECT 466.950 462.600 469.050 463.050 ;
        RECT 385.950 461.400 469.050 462.600 ;
        RECT 385.950 460.950 388.050 461.400 ;
        RECT 466.950 460.950 469.050 461.400 ;
        RECT 583.950 462.600 586.050 463.050 ;
        RECT 595.950 462.600 598.050 463.050 ;
        RECT 583.950 461.400 598.050 462.600 ;
        RECT 583.950 460.950 586.050 461.400 ;
        RECT 595.950 460.950 598.050 461.400 ;
        RECT 601.950 462.600 604.050 463.050 ;
        RECT 628.950 462.600 631.050 463.050 ;
        RECT 601.950 461.400 631.050 462.600 ;
        RECT 601.950 460.950 604.050 461.400 ;
        RECT 628.950 460.950 631.050 461.400 ;
        RECT 727.950 462.600 730.050 463.050 ;
        RECT 748.950 462.600 751.050 463.050 ;
        RECT 727.950 461.400 751.050 462.600 ;
        RECT 727.950 460.950 730.050 461.400 ;
        RECT 748.950 460.950 751.050 461.400 ;
        RECT 31.950 459.600 34.050 460.050 ;
        RECT 70.950 459.600 73.050 460.050 ;
        RECT 73.950 459.600 76.050 460.050 ;
        RECT 124.950 459.600 127.050 460.050 ;
        RECT 31.950 458.400 127.050 459.600 ;
        RECT 31.950 457.950 34.050 458.400 ;
        RECT 70.950 457.950 73.050 458.400 ;
        RECT 73.950 457.950 76.050 458.400 ;
        RECT 124.950 457.950 127.050 458.400 ;
        RECT 130.950 459.600 133.050 460.050 ;
        RECT 151.950 459.600 154.050 460.050 ;
        RECT 130.950 458.400 154.050 459.600 ;
        RECT 130.950 457.950 133.050 458.400 ;
        RECT 151.950 457.950 154.050 458.400 ;
        RECT 325.950 459.600 328.050 460.050 ;
        RECT 355.950 459.600 358.050 460.050 ;
        RECT 325.950 458.400 358.050 459.600 ;
        RECT 325.950 457.950 328.050 458.400 ;
        RECT 355.950 457.950 358.050 458.400 ;
        RECT 430.950 459.600 433.050 460.050 ;
        RECT 463.950 459.600 466.050 460.050 ;
        RECT 430.950 458.400 466.050 459.600 ;
        RECT 430.950 457.950 433.050 458.400 ;
        RECT 463.950 457.950 466.050 458.400 ;
        RECT 469.950 459.600 472.050 460.050 ;
        RECT 544.950 459.600 547.050 460.050 ;
        RECT 469.950 458.400 547.050 459.600 ;
        RECT 469.950 457.950 472.050 458.400 ;
        RECT 544.950 457.950 547.050 458.400 ;
        RECT 586.950 459.600 589.050 460.050 ;
        RECT 619.950 459.600 622.050 460.050 ;
        RECT 586.950 458.400 622.050 459.600 ;
        RECT 586.950 457.950 589.050 458.400 ;
        RECT 619.950 457.950 622.050 458.400 ;
        RECT 637.950 459.600 640.050 460.050 ;
        RECT 670.950 459.600 673.050 460.050 ;
        RECT 706.950 459.600 709.050 460.050 ;
        RECT 637.950 458.400 709.050 459.600 ;
        RECT 637.950 457.950 640.050 458.400 ;
        RECT 670.950 457.950 673.050 458.400 ;
        RECT 706.950 457.950 709.050 458.400 ;
        RECT 712.950 459.600 715.050 460.050 ;
        RECT 745.950 459.600 748.050 460.050 ;
        RECT 712.950 458.400 748.050 459.600 ;
        RECT 712.950 457.950 715.050 458.400 ;
        RECT 745.950 457.950 748.050 458.400 ;
        RECT 28.950 456.600 31.050 457.050 ;
        RECT 37.950 456.600 40.050 457.050 ;
        RECT 28.950 455.400 40.050 456.600 ;
        RECT 28.950 454.950 31.050 455.400 ;
        RECT 37.950 454.950 40.050 455.400 ;
        RECT 76.950 456.600 79.050 457.050 ;
        RECT 145.950 456.600 148.050 457.050 ;
        RECT 76.950 455.400 148.050 456.600 ;
        RECT 76.950 454.950 79.050 455.400 ;
        RECT 110.400 454.050 111.600 455.400 ;
        RECT 145.950 454.950 148.050 455.400 ;
        RECT 217.950 456.600 220.050 457.050 ;
        RECT 310.950 456.600 313.050 457.050 ;
        RECT 313.950 456.600 316.050 457.050 ;
        RECT 331.950 456.600 334.050 457.050 ;
        RECT 217.950 455.400 334.050 456.600 ;
        RECT 217.950 454.950 220.050 455.400 ;
        RECT 310.950 454.950 313.050 455.400 ;
        RECT 313.950 454.950 316.050 455.400 ;
        RECT 331.950 454.950 334.050 455.400 ;
        RECT 367.950 456.600 370.050 457.050 ;
        RECT 427.950 456.600 430.050 457.050 ;
        RECT 367.950 455.400 430.050 456.600 ;
        RECT 367.950 454.950 370.050 455.400 ;
        RECT 427.950 454.950 430.050 455.400 ;
        RECT 490.950 456.600 493.050 457.050 ;
        RECT 499.950 456.600 502.050 457.050 ;
        RECT 490.950 455.400 502.050 456.600 ;
        RECT 490.950 454.950 493.050 455.400 ;
        RECT 499.950 454.950 502.050 455.400 ;
        RECT 550.950 456.600 553.050 457.050 ;
        RECT 592.950 456.600 595.050 457.050 ;
        RECT 550.950 455.400 595.050 456.600 ;
        RECT 550.950 454.950 553.050 455.400 ;
        RECT 592.950 454.950 595.050 455.400 ;
        RECT 679.950 456.600 682.050 457.050 ;
        RECT 703.950 456.600 706.050 457.050 ;
        RECT 736.950 456.600 739.050 457.050 ;
        RECT 679.950 455.400 739.050 456.600 ;
        RECT 679.950 454.950 682.050 455.400 ;
        RECT 703.950 454.950 706.050 455.400 ;
        RECT 736.950 454.950 739.050 455.400 ;
        RECT 70.950 453.600 73.050 454.050 ;
        RECT 103.950 453.600 106.050 454.050 ;
        RECT 70.950 452.400 106.050 453.600 ;
        RECT 70.950 451.950 73.050 452.400 ;
        RECT 103.950 451.950 106.050 452.400 ;
        RECT 109.950 451.950 112.050 454.050 ;
        RECT 124.950 453.600 127.050 454.050 ;
        RECT 148.950 453.600 151.050 454.050 ;
        RECT 124.950 452.400 151.050 453.600 ;
        RECT 124.950 451.950 127.050 452.400 ;
        RECT 148.950 451.950 151.050 452.400 ;
        RECT 211.950 453.600 214.050 454.050 ;
        RECT 217.950 453.600 220.050 454.050 ;
        RECT 211.950 452.400 220.050 453.600 ;
        RECT 211.950 451.950 214.050 452.400 ;
        RECT 217.950 451.950 220.050 452.400 ;
        RECT 358.950 453.600 361.050 454.050 ;
        RECT 376.950 453.600 379.050 454.050 ;
        RECT 358.950 452.400 379.050 453.600 ;
        RECT 358.950 451.950 361.050 452.400 ;
        RECT 376.950 451.950 379.050 452.400 ;
        RECT 421.950 453.600 424.050 454.050 ;
        RECT 541.950 453.600 544.050 454.050 ;
        RECT 565.950 453.600 568.050 454.050 ;
        RECT 583.950 453.600 586.050 454.050 ;
        RECT 421.950 452.400 586.050 453.600 ;
        RECT 421.950 451.950 424.050 452.400 ;
        RECT 541.950 451.950 544.050 452.400 ;
        RECT 565.950 451.950 568.050 452.400 ;
        RECT 583.950 451.950 586.050 452.400 ;
        RECT 589.950 453.600 592.050 454.050 ;
        RECT 601.950 453.600 604.050 454.050 ;
        RECT 589.950 452.400 604.050 453.600 ;
        RECT 589.950 451.950 592.050 452.400 ;
        RECT 601.950 451.950 604.050 452.400 ;
        RECT 619.950 453.600 622.050 454.050 ;
        RECT 625.950 453.600 628.050 454.050 ;
        RECT 619.950 452.400 628.050 453.600 ;
        RECT 619.950 451.950 622.050 452.400 ;
        RECT 625.950 451.950 628.050 452.400 ;
        RECT 631.950 453.600 634.050 454.050 ;
        RECT 664.950 453.600 667.050 454.050 ;
        RECT 631.950 452.400 667.050 453.600 ;
        RECT 631.950 451.950 634.050 452.400 ;
        RECT 664.950 451.950 667.050 452.400 ;
        RECT 733.950 453.600 736.050 454.050 ;
        RECT 742.950 453.600 745.050 454.050 ;
        RECT 733.950 452.400 745.050 453.600 ;
        RECT 733.950 451.950 736.050 452.400 ;
        RECT 742.950 451.950 745.050 452.400 ;
        RECT 508.950 450.600 511.050 451.050 ;
        RECT 547.950 450.600 550.050 451.050 ;
        RECT 508.950 449.400 550.050 450.600 ;
        RECT 508.950 448.950 511.050 449.400 ;
        RECT 547.950 448.950 550.050 449.400 ;
        RECT 667.950 450.600 670.050 451.050 ;
        RECT 712.950 450.600 715.050 451.050 ;
        RECT 667.950 449.400 715.050 450.600 ;
        RECT 667.950 448.950 670.050 449.400 ;
        RECT 712.950 448.950 715.050 449.400 ;
        RECT 544.950 447.600 547.050 448.050 ;
        RECT 568.950 447.600 571.050 448.050 ;
        RECT 544.950 446.400 571.050 447.600 ;
        RECT 544.950 445.950 547.050 446.400 ;
        RECT 568.950 445.950 571.050 446.400 ;
        RECT 103.950 420.600 106.050 421.050 ;
        RECT 115.950 420.600 118.050 421.050 ;
        RECT 103.950 419.400 118.050 420.600 ;
        RECT 103.950 418.950 106.050 419.400 ;
        RECT 115.950 418.950 118.050 419.400 ;
        RECT 109.950 417.600 112.050 418.050 ;
        RECT 130.950 417.600 133.050 418.050 ;
        RECT 109.950 416.400 133.050 417.600 ;
        RECT 109.950 415.950 112.050 416.400 ;
        RECT 130.950 415.950 133.050 416.400 ;
        RECT 220.950 417.600 223.050 418.050 ;
        RECT 250.950 417.600 253.050 418.050 ;
        RECT 292.950 417.600 295.050 418.050 ;
        RECT 220.950 416.400 295.050 417.600 ;
        RECT 220.950 415.950 223.050 416.400 ;
        RECT 250.950 415.950 253.050 416.400 ;
        RECT 292.950 415.950 295.050 416.400 ;
        RECT 298.950 417.600 301.050 418.050 ;
        RECT 367.950 417.600 370.050 418.050 ;
        RECT 298.950 416.400 370.050 417.600 ;
        RECT 298.950 415.950 301.050 416.400 ;
        RECT 367.950 415.950 370.050 416.400 ;
        RECT 562.950 417.600 565.050 418.050 ;
        RECT 604.950 417.600 607.050 418.050 ;
        RECT 562.950 416.400 607.050 417.600 ;
        RECT 562.950 415.950 565.050 416.400 ;
        RECT 604.950 415.950 607.050 416.400 ;
        RECT 643.950 417.600 646.050 418.050 ;
        RECT 661.950 417.600 664.050 418.050 ;
        RECT 643.950 416.400 664.050 417.600 ;
        RECT 643.950 415.950 646.050 416.400 ;
        RECT 661.950 415.950 664.050 416.400 ;
        RECT 31.950 414.600 34.050 415.050 ;
        RECT 37.950 414.600 40.050 415.050 ;
        RECT 31.950 413.400 40.050 414.600 ;
        RECT 31.950 412.950 34.050 413.400 ;
        RECT 37.950 412.950 40.050 413.400 ;
        RECT 46.950 414.600 49.050 415.050 ;
        RECT 70.950 414.600 73.050 415.050 ;
        RECT 46.950 413.400 73.050 414.600 ;
        RECT 46.950 412.950 49.050 413.400 ;
        RECT 70.950 412.950 73.050 413.400 ;
        RECT 76.950 414.600 79.050 415.050 ;
        RECT 112.950 414.600 115.050 415.050 ;
        RECT 76.950 413.400 115.050 414.600 ;
        RECT 76.950 412.950 79.050 413.400 ;
        RECT 112.950 412.950 115.050 413.400 ;
        RECT 325.950 414.600 328.050 415.050 ;
        RECT 403.950 414.600 406.050 415.050 ;
        RECT 325.950 413.400 406.050 414.600 ;
        RECT 325.950 412.950 328.050 413.400 ;
        RECT 403.950 412.950 406.050 413.400 ;
        RECT 424.950 414.600 427.050 415.050 ;
        RECT 442.950 414.600 445.050 415.050 ;
        RECT 424.950 413.400 445.050 414.600 ;
        RECT 424.950 412.950 427.050 413.400 ;
        RECT 442.950 412.950 445.050 413.400 ;
        RECT 484.950 414.600 487.050 415.050 ;
        RECT 532.950 414.600 535.050 415.050 ;
        RECT 484.950 413.400 535.050 414.600 ;
        RECT 484.950 412.950 487.050 413.400 ;
        RECT 532.950 412.950 535.050 413.400 ;
        RECT 640.950 414.600 643.050 415.050 ;
        RECT 658.950 414.600 661.050 415.050 ;
        RECT 640.950 413.400 661.050 414.600 ;
        RECT 640.950 412.950 643.050 413.400 ;
        RECT 658.950 412.950 661.050 413.400 ;
        RECT 661.950 414.600 664.050 415.050 ;
        RECT 673.950 414.600 676.050 415.050 ;
        RECT 661.950 413.400 676.050 414.600 ;
        RECT 661.950 412.950 664.050 413.400 ;
        RECT 673.950 412.950 676.050 413.400 ;
        RECT 709.950 414.600 712.050 415.050 ;
        RECT 721.950 414.600 724.050 415.050 ;
        RECT 709.950 413.400 724.050 414.600 ;
        RECT 709.950 412.950 712.050 413.400 ;
        RECT 721.950 412.950 724.050 413.400 ;
        RECT 13.950 411.600 16.050 412.050 ;
        RECT 67.950 411.600 70.050 412.050 ;
        RECT 13.950 410.400 70.050 411.600 ;
        RECT 13.950 409.950 16.050 410.400 ;
        RECT 67.950 409.950 70.050 410.400 ;
        RECT 184.950 409.950 187.050 412.050 ;
        RECT 316.950 411.600 319.050 412.050 ;
        RECT 355.950 411.600 358.050 412.050 ;
        RECT 445.950 411.600 448.050 412.050 ;
        RECT 316.950 410.400 358.050 411.600 ;
        RECT 316.950 409.950 319.050 410.400 ;
        RECT 355.950 409.950 358.050 410.400 ;
        RECT 359.400 410.400 448.050 411.600 ;
        RECT 73.950 408.600 76.050 409.050 ;
        RECT 85.950 408.600 88.050 409.050 ;
        RECT 145.950 408.600 148.050 409.050 ;
        RECT 73.950 407.400 148.050 408.600 ;
        RECT 185.400 408.600 186.600 409.950 ;
        RECT 217.950 408.600 220.050 409.050 ;
        RECT 185.400 407.400 220.050 408.600 ;
        RECT 73.950 406.950 76.050 407.400 ;
        RECT 85.950 406.950 88.050 407.400 ;
        RECT 145.950 406.950 148.050 407.400 ;
        RECT 217.950 406.950 220.050 407.400 ;
        RECT 349.950 408.600 352.050 409.050 ;
        RECT 359.400 408.600 360.600 410.400 ;
        RECT 445.950 409.950 448.050 410.400 ;
        RECT 487.950 411.600 490.050 412.050 ;
        RECT 493.950 411.600 496.050 412.050 ;
        RECT 520.950 411.600 523.050 412.050 ;
        RECT 556.950 411.600 559.050 412.050 ;
        RECT 487.950 410.400 559.050 411.600 ;
        RECT 487.950 409.950 490.050 410.400 ;
        RECT 493.950 409.950 496.050 410.400 ;
        RECT 520.950 409.950 523.050 410.400 ;
        RECT 556.950 409.950 559.050 410.400 ;
        RECT 601.950 411.600 604.050 412.050 ;
        RECT 610.950 411.600 613.050 412.050 ;
        RECT 712.950 411.600 715.050 412.050 ;
        RECT 601.950 410.400 715.050 411.600 ;
        RECT 601.950 409.950 604.050 410.400 ;
        RECT 610.950 409.950 613.050 410.400 ;
        RECT 712.950 409.950 715.050 410.400 ;
        RECT 349.950 407.400 360.600 408.600 ;
        RECT 370.950 408.600 373.050 409.050 ;
        RECT 400.950 408.600 403.050 409.050 ;
        RECT 370.950 407.400 403.050 408.600 ;
        RECT 349.950 406.950 352.050 407.400 ;
        RECT 370.950 406.950 373.050 407.400 ;
        RECT 400.950 406.950 403.050 407.400 ;
        RECT 439.950 408.600 442.050 409.050 ;
        RECT 508.950 408.600 511.050 409.050 ;
        RECT 439.950 407.400 511.050 408.600 ;
        RECT 439.950 406.950 442.050 407.400 ;
        RECT 508.950 406.950 511.050 407.400 ;
        RECT 670.950 408.600 673.050 409.050 ;
        RECT 676.950 408.600 679.050 409.050 ;
        RECT 670.950 407.400 679.050 408.600 ;
        RECT 670.950 406.950 673.050 407.400 ;
        RECT 676.950 406.950 679.050 407.400 ;
        RECT 703.950 408.600 706.050 409.050 ;
        RECT 718.950 408.600 721.050 409.050 ;
        RECT 703.950 407.400 721.050 408.600 ;
        RECT 703.950 406.950 706.050 407.400 ;
        RECT 718.950 406.950 721.050 407.400 ;
        RECT 31.950 405.600 34.050 406.050 ;
        RECT 46.950 405.600 49.050 406.050 ;
        RECT 31.950 404.400 49.050 405.600 ;
        RECT 31.950 403.950 34.050 404.400 ;
        RECT 46.950 403.950 49.050 404.400 ;
        RECT 151.950 405.600 154.050 406.050 ;
        RECT 316.950 405.600 319.050 406.050 ;
        RECT 151.950 404.400 319.050 405.600 ;
        RECT 151.950 403.950 154.050 404.400 ;
        RECT 316.950 403.950 319.050 404.400 ;
        RECT 322.950 399.600 325.050 400.050 ;
        RECT 343.950 399.600 346.050 400.050 ;
        RECT 322.950 398.400 346.050 399.600 ;
        RECT 322.950 397.950 325.050 398.400 ;
        RECT 343.950 397.950 346.050 398.400 ;
        RECT 499.950 399.600 502.050 400.050 ;
        RECT 523.950 399.600 526.050 400.050 ;
        RECT 499.950 398.400 526.050 399.600 ;
        RECT 499.950 397.950 502.050 398.400 ;
        RECT 523.950 397.950 526.050 398.400 ;
        RECT 166.950 396.600 169.050 397.050 ;
        RECT 190.950 396.600 193.050 397.050 ;
        RECT 166.950 395.400 193.050 396.600 ;
        RECT 166.950 394.950 169.050 395.400 ;
        RECT 190.950 394.950 193.050 395.400 ;
        RECT 259.950 396.600 262.050 397.050 ;
        RECT 274.950 396.600 277.050 397.050 ;
        RECT 301.950 396.600 304.050 397.050 ;
        RECT 304.950 396.600 307.050 397.050 ;
        RECT 259.950 395.400 307.050 396.600 ;
        RECT 259.950 394.950 262.050 395.400 ;
        RECT 274.950 394.950 277.050 395.400 ;
        RECT 301.950 394.950 304.050 395.400 ;
        RECT 304.950 394.950 307.050 395.400 ;
        RECT 229.950 393.600 232.050 394.050 ;
        RECT 268.950 393.600 271.050 394.050 ;
        RECT 229.950 392.400 271.050 393.600 ;
        RECT 229.950 391.950 232.050 392.400 ;
        RECT 268.950 391.950 271.050 392.400 ;
        RECT 127.950 390.600 130.050 391.050 ;
        RECT 151.950 390.600 154.050 391.050 ;
        RECT 187.950 390.600 190.050 391.050 ;
        RECT 346.950 390.600 349.050 391.050 ;
        RECT 127.950 389.400 349.050 390.600 ;
        RECT 127.950 388.950 130.050 389.400 ;
        RECT 151.950 388.950 154.050 389.400 ;
        RECT 187.950 388.950 190.050 389.400 ;
        RECT 346.950 388.950 349.050 389.400 ;
        RECT 526.950 390.600 529.050 391.050 ;
        RECT 550.950 390.600 553.050 391.050 ;
        RECT 553.950 390.600 556.050 391.050 ;
        RECT 595.950 390.600 598.050 391.050 ;
        RECT 526.950 389.400 598.050 390.600 ;
        RECT 526.950 388.950 529.050 389.400 ;
        RECT 550.950 388.950 553.050 389.400 ;
        RECT 553.950 388.950 556.050 389.400 ;
        RECT 595.950 388.950 598.050 389.400 ;
        RECT 202.950 387.600 205.050 388.050 ;
        RECT 259.950 387.600 262.050 388.050 ;
        RECT 202.950 386.400 262.050 387.600 ;
        RECT 202.950 385.950 205.050 386.400 ;
        RECT 259.950 385.950 262.050 386.400 ;
        RECT 556.950 387.600 559.050 388.050 ;
        RECT 586.950 387.600 589.050 388.050 ;
        RECT 619.950 387.600 622.050 388.050 ;
        RECT 556.950 386.400 622.050 387.600 ;
        RECT 556.950 385.950 559.050 386.400 ;
        RECT 586.950 385.950 589.050 386.400 ;
        RECT 619.950 385.950 622.050 386.400 ;
        RECT 670.950 387.600 673.050 388.050 ;
        RECT 697.950 387.600 700.050 388.050 ;
        RECT 670.950 386.400 700.050 387.600 ;
        RECT 670.950 385.950 673.050 386.400 ;
        RECT 697.950 385.950 700.050 386.400 ;
        RECT 115.950 384.600 118.050 385.050 ;
        RECT 121.950 384.600 124.050 385.050 ;
        RECT 115.950 383.400 124.050 384.600 ;
        RECT 115.950 382.950 118.050 383.400 ;
        RECT 121.950 382.950 124.050 383.400 ;
        RECT 193.950 384.600 196.050 385.050 ;
        RECT 253.950 384.600 256.050 385.050 ;
        RECT 193.950 383.400 256.050 384.600 ;
        RECT 193.950 382.950 196.050 383.400 ;
        RECT 253.950 382.950 256.050 383.400 ;
        RECT 265.950 384.600 268.050 385.050 ;
        RECT 298.950 384.600 301.050 385.050 ;
        RECT 310.950 384.600 313.050 385.050 ;
        RECT 265.950 383.400 301.050 384.600 ;
        RECT 265.950 382.950 268.050 383.400 ;
        RECT 298.950 382.950 301.050 383.400 ;
        RECT 305.400 383.400 313.050 384.600 ;
        RECT 305.400 382.050 306.600 383.400 ;
        RECT 310.950 382.950 313.050 383.400 ;
        RECT 340.950 384.600 343.050 385.050 ;
        RECT 349.950 384.600 352.050 385.050 ;
        RECT 340.950 383.400 352.050 384.600 ;
        RECT 340.950 382.950 343.050 383.400 ;
        RECT 349.950 382.950 352.050 383.400 ;
        RECT 382.950 384.600 385.050 385.050 ;
        RECT 400.950 384.600 403.050 385.050 ;
        RECT 421.950 384.600 424.050 385.050 ;
        RECT 382.950 383.400 424.050 384.600 ;
        RECT 382.950 382.950 385.050 383.400 ;
        RECT 400.950 382.950 403.050 383.400 ;
        RECT 421.950 382.950 424.050 383.400 ;
        RECT 445.950 384.600 448.050 385.050 ;
        RECT 460.950 384.600 463.050 385.050 ;
        RECT 445.950 383.400 463.050 384.600 ;
        RECT 445.950 382.950 448.050 383.400 ;
        RECT 460.950 382.950 463.050 383.400 ;
        RECT 466.950 384.600 469.050 385.050 ;
        RECT 472.950 384.600 475.050 385.050 ;
        RECT 466.950 383.400 475.050 384.600 ;
        RECT 466.950 382.950 469.050 383.400 ;
        RECT 472.950 382.950 475.050 383.400 ;
        RECT 658.950 384.600 661.050 385.050 ;
        RECT 727.950 384.600 730.050 385.050 ;
        RECT 658.950 383.400 730.050 384.600 ;
        RECT 658.950 382.950 661.050 383.400 ;
        RECT 727.950 382.950 730.050 383.400 ;
        RECT 73.950 381.600 76.050 382.050 ;
        RECT 163.950 381.600 166.050 382.050 ;
        RECT 73.950 380.400 166.050 381.600 ;
        RECT 73.950 379.950 76.050 380.400 ;
        RECT 163.950 379.950 166.050 380.400 ;
        RECT 253.950 381.600 256.050 382.050 ;
        RECT 262.950 381.600 265.050 382.050 ;
        RECT 253.950 380.400 265.050 381.600 ;
        RECT 253.950 379.950 256.050 380.400 ;
        RECT 262.950 379.950 265.050 380.400 ;
        RECT 277.950 381.600 280.050 382.050 ;
        RECT 301.950 381.600 304.050 382.050 ;
        RECT 277.950 380.400 304.050 381.600 ;
        RECT 277.950 379.950 280.050 380.400 ;
        RECT 301.950 379.950 304.050 380.400 ;
        RECT 304.950 379.950 307.050 382.050 ;
        RECT 421.950 381.600 424.050 382.050 ;
        RECT 457.950 381.600 460.050 382.050 ;
        RECT 421.950 380.400 460.050 381.600 ;
        RECT 421.950 379.950 424.050 380.400 ;
        RECT 457.950 379.950 460.050 380.400 ;
        RECT 481.950 381.600 484.050 382.050 ;
        RECT 502.950 381.600 505.050 382.050 ;
        RECT 481.950 380.400 505.050 381.600 ;
        RECT 481.950 379.950 484.050 380.400 ;
        RECT 502.950 379.950 505.050 380.400 ;
        RECT 532.950 381.600 535.050 382.050 ;
        RECT 541.950 381.600 544.050 382.050 ;
        RECT 532.950 380.400 544.050 381.600 ;
        RECT 532.950 379.950 535.050 380.400 ;
        RECT 541.950 379.950 544.050 380.400 ;
        RECT 547.950 381.600 550.050 382.050 ;
        RECT 607.950 381.600 610.050 382.050 ;
        RECT 547.950 380.400 610.050 381.600 ;
        RECT 547.950 379.950 550.050 380.400 ;
        RECT 607.950 379.950 610.050 380.400 ;
        RECT 622.950 381.600 625.050 382.050 ;
        RECT 652.950 381.600 655.050 382.050 ;
        RECT 622.950 380.400 655.050 381.600 ;
        RECT 622.950 379.950 625.050 380.400 ;
        RECT 652.950 379.950 655.050 380.400 ;
        RECT 709.950 381.600 712.050 382.050 ;
        RECT 733.950 381.600 736.050 382.050 ;
        RECT 709.950 380.400 736.050 381.600 ;
        RECT 709.950 379.950 712.050 380.400 ;
        RECT 733.950 379.950 736.050 380.400 ;
        RECT 76.950 378.600 79.050 379.050 ;
        RECT 103.950 378.600 106.050 379.050 ;
        RECT 112.950 378.600 115.050 379.050 ;
        RECT 76.950 377.400 115.050 378.600 ;
        RECT 76.950 376.950 79.050 377.400 ;
        RECT 103.950 376.950 106.050 377.400 ;
        RECT 112.950 376.950 115.050 377.400 ;
        RECT 232.950 378.600 235.050 379.050 ;
        RECT 253.950 378.600 256.050 379.050 ;
        RECT 232.950 377.400 256.050 378.600 ;
        RECT 232.950 376.950 235.050 377.400 ;
        RECT 253.950 376.950 256.050 377.400 ;
        RECT 298.950 378.600 301.050 379.050 ;
        RECT 418.950 378.600 421.050 379.050 ;
        RECT 298.950 377.400 421.050 378.600 ;
        RECT 298.950 376.950 301.050 377.400 ;
        RECT 418.950 376.950 421.050 377.400 ;
        RECT 589.950 378.600 592.050 379.050 ;
        RECT 664.950 378.600 667.050 379.050 ;
        RECT 589.950 377.400 667.050 378.600 ;
        RECT 589.950 376.950 592.050 377.400 ;
        RECT 664.950 376.950 667.050 377.400 ;
        RECT 70.950 375.600 73.050 376.050 ;
        RECT 82.950 375.600 85.050 376.050 ;
        RECT 70.950 374.400 85.050 375.600 ;
        RECT 70.950 373.950 73.050 374.400 ;
        RECT 82.950 373.950 85.050 374.400 ;
        RECT 349.950 375.600 352.050 376.050 ;
        RECT 424.950 375.600 427.050 376.050 ;
        RECT 463.950 375.600 466.050 376.050 ;
        RECT 349.950 374.400 466.050 375.600 ;
        RECT 349.950 373.950 352.050 374.400 ;
        RECT 424.950 373.950 427.050 374.400 ;
        RECT 463.950 373.950 466.050 374.400 ;
        RECT 496.950 375.600 499.050 376.050 ;
        RECT 511.950 375.600 514.050 376.050 ;
        RECT 592.950 375.600 595.050 376.050 ;
        RECT 496.950 374.400 595.050 375.600 ;
        RECT 496.950 373.950 499.050 374.400 ;
        RECT 511.950 373.950 514.050 374.400 ;
        RECT 592.950 373.950 595.050 374.400 ;
        RECT 34.950 372.600 37.050 373.050 ;
        RECT 85.950 372.600 88.050 373.050 ;
        RECT 34.950 371.400 88.050 372.600 ;
        RECT 34.950 370.950 37.050 371.400 ;
        RECT 85.950 370.950 88.050 371.400 ;
        RECT 145.950 351.600 148.050 352.050 ;
        RECT 154.950 351.600 157.050 352.050 ;
        RECT 145.950 350.400 157.050 351.600 ;
        RECT 145.950 349.950 148.050 350.400 ;
        RECT 154.950 349.950 157.050 350.400 ;
        RECT 235.950 351.600 238.050 352.050 ;
        RECT 295.950 351.600 298.050 352.050 ;
        RECT 235.950 350.400 298.050 351.600 ;
        RECT 235.950 349.950 238.050 350.400 ;
        RECT 295.950 349.950 298.050 350.400 ;
        RECT 676.950 348.600 679.050 349.050 ;
        RECT 709.950 348.600 712.050 349.050 ;
        RECT 676.950 347.400 712.050 348.600 ;
        RECT 676.950 346.950 679.050 347.400 ;
        RECT 709.950 346.950 712.050 347.400 ;
        RECT 196.950 345.600 199.050 346.050 ;
        RECT 250.950 345.600 253.050 346.050 ;
        RECT 196.950 344.400 253.050 345.600 ;
        RECT 196.950 343.950 199.050 344.400 ;
        RECT 250.950 343.950 253.050 344.400 ;
        RECT 283.950 345.600 286.050 346.050 ;
        RECT 298.950 345.600 301.050 346.050 ;
        RECT 283.950 344.400 301.050 345.600 ;
        RECT 283.950 343.950 286.050 344.400 ;
        RECT 298.950 343.950 301.050 344.400 ;
        RECT 652.950 345.600 655.050 346.050 ;
        RECT 682.950 345.600 685.050 346.050 ;
        RECT 652.950 344.400 685.050 345.600 ;
        RECT 652.950 343.950 655.050 344.400 ;
        RECT 682.950 343.950 685.050 344.400 ;
        RECT 73.950 342.600 76.050 343.050 ;
        RECT 85.950 342.600 88.050 343.050 ;
        RECT 106.950 342.600 109.050 343.050 ;
        RECT 73.950 341.400 109.050 342.600 ;
        RECT 73.950 340.950 76.050 341.400 ;
        RECT 85.950 340.950 88.050 341.400 ;
        RECT 106.950 340.950 109.050 341.400 ;
        RECT 160.950 342.600 163.050 343.050 ;
        RECT 181.950 342.600 184.050 343.050 ;
        RECT 160.950 341.400 184.050 342.600 ;
        RECT 160.950 340.950 163.050 341.400 ;
        RECT 181.950 340.950 184.050 341.400 ;
        RECT 202.950 342.600 205.050 343.050 ;
        RECT 235.950 342.600 238.050 343.050 ;
        RECT 202.950 341.400 238.050 342.600 ;
        RECT 202.950 340.950 205.050 341.400 ;
        RECT 235.950 340.950 238.050 341.400 ;
        RECT 244.950 342.600 247.050 343.050 ;
        RECT 259.950 342.600 262.050 343.050 ;
        RECT 244.950 341.400 262.050 342.600 ;
        RECT 244.950 340.950 247.050 341.400 ;
        RECT 259.950 340.950 262.050 341.400 ;
        RECT 280.950 340.950 283.050 343.050 ;
        RECT 286.950 342.600 289.050 343.050 ;
        RECT 304.950 342.600 307.050 343.050 ;
        RECT 286.950 341.400 307.050 342.600 ;
        RECT 286.950 340.950 289.050 341.400 ;
        RECT 304.950 340.950 307.050 341.400 ;
        RECT 439.950 342.600 442.050 343.050 ;
        RECT 454.950 342.600 457.050 343.050 ;
        RECT 439.950 341.400 457.050 342.600 ;
        RECT 439.950 340.950 442.050 341.400 ;
        RECT 454.950 340.950 457.050 341.400 ;
        RECT 481.950 340.950 484.050 343.050 ;
        RECT 508.950 342.600 511.050 343.050 ;
        RECT 589.950 342.600 592.050 343.050 ;
        RECT 598.950 342.600 601.050 343.050 ;
        RECT 508.950 341.400 601.050 342.600 ;
        RECT 508.950 340.950 511.050 341.400 ;
        RECT 589.950 340.950 592.050 341.400 ;
        RECT 598.950 340.950 601.050 341.400 ;
        RECT 604.950 340.950 607.050 343.050 ;
        RECT 670.950 342.600 673.050 343.050 ;
        RECT 679.950 342.600 682.050 343.050 ;
        RECT 670.950 341.400 682.050 342.600 ;
        RECT 670.950 340.950 673.050 341.400 ;
        RECT 679.950 340.950 682.050 341.400 ;
        RECT 718.950 342.600 721.050 343.050 ;
        RECT 730.950 342.600 733.050 343.050 ;
        RECT 718.950 341.400 733.050 342.600 ;
        RECT 718.950 340.950 721.050 341.400 ;
        RECT 730.950 340.950 733.050 341.400 ;
        RECT 52.950 339.600 55.050 340.050 ;
        RECT 115.950 339.600 118.050 340.050 ;
        RECT 142.950 339.600 145.050 340.050 ;
        RECT 172.950 339.600 175.050 340.050 ;
        RECT 52.950 338.400 175.050 339.600 ;
        RECT 52.950 337.950 55.050 338.400 ;
        RECT 115.950 337.950 118.050 338.400 ;
        RECT 142.950 337.950 145.050 338.400 ;
        RECT 172.950 337.950 175.050 338.400 ;
        RECT 181.950 339.600 184.050 340.050 ;
        RECT 193.950 339.600 196.050 340.050 ;
        RECT 181.950 338.400 196.050 339.600 ;
        RECT 181.950 337.950 184.050 338.400 ;
        RECT 193.950 337.950 196.050 338.400 ;
        RECT 199.950 339.600 202.050 340.050 ;
        RECT 226.950 339.600 229.050 340.050 ;
        RECT 199.950 338.400 229.050 339.600 ;
        RECT 199.950 337.950 202.050 338.400 ;
        RECT 226.950 337.950 229.050 338.400 ;
        RECT 241.950 339.600 244.050 340.050 ;
        RECT 281.400 339.600 282.600 340.950 ;
        RECT 241.950 338.400 282.600 339.600 ;
        RECT 283.950 339.600 286.050 340.050 ;
        RECT 319.950 339.600 322.050 340.050 ;
        RECT 283.950 338.400 322.050 339.600 ;
        RECT 241.950 337.950 244.050 338.400 ;
        RECT 283.950 337.950 286.050 338.400 ;
        RECT 319.950 337.950 322.050 338.400 ;
        RECT 328.950 339.600 331.050 340.050 ;
        RECT 349.950 339.600 352.050 340.050 ;
        RECT 328.950 338.400 352.050 339.600 ;
        RECT 328.950 337.950 331.050 338.400 ;
        RECT 349.950 337.950 352.050 338.400 ;
        RECT 352.950 339.600 355.050 340.050 ;
        RECT 397.950 339.600 400.050 340.050 ;
        RECT 352.950 338.400 400.050 339.600 ;
        RECT 352.950 337.950 355.050 338.400 ;
        RECT 397.950 337.950 400.050 338.400 ;
        RECT 442.950 339.600 445.050 340.050 ;
        RECT 482.400 339.600 483.600 340.950 ;
        RECT 442.950 338.400 483.600 339.600 ;
        RECT 484.950 339.600 487.050 340.050 ;
        RECT 520.950 339.600 523.050 340.050 ;
        RECT 535.950 339.600 538.050 340.050 ;
        RECT 484.950 338.400 523.050 339.600 ;
        RECT 442.950 337.950 445.050 338.400 ;
        RECT 484.950 337.950 487.050 338.400 ;
        RECT 520.950 337.950 523.050 338.400 ;
        RECT 530.400 338.400 538.050 339.600 ;
        RECT 605.400 339.600 606.600 340.950 ;
        RECT 646.950 339.600 649.050 340.050 ;
        RECT 694.950 339.600 697.050 340.050 ;
        RECT 605.400 338.400 697.050 339.600 ;
        RECT 130.950 336.600 133.050 337.050 ;
        RECT 157.950 336.600 160.050 337.050 ;
        RECT 130.950 335.400 160.050 336.600 ;
        RECT 130.950 334.950 133.050 335.400 ;
        RECT 157.950 334.950 160.050 335.400 ;
        RECT 373.950 336.600 376.050 337.050 ;
        RECT 385.950 336.600 388.050 337.050 ;
        RECT 406.950 336.600 409.050 337.050 ;
        RECT 448.950 336.600 451.050 337.050 ;
        RECT 373.950 335.400 451.050 336.600 ;
        RECT 373.950 334.950 376.050 335.400 ;
        RECT 385.950 334.950 388.050 335.400 ;
        RECT 406.950 334.950 409.050 335.400 ;
        RECT 448.950 334.950 451.050 335.400 ;
        RECT 478.950 336.600 481.050 337.050 ;
        RECT 530.400 336.600 531.600 338.400 ;
        RECT 535.950 337.950 538.050 338.400 ;
        RECT 646.950 337.950 649.050 338.400 ;
        RECT 694.950 337.950 697.050 338.400 ;
        RECT 721.950 339.600 724.050 340.050 ;
        RECT 727.950 339.600 730.050 340.050 ;
        RECT 721.950 338.400 730.050 339.600 ;
        RECT 721.950 337.950 724.050 338.400 ;
        RECT 727.950 337.950 730.050 338.400 ;
        RECT 478.950 335.400 531.600 336.600 ;
        RECT 607.950 336.600 610.050 337.050 ;
        RECT 640.950 336.600 643.050 337.050 ;
        RECT 715.950 336.600 718.050 337.050 ;
        RECT 736.950 336.600 739.050 337.050 ;
        RECT 607.950 335.400 739.050 336.600 ;
        RECT 478.950 334.950 481.050 335.400 ;
        RECT 607.950 334.950 610.050 335.400 ;
        RECT 640.950 334.950 643.050 335.400 ;
        RECT 715.950 334.950 718.050 335.400 ;
        RECT 736.950 334.950 739.050 335.400 ;
        RECT 25.950 333.600 28.050 334.050 ;
        RECT 91.950 333.600 94.050 334.050 ;
        RECT 145.950 333.600 148.050 334.050 ;
        RECT 196.950 333.600 199.050 334.050 ;
        RECT 226.950 333.600 229.050 334.050 ;
        RECT 25.950 332.400 229.050 333.600 ;
        RECT 25.950 331.950 28.050 332.400 ;
        RECT 91.950 331.950 94.050 332.400 ;
        RECT 145.950 331.950 148.050 332.400 ;
        RECT 196.950 331.950 199.050 332.400 ;
        RECT 226.950 331.950 229.050 332.400 ;
        RECT 307.950 327.600 310.050 328.050 ;
        RECT 331.950 327.600 334.050 328.050 ;
        RECT 337.950 327.600 340.050 328.050 ;
        RECT 307.950 326.400 340.050 327.600 ;
        RECT 307.950 325.950 310.050 326.400 ;
        RECT 331.950 325.950 334.050 326.400 ;
        RECT 337.950 325.950 340.050 326.400 ;
        RECT 109.950 318.600 112.050 319.050 ;
        RECT 184.950 318.600 187.050 319.050 ;
        RECT 109.950 317.400 187.050 318.600 ;
        RECT 109.950 316.950 112.050 317.400 ;
        RECT 184.950 316.950 187.050 317.400 ;
        RECT 298.950 318.600 301.050 319.050 ;
        RECT 490.950 318.600 493.050 319.050 ;
        RECT 298.950 317.400 493.050 318.600 ;
        RECT 298.950 316.950 301.050 317.400 ;
        RECT 490.950 316.950 493.050 317.400 ;
        RECT 19.950 315.600 22.050 316.050 ;
        RECT 52.950 315.600 55.050 316.050 ;
        RECT 19.950 314.400 55.050 315.600 ;
        RECT 19.950 313.950 22.050 314.400 ;
        RECT 52.950 313.950 55.050 314.400 ;
        RECT 190.950 315.600 193.050 316.050 ;
        RECT 202.950 315.600 205.050 316.050 ;
        RECT 190.950 314.400 205.050 315.600 ;
        RECT 190.950 313.950 193.050 314.400 ;
        RECT 202.950 313.950 205.050 314.400 ;
        RECT 247.950 315.600 250.050 316.050 ;
        RECT 262.950 315.600 265.050 316.050 ;
        RECT 247.950 314.400 265.050 315.600 ;
        RECT 247.950 313.950 250.050 314.400 ;
        RECT 262.950 313.950 265.050 314.400 ;
        RECT 622.950 315.600 625.050 316.050 ;
        RECT 643.950 315.600 646.050 316.050 ;
        RECT 652.950 315.600 655.050 316.050 ;
        RECT 622.950 314.400 655.050 315.600 ;
        RECT 622.950 313.950 625.050 314.400 ;
        RECT 643.950 313.950 646.050 314.400 ;
        RECT 652.950 313.950 655.050 314.400 ;
        RECT 58.950 312.600 61.050 313.050 ;
        RECT 103.950 312.600 106.050 313.050 ;
        RECT 58.950 311.400 106.050 312.600 ;
        RECT 58.950 310.950 61.050 311.400 ;
        RECT 103.950 310.950 106.050 311.400 ;
        RECT 199.950 312.600 202.050 313.050 ;
        RECT 229.950 312.600 232.050 313.050 ;
        RECT 199.950 311.400 232.050 312.600 ;
        RECT 199.950 310.950 202.050 311.400 ;
        RECT 229.950 310.950 232.050 311.400 ;
        RECT 283.950 312.600 286.050 313.050 ;
        RECT 298.950 312.600 301.050 313.050 ;
        RECT 283.950 311.400 301.050 312.600 ;
        RECT 283.950 310.950 286.050 311.400 ;
        RECT 298.950 310.950 301.050 311.400 ;
        RECT 304.950 312.600 307.050 313.050 ;
        RECT 310.950 312.600 313.050 313.050 ;
        RECT 304.950 311.400 313.050 312.600 ;
        RECT 304.950 310.950 307.050 311.400 ;
        RECT 310.950 310.950 313.050 311.400 ;
        RECT 379.950 312.600 382.050 313.050 ;
        RECT 424.950 312.600 427.050 313.050 ;
        RECT 478.950 312.600 481.050 313.050 ;
        RECT 379.950 311.400 423.600 312.600 ;
        RECT 379.950 310.950 382.050 311.400 ;
        RECT 422.400 310.050 423.600 311.400 ;
        RECT 424.950 311.400 481.050 312.600 ;
        RECT 424.950 310.950 427.050 311.400 ;
        RECT 478.950 310.950 481.050 311.400 ;
        RECT 541.950 312.600 544.050 313.050 ;
        RECT 586.950 312.600 589.050 313.050 ;
        RECT 541.950 311.400 589.050 312.600 ;
        RECT 541.950 310.950 544.050 311.400 ;
        RECT 586.950 310.950 589.050 311.400 ;
        RECT 40.950 309.600 43.050 310.050 ;
        RECT 82.950 309.600 85.050 310.050 ;
        RECT 40.950 308.400 85.050 309.600 ;
        RECT 40.950 307.950 43.050 308.400 ;
        RECT 82.950 307.950 85.050 308.400 ;
        RECT 88.950 309.600 91.050 310.050 ;
        RECT 106.950 309.600 109.050 310.050 ;
        RECT 88.950 308.400 109.050 309.600 ;
        RECT 88.950 307.950 91.050 308.400 ;
        RECT 106.950 307.950 109.050 308.400 ;
        RECT 181.950 309.600 184.050 310.050 ;
        RECT 193.950 309.600 196.050 310.050 ;
        RECT 181.950 308.400 196.050 309.600 ;
        RECT 181.950 307.950 184.050 308.400 ;
        RECT 193.950 307.950 196.050 308.400 ;
        RECT 202.950 309.600 205.050 310.050 ;
        RECT 232.950 309.600 235.050 310.050 ;
        RECT 256.950 309.600 259.050 310.050 ;
        RECT 310.950 309.600 313.050 310.050 ;
        RECT 202.950 308.400 313.050 309.600 ;
        RECT 202.950 307.950 205.050 308.400 ;
        RECT 232.950 307.950 235.050 308.400 ;
        RECT 256.950 307.950 259.050 308.400 ;
        RECT 310.950 307.950 313.050 308.400 ;
        RECT 328.950 309.600 331.050 310.050 ;
        RECT 340.950 309.600 343.050 310.050 ;
        RECT 328.950 308.400 343.050 309.600 ;
        RECT 328.950 307.950 331.050 308.400 ;
        RECT 340.950 307.950 343.050 308.400 ;
        RECT 382.950 307.950 385.050 310.050 ;
        RECT 415.950 307.950 418.050 310.050 ;
        RECT 421.950 307.950 424.050 310.050 ;
        RECT 640.950 309.600 643.050 310.050 ;
        RECT 655.950 309.600 658.050 310.050 ;
        RECT 640.950 308.400 658.050 309.600 ;
        RECT 640.950 307.950 643.050 308.400 ;
        RECT 655.950 307.950 658.050 308.400 ;
        RECT 187.950 306.600 190.050 307.050 ;
        RECT 199.950 306.600 202.050 307.050 ;
        RECT 187.950 305.400 202.050 306.600 ;
        RECT 187.950 304.950 190.050 305.400 ;
        RECT 199.950 304.950 202.050 305.400 ;
        RECT 322.950 306.600 325.050 307.050 ;
        RECT 376.950 306.600 379.050 307.050 ;
        RECT 322.950 305.400 379.050 306.600 ;
        RECT 322.950 304.950 325.050 305.400 ;
        RECT 376.950 304.950 379.050 305.400 ;
        RECT 379.950 306.600 382.050 307.050 ;
        RECT 383.400 306.600 384.600 307.950 ;
        RECT 379.950 305.400 384.600 306.600 ;
        RECT 416.400 306.600 417.600 307.950 ;
        RECT 418.950 306.600 421.050 307.050 ;
        RECT 416.400 305.400 421.050 306.600 ;
        RECT 379.950 304.950 382.050 305.400 ;
        RECT 418.950 304.950 421.050 305.400 ;
        RECT 574.950 306.600 577.050 307.050 ;
        RECT 586.950 306.600 589.050 307.050 ;
        RECT 574.950 305.400 589.050 306.600 ;
        RECT 574.950 304.950 577.050 305.400 ;
        RECT 586.950 304.950 589.050 305.400 ;
        RECT 613.950 306.600 616.050 307.050 ;
        RECT 649.950 306.600 652.050 307.050 ;
        RECT 613.950 305.400 652.050 306.600 ;
        RECT 613.950 304.950 616.050 305.400 ;
        RECT 649.950 304.950 652.050 305.400 ;
        RECT 238.950 303.600 241.050 304.050 ;
        RECT 514.950 303.600 517.050 304.050 ;
        RECT 541.950 303.600 544.050 304.050 ;
        RECT 688.950 303.600 691.050 304.050 ;
        RECT 724.950 303.600 727.050 304.050 ;
        RECT 238.950 302.400 727.050 303.600 ;
        RECT 238.950 301.950 241.050 302.400 ;
        RECT 514.950 301.950 517.050 302.400 ;
        RECT 541.950 301.950 544.050 302.400 ;
        RECT 688.950 301.950 691.050 302.400 ;
        RECT 724.950 301.950 727.050 302.400 ;
        RECT 535.950 300.600 538.050 301.050 ;
        RECT 580.950 300.600 583.050 301.050 ;
        RECT 535.950 299.400 583.050 300.600 ;
        RECT 535.950 298.950 538.050 299.400 ;
        RECT 580.950 298.950 583.050 299.400 ;
        RECT 31.950 294.600 34.050 295.050 ;
        RECT 43.950 294.600 46.050 295.050 ;
        RECT 31.950 293.400 46.050 294.600 ;
        RECT 31.950 292.950 34.050 293.400 ;
        RECT 43.950 292.950 46.050 293.400 ;
        RECT 40.950 279.600 43.050 280.050 ;
        RECT 46.950 279.600 49.050 280.050 ;
        RECT 40.950 278.400 49.050 279.600 ;
        RECT 40.950 277.950 43.050 278.400 ;
        RECT 46.950 277.950 49.050 278.400 ;
        RECT 142.950 276.600 145.050 277.050 ;
        RECT 214.950 276.600 217.050 277.050 ;
        RECT 142.950 275.400 217.050 276.600 ;
        RECT 142.950 274.950 145.050 275.400 ;
        RECT 214.950 274.950 217.050 275.400 ;
        RECT 310.950 276.600 313.050 277.050 ;
        RECT 358.950 276.600 361.050 277.050 ;
        RECT 310.950 275.400 361.050 276.600 ;
        RECT 310.950 274.950 313.050 275.400 ;
        RECT 358.950 274.950 361.050 275.400 ;
        RECT 436.950 276.600 439.050 277.050 ;
        RECT 448.950 276.600 451.050 277.050 ;
        RECT 436.950 275.400 451.050 276.600 ;
        RECT 436.950 274.950 439.050 275.400 ;
        RECT 448.950 274.950 451.050 275.400 ;
        RECT 34.950 273.600 37.050 274.050 ;
        RECT 73.950 273.600 76.050 274.050 ;
        RECT 181.950 273.600 184.050 274.050 ;
        RECT 187.950 273.600 190.050 274.050 ;
        RECT 34.950 272.400 45.600 273.600 ;
        RECT 34.950 271.950 37.050 272.400 ;
        RECT 40.950 268.950 43.050 271.050 ;
        RECT 44.400 270.600 45.600 272.400 ;
        RECT 73.950 272.400 190.050 273.600 ;
        RECT 73.950 271.950 76.050 272.400 ;
        RECT 181.950 271.950 184.050 272.400 ;
        RECT 187.950 271.950 190.050 272.400 ;
        RECT 355.950 273.600 358.050 274.050 ;
        RECT 391.950 273.600 394.050 274.050 ;
        RECT 427.950 273.600 430.050 274.050 ;
        RECT 355.950 272.400 430.050 273.600 ;
        RECT 355.950 271.950 358.050 272.400 ;
        RECT 391.950 271.950 394.050 272.400 ;
        RECT 427.950 271.950 430.050 272.400 ;
        RECT 502.950 273.600 505.050 274.050 ;
        RECT 529.950 273.600 532.050 274.050 ;
        RECT 502.950 272.400 532.050 273.600 ;
        RECT 502.950 271.950 505.050 272.400 ;
        RECT 529.950 271.950 532.050 272.400 ;
        RECT 601.950 273.600 604.050 274.050 ;
        RECT 610.950 273.600 613.050 274.050 ;
        RECT 601.950 272.400 613.050 273.600 ;
        RECT 601.950 271.950 604.050 272.400 ;
        RECT 610.950 271.950 613.050 272.400 ;
        RECT 79.950 270.600 82.050 271.050 ;
        RECT 91.950 270.600 94.050 271.050 ;
        RECT 44.400 269.400 75.600 270.600 ;
        RECT 16.950 267.600 19.050 268.050 ;
        RECT 31.950 267.600 34.050 268.050 ;
        RECT 16.950 266.400 34.050 267.600 ;
        RECT 16.950 265.950 19.050 266.400 ;
        RECT 31.950 265.950 34.050 266.400 ;
        RECT 41.400 261.600 42.600 268.950 ;
        RECT 43.950 267.600 46.050 268.050 ;
        RECT 70.950 267.600 73.050 268.050 ;
        RECT 43.950 266.400 73.050 267.600 ;
        RECT 74.400 267.600 75.600 269.400 ;
        RECT 79.950 269.400 94.050 270.600 ;
        RECT 79.950 268.950 82.050 269.400 ;
        RECT 91.950 268.950 94.050 269.400 ;
        RECT 268.950 268.950 271.050 271.050 ;
        RECT 349.950 268.950 352.050 271.050 ;
        RECT 379.950 270.600 382.050 271.050 ;
        RECT 388.950 270.600 391.050 271.050 ;
        RECT 379.950 269.400 391.050 270.600 ;
        RECT 379.950 268.950 382.050 269.400 ;
        RECT 388.950 268.950 391.050 269.400 ;
        RECT 592.950 270.600 595.050 271.050 ;
        RECT 637.950 270.600 640.050 271.050 ;
        RECT 655.950 270.600 658.050 271.050 ;
        RECT 592.950 269.400 658.050 270.600 ;
        RECT 592.950 268.950 595.050 269.400 ;
        RECT 637.950 268.950 640.050 269.400 ;
        RECT 655.950 268.950 658.050 269.400 ;
        RECT 76.950 267.600 79.050 268.050 ;
        RECT 74.400 266.400 79.050 267.600 ;
        RECT 43.950 265.950 46.050 266.400 ;
        RECT 70.950 265.950 73.050 266.400 ;
        RECT 76.950 265.950 79.050 266.400 ;
        RECT 136.950 267.600 139.050 268.050 ;
        RECT 151.950 267.600 154.050 268.050 ;
        RECT 184.950 267.600 187.050 268.050 ;
        RECT 136.950 266.400 187.050 267.600 ;
        RECT 136.950 265.950 139.050 266.400 ;
        RECT 151.950 265.950 154.050 266.400 ;
        RECT 184.950 265.950 187.050 266.400 ;
        RECT 229.950 267.600 232.050 268.050 ;
        RECT 247.950 267.600 250.050 268.050 ;
        RECT 229.950 266.400 250.050 267.600 ;
        RECT 269.400 267.600 270.600 268.950 ;
        RECT 307.950 267.600 310.050 268.050 ;
        RECT 269.400 266.400 310.050 267.600 ;
        RECT 229.950 265.950 232.050 266.400 ;
        RECT 247.950 265.950 250.050 266.400 ;
        RECT 307.950 265.950 310.050 266.400 ;
        RECT 350.400 265.050 351.600 268.950 ;
        RECT 454.950 267.600 457.050 268.050 ;
        RECT 499.950 267.600 502.050 268.050 ;
        RECT 454.950 266.400 502.050 267.600 ;
        RECT 454.950 265.950 457.050 266.400 ;
        RECT 499.950 265.950 502.050 266.400 ;
        RECT 550.950 267.600 553.050 268.050 ;
        RECT 556.950 267.600 559.050 268.050 ;
        RECT 550.950 266.400 559.050 267.600 ;
        RECT 550.950 265.950 553.050 266.400 ;
        RECT 556.950 265.950 559.050 266.400 ;
        RECT 73.950 264.600 76.050 265.050 ;
        RECT 112.950 264.600 115.050 265.050 ;
        RECT 73.950 263.400 115.050 264.600 ;
        RECT 73.950 262.950 76.050 263.400 ;
        RECT 112.950 262.950 115.050 263.400 ;
        RECT 118.950 264.600 121.050 265.050 ;
        RECT 256.950 264.600 259.050 265.050 ;
        RECT 265.950 264.600 268.050 265.050 ;
        RECT 118.950 263.400 268.050 264.600 ;
        RECT 118.950 262.950 121.050 263.400 ;
        RECT 256.950 262.950 259.050 263.400 ;
        RECT 265.950 262.950 268.050 263.400 ;
        RECT 349.950 262.950 352.050 265.050 ;
        RECT 352.950 264.600 355.050 265.050 ;
        RECT 358.950 264.600 361.050 265.050 ;
        RECT 352.950 263.400 361.050 264.600 ;
        RECT 352.950 262.950 355.050 263.400 ;
        RECT 358.950 262.950 361.050 263.400 ;
        RECT 478.950 264.600 481.050 265.050 ;
        RECT 508.950 264.600 511.050 265.050 ;
        RECT 478.950 263.400 511.050 264.600 ;
        RECT 478.950 262.950 481.050 263.400 ;
        RECT 508.950 262.950 511.050 263.400 ;
        RECT 532.950 264.600 535.050 265.050 ;
        RECT 571.950 264.600 574.050 265.050 ;
        RECT 532.950 263.400 574.050 264.600 ;
        RECT 532.950 262.950 535.050 263.400 ;
        RECT 571.950 262.950 574.050 263.400 ;
        RECT 694.950 264.600 697.050 265.050 ;
        RECT 697.950 264.600 700.050 265.050 ;
        RECT 760.950 264.600 763.050 265.050 ;
        RECT 694.950 263.400 763.050 264.600 ;
        RECT 694.950 262.950 697.050 263.400 ;
        RECT 697.950 262.950 700.050 263.400 ;
        RECT 760.950 262.950 763.050 263.400 ;
        RECT 115.950 261.600 118.050 262.050 ;
        RECT 41.400 260.400 118.050 261.600 ;
        RECT 115.950 259.950 118.050 260.400 ;
        RECT 133.950 261.600 136.050 262.050 ;
        RECT 184.950 261.600 187.050 262.050 ;
        RECT 133.950 260.400 187.050 261.600 ;
        RECT 133.950 259.950 136.050 260.400 ;
        RECT 184.950 259.950 187.050 260.400 ;
        RECT 211.950 261.600 214.050 262.050 ;
        RECT 271.950 261.600 274.050 262.050 ;
        RECT 211.950 260.400 274.050 261.600 ;
        RECT 211.950 259.950 214.050 260.400 ;
        RECT 271.950 259.950 274.050 260.400 ;
        RECT 457.950 261.600 460.050 262.050 ;
        RECT 478.950 261.600 481.050 262.050 ;
        RECT 457.950 260.400 481.050 261.600 ;
        RECT 457.950 259.950 460.050 260.400 ;
        RECT 478.950 259.950 481.050 260.400 ;
        RECT 526.950 261.600 529.050 262.050 ;
        RECT 547.950 261.600 550.050 262.050 ;
        RECT 562.950 261.600 565.050 262.050 ;
        RECT 526.950 260.400 565.050 261.600 ;
        RECT 526.950 259.950 529.050 260.400 ;
        RECT 547.950 259.950 550.050 260.400 ;
        RECT 562.950 259.950 565.050 260.400 ;
        RECT 658.950 261.600 661.050 262.050 ;
        RECT 661.950 261.600 664.050 262.050 ;
        RECT 709.950 261.600 712.050 262.050 ;
        RECT 733.950 261.600 736.050 262.050 ;
        RECT 658.950 260.400 736.050 261.600 ;
        RECT 658.950 259.950 661.050 260.400 ;
        RECT 661.950 259.950 664.050 260.400 ;
        RECT 709.950 259.950 712.050 260.400 ;
        RECT 733.950 259.950 736.050 260.400 ;
        RECT 229.950 258.600 232.050 259.050 ;
        RECT 493.950 258.600 496.050 259.050 ;
        RECT 229.950 257.400 496.050 258.600 ;
        RECT 229.950 256.950 232.050 257.400 ;
        RECT 493.950 256.950 496.050 257.400 ;
        RECT 580.950 258.600 583.050 259.050 ;
        RECT 679.950 258.600 682.050 259.050 ;
        RECT 580.950 257.400 682.050 258.600 ;
        RECT 580.950 256.950 583.050 257.400 ;
        RECT 679.950 256.950 682.050 257.400 ;
        RECT 313.950 255.600 316.050 256.050 ;
        RECT 556.950 255.600 559.050 256.050 ;
        RECT 313.950 254.400 559.050 255.600 ;
        RECT 313.950 253.950 316.050 254.400 ;
        RECT 556.950 253.950 559.050 254.400 ;
        RECT 487.950 252.600 490.050 253.050 ;
        RECT 493.950 252.600 496.050 253.050 ;
        RECT 487.950 251.400 496.050 252.600 ;
        RECT 487.950 250.950 490.050 251.400 ;
        RECT 493.950 250.950 496.050 251.400 ;
        RECT 583.950 252.600 586.050 253.050 ;
        RECT 613.950 252.600 616.050 253.050 ;
        RECT 583.950 251.400 616.050 252.600 ;
        RECT 583.950 250.950 586.050 251.400 ;
        RECT 613.950 250.950 616.050 251.400 ;
        RECT 568.950 249.600 571.050 250.050 ;
        RECT 613.950 249.600 616.050 250.050 ;
        RECT 568.950 248.400 616.050 249.600 ;
        RECT 568.950 247.950 571.050 248.400 ;
        RECT 613.950 247.950 616.050 248.400 ;
        RECT 181.950 246.600 184.050 247.050 ;
        RECT 190.950 246.600 193.050 247.050 ;
        RECT 181.950 245.400 193.050 246.600 ;
        RECT 181.950 244.950 184.050 245.400 ;
        RECT 190.950 244.950 193.050 245.400 ;
        RECT 385.950 246.600 388.050 247.050 ;
        RECT 430.950 246.600 433.050 247.050 ;
        RECT 385.950 245.400 433.050 246.600 ;
        RECT 385.950 244.950 388.050 245.400 ;
        RECT 430.950 244.950 433.050 245.400 ;
        RECT 547.950 246.600 550.050 247.050 ;
        RECT 694.950 246.600 697.050 247.050 ;
        RECT 547.950 245.400 697.050 246.600 ;
        RECT 547.950 244.950 550.050 245.400 ;
        RECT 694.950 244.950 697.050 245.400 ;
        RECT 187.950 241.950 190.050 244.050 ;
        RECT 346.950 243.600 349.050 244.050 ;
        RECT 364.950 243.600 367.050 244.050 ;
        RECT 346.950 242.400 367.050 243.600 ;
        RECT 346.950 241.950 349.050 242.400 ;
        RECT 364.950 241.950 367.050 242.400 ;
        RECT 370.950 243.600 373.050 244.050 ;
        RECT 445.950 243.600 448.050 244.050 ;
        RECT 448.950 243.600 451.050 244.050 ;
        RECT 526.950 243.600 529.050 244.050 ;
        RECT 370.950 242.400 529.050 243.600 ;
        RECT 370.950 241.950 373.050 242.400 ;
        RECT 445.950 241.950 448.050 242.400 ;
        RECT 448.950 241.950 451.050 242.400 ;
        RECT 526.950 241.950 529.050 242.400 ;
        RECT 553.950 243.600 556.050 244.050 ;
        RECT 577.950 243.600 580.050 244.050 ;
        RECT 553.950 242.400 580.050 243.600 ;
        RECT 553.950 241.950 556.050 242.400 ;
        RECT 577.950 241.950 580.050 242.400 ;
        RECT 619.950 243.600 622.050 244.050 ;
        RECT 652.950 243.600 655.050 244.050 ;
        RECT 619.950 242.400 655.050 243.600 ;
        RECT 619.950 241.950 622.050 242.400 ;
        RECT 652.950 241.950 655.050 242.400 ;
        RECT 64.950 240.600 67.050 241.050 ;
        RECT 70.950 240.600 73.050 241.050 ;
        RECT 64.950 239.400 73.050 240.600 ;
        RECT 64.950 238.950 67.050 239.400 ;
        RECT 70.950 238.950 73.050 239.400 ;
        RECT 76.950 240.600 79.050 241.050 ;
        RECT 79.950 240.600 82.050 241.050 ;
        RECT 139.950 240.600 142.050 241.050 ;
        RECT 76.950 239.400 142.050 240.600 ;
        RECT 76.950 238.950 79.050 239.400 ;
        RECT 79.950 238.950 82.050 239.400 ;
        RECT 139.950 238.950 142.050 239.400 ;
        RECT 188.400 238.050 189.600 241.950 ;
        RECT 217.950 240.600 220.050 241.050 ;
        RECT 223.950 240.600 226.050 241.050 ;
        RECT 217.950 239.400 226.050 240.600 ;
        RECT 217.950 238.950 220.050 239.400 ;
        RECT 223.950 238.950 226.050 239.400 ;
        RECT 409.950 240.600 412.050 241.050 ;
        RECT 439.950 240.600 442.050 241.050 ;
        RECT 409.950 239.400 442.050 240.600 ;
        RECT 409.950 238.950 412.050 239.400 ;
        RECT 439.950 238.950 442.050 239.400 ;
        RECT 532.950 240.600 535.050 241.050 ;
        RECT 685.950 240.600 688.050 241.050 ;
        RECT 703.950 240.600 706.050 241.050 ;
        RECT 532.950 239.400 576.600 240.600 ;
        RECT 532.950 238.950 535.050 239.400 ;
        RECT 575.400 238.050 576.600 239.400 ;
        RECT 685.950 239.400 706.050 240.600 ;
        RECT 685.950 238.950 688.050 239.400 ;
        RECT 703.950 238.950 706.050 239.400 ;
        RECT 724.950 240.600 727.050 241.050 ;
        RECT 736.950 240.600 739.050 241.050 ;
        RECT 724.950 239.400 739.050 240.600 ;
        RECT 724.950 238.950 727.050 239.400 ;
        RECT 736.950 238.950 739.050 239.400 ;
        RECT 115.950 237.600 118.050 238.050 ;
        RECT 145.950 237.600 148.050 238.050 ;
        RECT 115.950 236.400 148.050 237.600 ;
        RECT 115.950 235.950 118.050 236.400 ;
        RECT 145.950 235.950 148.050 236.400 ;
        RECT 187.950 235.950 190.050 238.050 ;
        RECT 343.950 237.600 346.050 238.050 ;
        RECT 346.950 237.600 349.050 238.050 ;
        RECT 367.950 237.600 370.050 238.050 ;
        RECT 343.950 236.400 370.050 237.600 ;
        RECT 343.950 235.950 346.050 236.400 ;
        RECT 346.950 235.950 349.050 236.400 ;
        RECT 367.950 235.950 370.050 236.400 ;
        RECT 574.950 235.950 577.050 238.050 ;
        RECT 622.950 237.600 625.050 238.050 ;
        RECT 655.950 237.600 658.050 238.050 ;
        RECT 622.950 236.400 658.050 237.600 ;
        RECT 622.950 235.950 625.050 236.400 ;
        RECT 655.950 235.950 658.050 236.400 ;
        RECT 37.950 234.600 40.050 235.050 ;
        RECT 79.950 234.600 82.050 235.050 ;
        RECT 37.950 233.400 82.050 234.600 ;
        RECT 37.950 232.950 40.050 233.400 ;
        RECT 79.950 232.950 82.050 233.400 ;
        RECT 148.950 234.600 151.050 235.050 ;
        RECT 163.950 234.600 166.050 235.050 ;
        RECT 148.950 233.400 166.050 234.600 ;
        RECT 148.950 232.950 151.050 233.400 ;
        RECT 163.950 232.950 166.050 233.400 ;
        RECT 349.950 234.600 352.050 235.050 ;
        RECT 367.950 234.600 370.050 235.050 ;
        RECT 349.950 233.400 370.050 234.600 ;
        RECT 349.950 232.950 352.050 233.400 ;
        RECT 367.950 232.950 370.050 233.400 ;
        RECT 403.950 234.600 406.050 235.050 ;
        RECT 421.950 234.600 424.050 235.050 ;
        RECT 403.950 233.400 424.050 234.600 ;
        RECT 403.950 232.950 406.050 233.400 ;
        RECT 421.950 232.950 424.050 233.400 ;
        RECT 457.950 234.600 460.050 235.050 ;
        RECT 490.950 234.600 493.050 235.050 ;
        RECT 457.950 233.400 493.050 234.600 ;
        RECT 457.950 232.950 460.050 233.400 ;
        RECT 490.950 232.950 493.050 233.400 ;
        RECT 496.950 234.600 499.050 235.050 ;
        RECT 508.950 234.600 511.050 235.050 ;
        RECT 496.950 233.400 511.050 234.600 ;
        RECT 496.950 232.950 499.050 233.400 ;
        RECT 508.950 232.950 511.050 233.400 ;
        RECT 31.950 231.600 34.050 232.050 ;
        RECT 64.950 231.600 67.050 232.050 ;
        RECT 31.950 230.400 67.050 231.600 ;
        RECT 31.950 229.950 34.050 230.400 ;
        RECT 64.950 229.950 67.050 230.400 ;
        RECT 415.950 231.600 418.050 232.050 ;
        RECT 496.950 231.600 499.050 232.050 ;
        RECT 415.950 230.400 499.050 231.600 ;
        RECT 415.950 229.950 418.050 230.400 ;
        RECT 496.950 229.950 499.050 230.400 ;
        RECT 100.950 207.600 103.050 208.050 ;
        RECT 106.950 207.600 109.050 208.050 ;
        RECT 100.950 206.400 109.050 207.600 ;
        RECT 100.950 205.950 103.050 206.400 ;
        RECT 106.950 205.950 109.050 206.400 ;
        RECT 115.950 207.600 118.050 208.050 ;
        RECT 121.950 207.600 124.050 208.050 ;
        RECT 226.950 207.600 229.050 208.050 ;
        RECT 115.950 206.400 229.050 207.600 ;
        RECT 115.950 205.950 118.050 206.400 ;
        RECT 121.950 205.950 124.050 206.400 ;
        RECT 226.950 205.950 229.050 206.400 ;
        RECT 118.950 204.600 121.050 205.050 ;
        RECT 142.950 204.600 145.050 205.050 ;
        RECT 145.950 204.600 148.050 205.050 ;
        RECT 118.950 203.400 148.050 204.600 ;
        RECT 118.950 202.950 121.050 203.400 ;
        RECT 142.950 202.950 145.050 203.400 ;
        RECT 145.950 202.950 148.050 203.400 ;
        RECT 220.950 204.600 223.050 205.050 ;
        RECT 229.950 204.600 232.050 205.050 ;
        RECT 220.950 203.400 232.050 204.600 ;
        RECT 220.950 202.950 223.050 203.400 ;
        RECT 229.950 202.950 232.050 203.400 ;
        RECT 691.950 204.600 694.050 205.050 ;
        RECT 754.950 204.600 757.050 205.050 ;
        RECT 691.950 203.400 757.050 204.600 ;
        RECT 691.950 202.950 694.050 203.400 ;
        RECT 754.950 202.950 757.050 203.400 ;
        RECT 139.950 201.600 142.050 202.050 ;
        RECT 151.950 201.600 154.050 202.050 ;
        RECT 139.950 200.400 154.050 201.600 ;
        RECT 139.950 199.950 142.050 200.400 ;
        RECT 151.950 199.950 154.050 200.400 ;
        RECT 199.950 201.600 202.050 202.050 ;
        RECT 226.950 201.600 229.050 202.050 ;
        RECT 199.950 200.400 229.050 201.600 ;
        RECT 199.950 199.950 202.050 200.400 ;
        RECT 226.950 199.950 229.050 200.400 ;
        RECT 250.950 201.600 253.050 202.050 ;
        RECT 265.950 201.600 268.050 202.050 ;
        RECT 250.950 200.400 268.050 201.600 ;
        RECT 250.950 199.950 253.050 200.400 ;
        RECT 265.950 199.950 268.050 200.400 ;
        RECT 373.950 201.600 376.050 202.050 ;
        RECT 547.950 201.600 550.050 202.050 ;
        RECT 568.950 201.600 571.050 202.050 ;
        RECT 373.950 200.400 571.050 201.600 ;
        RECT 373.950 199.950 376.050 200.400 ;
        RECT 547.950 199.950 550.050 200.400 ;
        RECT 568.950 199.950 571.050 200.400 ;
        RECT 649.950 201.600 652.050 202.050 ;
        RECT 685.950 201.600 688.050 202.050 ;
        RECT 649.950 200.400 688.050 201.600 ;
        RECT 649.950 199.950 652.050 200.400 ;
        RECT 685.950 199.950 688.050 200.400 ;
        RECT 730.950 199.950 733.050 202.050 ;
        RECT 97.950 198.600 100.050 199.050 ;
        RECT 106.950 198.600 109.050 199.050 ;
        RECT 97.950 197.400 109.050 198.600 ;
        RECT 97.950 196.950 100.050 197.400 ;
        RECT 106.950 196.950 109.050 197.400 ;
        RECT 217.950 198.600 220.050 199.050 ;
        RECT 223.950 198.600 226.050 199.050 ;
        RECT 217.950 197.400 226.050 198.600 ;
        RECT 217.950 196.950 220.050 197.400 ;
        RECT 223.950 196.950 226.050 197.400 ;
        RECT 478.950 198.600 481.050 199.050 ;
        RECT 496.950 198.600 499.050 199.050 ;
        RECT 478.950 197.400 499.050 198.600 ;
        RECT 478.950 196.950 481.050 197.400 ;
        RECT 496.950 196.950 499.050 197.400 ;
        RECT 526.950 198.600 529.050 199.050 ;
        RECT 532.950 198.600 535.050 199.050 ;
        RECT 526.950 197.400 535.050 198.600 ;
        RECT 526.950 196.950 529.050 197.400 ;
        RECT 532.950 196.950 535.050 197.400 ;
        RECT 538.950 198.600 541.050 199.050 ;
        RECT 553.950 198.600 556.050 199.050 ;
        RECT 538.950 197.400 556.050 198.600 ;
        RECT 538.950 196.950 541.050 197.400 ;
        RECT 553.950 196.950 556.050 197.400 ;
        RECT 556.950 198.600 559.050 199.050 ;
        RECT 724.950 198.600 727.050 199.050 ;
        RECT 556.950 197.400 727.050 198.600 ;
        RECT 556.950 196.950 559.050 197.400 ;
        RECT 724.950 196.950 727.050 197.400 ;
        RECT 34.950 195.600 37.050 196.050 ;
        RECT 40.950 195.600 43.050 196.050 ;
        RECT 46.950 195.600 49.050 196.050 ;
        RECT 34.950 194.400 49.050 195.600 ;
        RECT 34.950 193.950 37.050 194.400 ;
        RECT 40.950 193.950 43.050 194.400 ;
        RECT 46.950 193.950 49.050 194.400 ;
        RECT 100.950 195.600 103.050 196.050 ;
        RECT 109.950 195.600 112.050 196.050 ;
        RECT 100.950 194.400 112.050 195.600 ;
        RECT 100.950 193.950 103.050 194.400 ;
        RECT 109.950 193.950 112.050 194.400 ;
        RECT 148.950 195.600 151.050 196.050 ;
        RECT 184.950 195.600 187.050 196.050 ;
        RECT 148.950 194.400 187.050 195.600 ;
        RECT 148.950 193.950 151.050 194.400 ;
        RECT 184.950 193.950 187.050 194.400 ;
        RECT 193.950 195.600 196.050 196.050 ;
        RECT 262.950 195.600 265.050 196.050 ;
        RECT 193.950 194.400 265.050 195.600 ;
        RECT 193.950 193.950 196.050 194.400 ;
        RECT 262.950 193.950 265.050 194.400 ;
        RECT 463.950 195.600 466.050 196.050 ;
        RECT 490.950 195.600 493.050 196.050 ;
        RECT 463.950 194.400 493.050 195.600 ;
        RECT 463.950 193.950 466.050 194.400 ;
        RECT 490.950 193.950 493.050 194.400 ;
        RECT 541.950 195.600 544.050 196.050 ;
        RECT 557.400 195.600 558.600 196.950 ;
        RECT 731.400 196.050 732.600 199.950 ;
        RECT 616.950 195.600 619.050 196.050 ;
        RECT 541.950 194.400 558.600 195.600 ;
        RECT 605.400 194.400 619.050 195.600 ;
        RECT 541.950 193.950 544.050 194.400 ;
        RECT 31.950 192.600 34.050 193.050 ;
        RECT 73.950 192.600 76.050 193.050 ;
        RECT 97.950 192.600 100.050 193.050 ;
        RECT 31.950 191.400 100.050 192.600 ;
        RECT 31.950 190.950 34.050 191.400 ;
        RECT 73.950 190.950 76.050 191.400 ;
        RECT 97.950 190.950 100.050 191.400 ;
        RECT 142.950 192.600 145.050 193.050 ;
        RECT 190.950 192.600 193.050 193.050 ;
        RECT 142.950 191.400 193.050 192.600 ;
        RECT 142.950 190.950 145.050 191.400 ;
        RECT 190.950 190.950 193.050 191.400 ;
        RECT 307.950 192.600 310.050 193.050 ;
        RECT 316.950 192.600 319.050 193.050 ;
        RECT 415.950 192.600 418.050 193.050 ;
        RECT 307.950 191.400 418.050 192.600 ;
        RECT 307.950 190.950 310.050 191.400 ;
        RECT 316.950 190.950 319.050 191.400 ;
        RECT 415.950 190.950 418.050 191.400 ;
        RECT 535.950 192.600 538.050 193.050 ;
        RECT 605.400 192.600 606.600 194.400 ;
        RECT 616.950 193.950 619.050 194.400 ;
        RECT 640.950 195.600 643.050 196.050 ;
        RECT 697.950 195.600 700.050 196.050 ;
        RECT 640.950 194.400 700.050 195.600 ;
        RECT 640.950 193.950 643.050 194.400 ;
        RECT 697.950 193.950 700.050 194.400 ;
        RECT 730.950 193.950 733.050 196.050 ;
        RECT 535.950 191.400 606.600 192.600 ;
        RECT 607.950 192.600 610.050 193.050 ;
        RECT 622.950 192.600 625.050 193.050 ;
        RECT 643.950 192.600 646.050 193.050 ;
        RECT 607.950 191.400 646.050 192.600 ;
        RECT 535.950 190.950 538.050 191.400 ;
        RECT 607.950 190.950 610.050 191.400 ;
        RECT 622.950 190.950 625.050 191.400 ;
        RECT 643.950 190.950 646.050 191.400 ;
        RECT 688.950 192.600 691.050 193.050 ;
        RECT 721.950 192.600 724.050 193.050 ;
        RECT 733.950 192.600 736.050 193.050 ;
        RECT 688.950 191.400 736.050 192.600 ;
        RECT 688.950 190.950 691.050 191.400 ;
        RECT 721.950 190.950 724.050 191.400 ;
        RECT 733.950 190.950 736.050 191.400 ;
        RECT 31.950 189.600 34.050 190.050 ;
        RECT 67.950 189.600 70.050 190.050 ;
        RECT 103.950 189.600 106.050 190.050 ;
        RECT 31.950 188.400 106.050 189.600 ;
        RECT 31.950 187.950 34.050 188.400 ;
        RECT 67.950 187.950 70.050 188.400 ;
        RECT 103.950 187.950 106.050 188.400 ;
        RECT 304.950 189.600 307.050 190.050 ;
        RECT 343.950 189.600 346.050 190.050 ;
        RECT 526.950 189.600 529.050 190.050 ;
        RECT 304.950 188.400 529.050 189.600 ;
        RECT 304.950 187.950 307.050 188.400 ;
        RECT 343.950 187.950 346.050 188.400 ;
        RECT 526.950 187.950 529.050 188.400 ;
        RECT 565.950 189.600 568.050 190.050 ;
        RECT 601.950 189.600 604.050 190.050 ;
        RECT 565.950 188.400 604.050 189.600 ;
        RECT 565.950 187.950 568.050 188.400 ;
        RECT 601.950 187.950 604.050 188.400 ;
        RECT 64.950 186.600 67.050 187.050 ;
        RECT 73.950 186.600 76.050 187.050 ;
        RECT 64.950 185.400 76.050 186.600 ;
        RECT 64.950 184.950 67.050 185.400 ;
        RECT 73.950 184.950 76.050 185.400 ;
        RECT 157.950 180.600 160.050 181.050 ;
        RECT 502.950 180.600 505.050 181.050 ;
        RECT 544.950 180.600 547.050 181.050 ;
        RECT 157.950 179.400 547.050 180.600 ;
        RECT 157.950 178.950 160.050 179.400 ;
        RECT 502.950 178.950 505.050 179.400 ;
        RECT 544.950 178.950 547.050 179.400 ;
        RECT 268.950 177.600 271.050 178.050 ;
        RECT 475.950 177.600 478.050 178.050 ;
        RECT 481.950 177.600 484.050 178.050 ;
        RECT 559.950 177.600 562.050 178.050 ;
        RECT 268.950 176.400 562.050 177.600 ;
        RECT 268.950 175.950 271.050 176.400 ;
        RECT 475.950 175.950 478.050 176.400 ;
        RECT 481.950 175.950 484.050 176.400 ;
        RECT 559.950 175.950 562.050 176.400 ;
        RECT 79.950 174.600 82.050 175.050 ;
        RECT 112.950 174.600 115.050 175.050 ;
        RECT 118.950 174.600 121.050 175.050 ;
        RECT 79.950 173.400 121.050 174.600 ;
        RECT 79.950 172.950 82.050 173.400 ;
        RECT 112.950 172.950 115.050 173.400 ;
        RECT 118.950 172.950 121.050 173.400 ;
        RECT 121.950 174.600 124.050 175.050 ;
        RECT 199.950 174.600 202.050 175.050 ;
        RECT 121.950 173.400 202.050 174.600 ;
        RECT 121.950 172.950 124.050 173.400 ;
        RECT 199.950 172.950 202.050 173.400 ;
        RECT 364.950 174.600 367.050 175.050 ;
        RECT 382.950 174.600 385.050 175.050 ;
        RECT 364.950 173.400 385.050 174.600 ;
        RECT 364.950 172.950 367.050 173.400 ;
        RECT 382.950 172.950 385.050 173.400 ;
        RECT 412.950 174.600 415.050 175.050 ;
        RECT 460.950 174.600 463.050 175.050 ;
        RECT 412.950 173.400 463.050 174.600 ;
        RECT 412.950 172.950 415.050 173.400 ;
        RECT 460.950 172.950 463.050 173.400 ;
        RECT 613.950 174.600 616.050 175.050 ;
        RECT 649.950 174.600 652.050 175.050 ;
        RECT 685.950 174.600 688.050 175.050 ;
        RECT 613.950 173.400 688.050 174.600 ;
        RECT 613.950 172.950 616.050 173.400 ;
        RECT 649.950 172.950 652.050 173.400 ;
        RECT 685.950 172.950 688.050 173.400 ;
        RECT 70.950 171.600 73.050 172.050 ;
        RECT 79.950 171.600 82.050 172.050 ;
        RECT 70.950 170.400 82.050 171.600 ;
        RECT 70.950 169.950 73.050 170.400 ;
        RECT 79.950 169.950 82.050 170.400 ;
        RECT 85.950 171.600 88.050 172.050 ;
        RECT 163.950 171.600 166.050 172.050 ;
        RECT 193.950 171.600 196.050 172.050 ;
        RECT 85.950 170.400 196.050 171.600 ;
        RECT 85.950 169.950 88.050 170.400 ;
        RECT 163.950 169.950 166.050 170.400 ;
        RECT 193.950 169.950 196.050 170.400 ;
        RECT 205.950 171.600 208.050 172.050 ;
        RECT 238.950 171.600 241.050 172.050 ;
        RECT 259.950 171.600 262.050 172.050 ;
        RECT 205.950 170.400 262.050 171.600 ;
        RECT 205.950 169.950 208.050 170.400 ;
        RECT 238.950 169.950 241.050 170.400 ;
        RECT 259.950 169.950 262.050 170.400 ;
        RECT 283.950 171.600 286.050 172.050 ;
        RECT 322.950 171.600 325.050 172.050 ;
        RECT 283.950 170.400 325.050 171.600 ;
        RECT 283.950 169.950 286.050 170.400 ;
        RECT 322.950 169.950 325.050 170.400 ;
        RECT 379.950 171.600 382.050 172.050 ;
        RECT 445.950 171.600 448.050 172.050 ;
        RECT 379.950 170.400 448.050 171.600 ;
        RECT 379.950 169.950 382.050 170.400 ;
        RECT 445.950 169.950 448.050 170.400 ;
        RECT 607.950 171.600 610.050 172.050 ;
        RECT 643.950 171.600 646.050 172.050 ;
        RECT 607.950 170.400 646.050 171.600 ;
        RECT 607.950 169.950 610.050 170.400 ;
        RECT 643.950 169.950 646.050 170.400 ;
        RECT 289.950 168.600 292.050 169.050 ;
        RECT 301.950 168.600 304.050 169.050 ;
        RECT 325.950 168.600 328.050 169.050 ;
        RECT 289.950 167.400 328.050 168.600 ;
        RECT 289.950 166.950 292.050 167.400 ;
        RECT 301.950 166.950 304.050 167.400 ;
        RECT 325.950 166.950 328.050 167.400 ;
        RECT 328.950 168.600 331.050 169.050 ;
        RECT 349.950 168.600 352.050 169.050 ;
        RECT 376.950 168.600 379.050 169.050 ;
        RECT 406.950 168.600 409.050 169.050 ;
        RECT 328.950 167.400 372.600 168.600 ;
        RECT 328.950 166.950 331.050 167.400 ;
        RECT 349.950 166.950 352.050 167.400 ;
        RECT 371.400 166.050 372.600 167.400 ;
        RECT 376.950 167.400 409.050 168.600 ;
        RECT 376.950 166.950 379.050 167.400 ;
        RECT 406.950 166.950 409.050 167.400 ;
        RECT 451.950 168.600 454.050 169.050 ;
        RECT 469.950 168.600 472.050 169.050 ;
        RECT 523.950 168.600 526.050 169.050 ;
        RECT 451.950 167.400 472.050 168.600 ;
        RECT 451.950 166.950 454.050 167.400 ;
        RECT 469.950 166.950 472.050 167.400 ;
        RECT 473.400 167.400 526.050 168.600 ;
        RECT 67.950 165.600 70.050 166.050 ;
        RECT 76.950 165.600 79.050 166.050 ;
        RECT 67.950 164.400 79.050 165.600 ;
        RECT 67.950 163.950 70.050 164.400 ;
        RECT 76.950 163.950 79.050 164.400 ;
        RECT 166.950 165.600 169.050 166.050 ;
        RECT 187.950 165.600 190.050 166.050 ;
        RECT 166.950 164.400 190.050 165.600 ;
        RECT 166.950 163.950 169.050 164.400 ;
        RECT 187.950 163.950 190.050 164.400 ;
        RECT 370.950 165.600 373.050 166.050 ;
        RECT 379.950 165.600 382.050 166.050 ;
        RECT 370.950 164.400 382.050 165.600 ;
        RECT 370.950 163.950 373.050 164.400 ;
        RECT 379.950 163.950 382.050 164.400 ;
        RECT 448.950 165.600 451.050 166.050 ;
        RECT 473.400 165.600 474.600 167.400 ;
        RECT 523.950 166.950 526.050 167.400 ;
        RECT 562.950 168.600 565.050 169.050 ;
        RECT 562.950 167.400 606.600 168.600 ;
        RECT 562.950 166.950 565.050 167.400 ;
        RECT 605.400 166.050 606.600 167.400 ;
        RECT 448.950 164.400 474.600 165.600 ;
        RECT 526.950 165.600 529.050 166.050 ;
        RECT 529.950 165.600 532.050 166.050 ;
        RECT 559.950 165.600 562.050 166.050 ;
        RECT 526.950 164.400 562.050 165.600 ;
        RECT 448.950 163.950 451.050 164.400 ;
        RECT 526.950 163.950 529.050 164.400 ;
        RECT 529.950 163.950 532.050 164.400 ;
        RECT 559.950 163.950 562.050 164.400 ;
        RECT 604.950 163.950 607.050 166.050 ;
        RECT 610.950 165.600 613.050 166.050 ;
        RECT 652.950 165.600 655.050 166.050 ;
        RECT 679.950 165.600 682.050 166.050 ;
        RECT 610.950 164.400 651.600 165.600 ;
        RECT 610.950 163.950 613.050 164.400 ;
        RECT 118.950 162.600 121.050 163.050 ;
        RECT 139.950 162.600 142.050 163.050 ;
        RECT 118.950 161.400 142.050 162.600 ;
        RECT 118.950 160.950 121.050 161.400 ;
        RECT 139.950 160.950 142.050 161.400 ;
        RECT 442.950 162.600 445.050 163.050 ;
        RECT 478.950 162.600 481.050 163.050 ;
        RECT 442.950 161.400 481.050 162.600 ;
        RECT 442.950 160.950 445.050 161.400 ;
        RECT 478.950 160.950 481.050 161.400 ;
        RECT 520.950 162.600 523.050 163.050 ;
        RECT 637.950 162.600 640.050 163.050 ;
        RECT 646.950 162.600 649.050 163.050 ;
        RECT 520.950 161.400 649.050 162.600 ;
        RECT 650.400 162.600 651.600 164.400 ;
        RECT 652.950 164.400 682.050 165.600 ;
        RECT 652.950 163.950 655.050 164.400 ;
        RECT 679.950 163.950 682.050 164.400 ;
        RECT 691.950 162.600 694.050 163.050 ;
        RECT 650.400 161.400 694.050 162.600 ;
        RECT 520.950 160.950 523.050 161.400 ;
        RECT 637.950 160.950 640.050 161.400 ;
        RECT 646.950 160.950 649.050 161.400 ;
        RECT 691.950 160.950 694.050 161.400 ;
        RECT 586.950 159.600 589.050 160.050 ;
        RECT 610.950 159.600 613.050 160.050 ;
        RECT 586.950 158.400 613.050 159.600 ;
        RECT 586.950 157.950 589.050 158.400 ;
        RECT 610.950 157.950 613.050 158.400 ;
        RECT 124.950 132.600 127.050 133.050 ;
        RECT 202.950 132.600 205.050 133.050 ;
        RECT 124.950 131.400 205.050 132.600 ;
        RECT 124.950 130.950 127.050 131.400 ;
        RECT 202.950 130.950 205.050 131.400 ;
        RECT 370.950 132.600 373.050 133.050 ;
        RECT 376.950 132.600 379.050 133.050 ;
        RECT 370.950 131.400 379.050 132.600 ;
        RECT 370.950 130.950 373.050 131.400 ;
        RECT 376.950 130.950 379.050 131.400 ;
        RECT 424.950 132.600 427.050 133.050 ;
        RECT 538.950 132.600 541.050 133.050 ;
        RECT 553.950 132.600 556.050 133.050 ;
        RECT 565.950 132.600 568.050 133.050 ;
        RECT 424.950 131.400 568.050 132.600 ;
        RECT 424.950 130.950 427.050 131.400 ;
        RECT 538.950 130.950 541.050 131.400 ;
        RECT 553.950 130.950 556.050 131.400 ;
        RECT 565.950 130.950 568.050 131.400 ;
        RECT 649.950 132.600 652.050 133.050 ;
        RECT 694.950 132.600 697.050 133.050 ;
        RECT 649.950 131.400 697.050 132.600 ;
        RECT 649.950 130.950 652.050 131.400 ;
        RECT 694.950 130.950 697.050 131.400 ;
        RECT 196.950 129.600 199.050 130.050 ;
        RECT 223.950 129.600 226.050 130.050 ;
        RECT 196.950 128.400 226.050 129.600 ;
        RECT 196.950 127.950 199.050 128.400 ;
        RECT 223.950 127.950 226.050 128.400 ;
        RECT 253.950 129.600 256.050 130.050 ;
        RECT 268.950 129.600 271.050 130.050 ;
        RECT 286.950 129.600 289.050 130.050 ;
        RECT 253.950 128.400 289.050 129.600 ;
        RECT 253.950 127.950 256.050 128.400 ;
        RECT 268.950 127.950 271.050 128.400 ;
        RECT 286.950 127.950 289.050 128.400 ;
        RECT 457.950 129.600 460.050 130.050 ;
        RECT 490.950 129.600 493.050 130.050 ;
        RECT 457.950 128.400 493.050 129.600 ;
        RECT 457.950 127.950 460.050 128.400 ;
        RECT 490.950 127.950 493.050 128.400 ;
        RECT 655.950 129.600 658.050 130.050 ;
        RECT 664.950 129.600 667.050 130.050 ;
        RECT 655.950 128.400 667.050 129.600 ;
        RECT 655.950 127.950 658.050 128.400 ;
        RECT 664.950 127.950 667.050 128.400 ;
        RECT 688.950 129.600 691.050 130.050 ;
        RECT 688.950 128.400 696.600 129.600 ;
        RECT 688.950 127.950 691.050 128.400 ;
        RECT 70.950 126.600 73.050 127.050 ;
        RECT 103.950 126.600 106.050 127.050 ;
        RECT 70.950 125.400 106.050 126.600 ;
        RECT 70.950 124.950 73.050 125.400 ;
        RECT 103.950 124.950 106.050 125.400 ;
        RECT 142.950 124.950 145.050 127.050 ;
        RECT 148.950 126.600 151.050 127.050 ;
        RECT 184.950 126.600 187.050 127.050 ;
        RECT 148.950 125.400 187.050 126.600 ;
        RECT 148.950 124.950 151.050 125.400 ;
        RECT 184.950 124.950 187.050 125.400 ;
        RECT 217.950 126.600 220.050 127.050 ;
        RECT 229.950 126.600 232.050 127.050 ;
        RECT 217.950 125.400 232.050 126.600 ;
        RECT 217.950 124.950 220.050 125.400 ;
        RECT 229.950 124.950 232.050 125.400 ;
        RECT 361.950 126.600 364.050 127.050 ;
        RECT 373.950 126.600 376.050 127.050 ;
        RECT 361.950 125.400 376.050 126.600 ;
        RECT 361.950 124.950 364.050 125.400 ;
        RECT 373.950 124.950 376.050 125.400 ;
        RECT 415.950 124.950 418.050 127.050 ;
        RECT 421.950 126.600 424.050 127.050 ;
        RECT 454.950 126.600 457.050 127.050 ;
        RECT 421.950 125.400 457.050 126.600 ;
        RECT 421.950 124.950 424.050 125.400 ;
        RECT 454.950 124.950 457.050 125.400 ;
        RECT 568.950 126.600 571.050 127.050 ;
        RECT 574.950 126.600 577.050 127.050 ;
        RECT 568.950 125.400 577.050 126.600 ;
        RECT 568.950 124.950 571.050 125.400 ;
        RECT 574.950 124.950 577.050 125.400 ;
        RECT 580.950 126.600 583.050 127.050 ;
        RECT 652.950 126.600 655.050 127.050 ;
        RECT 580.950 125.400 655.050 126.600 ;
        RECT 580.950 124.950 583.050 125.400 ;
        RECT 652.950 124.950 655.050 125.400 ;
        RECT 679.950 126.600 682.050 127.050 ;
        RECT 691.950 126.600 694.050 127.050 ;
        RECT 679.950 125.400 694.050 126.600 ;
        RECT 695.400 126.600 696.600 128.400 ;
        RECT 730.950 126.600 733.050 127.050 ;
        RECT 695.400 125.400 733.050 126.600 ;
        RECT 679.950 124.950 682.050 125.400 ;
        RECT 691.950 124.950 694.050 125.400 ;
        RECT 730.950 124.950 733.050 125.400 ;
        RECT 37.950 123.600 40.050 124.050 ;
        RECT 100.950 123.600 103.050 124.050 ;
        RECT 37.950 122.400 103.050 123.600 ;
        RECT 37.950 121.950 40.050 122.400 ;
        RECT 100.950 121.950 103.050 122.400 ;
        RECT 106.950 123.600 109.050 124.050 ;
        RECT 124.950 123.600 127.050 124.050 ;
        RECT 106.950 122.400 127.050 123.600 ;
        RECT 106.950 121.950 109.050 122.400 ;
        RECT 124.950 121.950 127.050 122.400 ;
        RECT 143.400 121.050 144.600 124.950 ;
        RECT 145.950 123.600 148.050 124.050 ;
        RECT 160.950 123.600 163.050 124.050 ;
        RECT 145.950 122.400 163.050 123.600 ;
        RECT 145.950 121.950 148.050 122.400 ;
        RECT 160.950 121.950 163.050 122.400 ;
        RECT 226.950 123.600 229.050 124.050 ;
        RECT 235.950 123.600 238.050 124.050 ;
        RECT 226.950 122.400 238.050 123.600 ;
        RECT 226.950 121.950 229.050 122.400 ;
        RECT 235.950 121.950 238.050 122.400 ;
        RECT 244.950 123.600 247.050 124.050 ;
        RECT 262.950 123.600 265.050 124.050 ;
        RECT 244.950 122.400 265.050 123.600 ;
        RECT 244.950 121.950 247.050 122.400 ;
        RECT 262.950 121.950 265.050 122.400 ;
        RECT 301.950 123.600 304.050 124.050 ;
        RECT 334.950 123.600 337.050 124.050 ;
        RECT 403.950 123.600 406.050 124.050 ;
        RECT 301.950 122.400 406.050 123.600 ;
        RECT 416.400 123.600 417.600 124.950 ;
        RECT 466.950 123.600 469.050 124.050 ;
        RECT 416.400 122.400 469.050 123.600 ;
        RECT 301.950 121.950 304.050 122.400 ;
        RECT 334.950 121.950 337.050 122.400 ;
        RECT 403.950 121.950 406.050 122.400 ;
        RECT 466.950 121.950 469.050 122.400 ;
        RECT 514.950 123.600 517.050 124.050 ;
        RECT 541.950 123.600 544.050 124.050 ;
        RECT 550.950 123.600 553.050 124.050 ;
        RECT 514.950 122.400 553.050 123.600 ;
        RECT 514.950 121.950 517.050 122.400 ;
        RECT 541.950 121.950 544.050 122.400 ;
        RECT 550.950 121.950 553.050 122.400 ;
        RECT 565.950 123.600 568.050 124.050 ;
        RECT 613.950 123.600 616.050 124.050 ;
        RECT 622.950 123.600 625.050 124.050 ;
        RECT 655.950 123.600 658.050 124.050 ;
        RECT 565.950 122.400 579.600 123.600 ;
        RECT 565.950 121.950 568.050 122.400 ;
        RECT 578.400 121.050 579.600 122.400 ;
        RECT 613.950 122.400 658.050 123.600 ;
        RECT 613.950 121.950 616.050 122.400 ;
        RECT 622.950 121.950 625.050 122.400 ;
        RECT 655.950 121.950 658.050 122.400 ;
        RECT 67.950 120.600 70.050 121.050 ;
        RECT 73.950 120.600 76.050 121.050 ;
        RECT 67.950 119.400 76.050 120.600 ;
        RECT 67.950 118.950 70.050 119.400 ;
        RECT 73.950 118.950 76.050 119.400 ;
        RECT 142.950 118.950 145.050 121.050 ;
        RECT 187.950 120.600 190.050 121.050 ;
        RECT 196.950 120.600 199.050 121.050 ;
        RECT 187.950 119.400 199.050 120.600 ;
        RECT 187.950 118.950 190.050 119.400 ;
        RECT 196.950 118.950 199.050 119.400 ;
        RECT 202.950 120.600 205.050 121.050 ;
        RECT 220.950 120.600 223.050 121.050 ;
        RECT 202.950 119.400 223.050 120.600 ;
        RECT 202.950 118.950 205.050 119.400 ;
        RECT 220.950 118.950 223.050 119.400 ;
        RECT 229.950 120.600 232.050 121.050 ;
        RECT 265.950 120.600 268.050 121.050 ;
        RECT 229.950 119.400 268.050 120.600 ;
        RECT 229.950 118.950 232.050 119.400 ;
        RECT 265.950 118.950 268.050 119.400 ;
        RECT 325.950 120.600 328.050 121.050 ;
        RECT 340.950 120.600 343.050 121.050 ;
        RECT 325.950 119.400 343.050 120.600 ;
        RECT 325.950 118.950 328.050 119.400 ;
        RECT 340.950 118.950 343.050 119.400 ;
        RECT 418.950 120.600 421.050 121.050 ;
        RECT 424.950 120.600 427.050 121.050 ;
        RECT 418.950 119.400 427.050 120.600 ;
        RECT 418.950 118.950 421.050 119.400 ;
        RECT 424.950 118.950 427.050 119.400 ;
        RECT 535.950 120.600 538.050 121.050 ;
        RECT 568.950 120.600 571.050 121.050 ;
        RECT 535.950 119.400 571.050 120.600 ;
        RECT 535.950 118.950 538.050 119.400 ;
        RECT 568.950 118.950 571.050 119.400 ;
        RECT 577.950 118.950 580.050 121.050 ;
        RECT 34.950 117.600 37.050 118.050 ;
        RECT 118.950 117.600 121.050 118.050 ;
        RECT 34.950 116.400 121.050 117.600 ;
        RECT 34.950 115.950 37.050 116.400 ;
        RECT 118.950 115.950 121.050 116.400 ;
        RECT 382.950 117.600 385.050 118.050 ;
        RECT 430.950 117.600 433.050 118.050 ;
        RECT 382.950 116.400 433.050 117.600 ;
        RECT 382.950 115.950 385.050 116.400 ;
        RECT 430.950 115.950 433.050 116.400 ;
        RECT 448.950 117.600 451.050 118.050 ;
        RECT 541.950 117.600 544.050 118.050 ;
        RECT 448.950 116.400 544.050 117.600 ;
        RECT 448.950 115.950 451.050 116.400 ;
        RECT 541.950 115.950 544.050 116.400 ;
        RECT 607.950 117.600 610.050 118.050 ;
        RECT 619.950 117.600 622.050 118.050 ;
        RECT 607.950 116.400 622.050 117.600 ;
        RECT 607.950 115.950 610.050 116.400 ;
        RECT 619.950 115.950 622.050 116.400 ;
        RECT 283.950 114.600 286.050 115.050 ;
        RECT 424.950 114.600 427.050 115.050 ;
        RECT 283.950 113.400 427.050 114.600 ;
        RECT 283.950 112.950 286.050 113.400 ;
        RECT 424.950 112.950 427.050 113.400 ;
        RECT 361.950 111.600 364.050 112.050 ;
        RECT 463.950 111.600 466.050 112.050 ;
        RECT 361.950 110.400 466.050 111.600 ;
        RECT 361.950 109.950 364.050 110.400 ;
        RECT 463.950 109.950 466.050 110.400 ;
        RECT 481.950 108.600 484.050 109.050 ;
        RECT 490.950 108.600 493.050 109.050 ;
        RECT 568.950 108.600 571.050 109.050 ;
        RECT 481.950 107.400 571.050 108.600 ;
        RECT 481.950 106.950 484.050 107.400 ;
        RECT 490.950 106.950 493.050 107.400 ;
        RECT 568.950 106.950 571.050 107.400 ;
        RECT 223.950 102.600 226.050 103.050 ;
        RECT 298.950 102.600 301.050 103.050 ;
        RECT 334.950 102.600 337.050 103.050 ;
        RECT 223.950 101.400 337.050 102.600 ;
        RECT 223.950 100.950 226.050 101.400 ;
        RECT 298.950 100.950 301.050 101.400 ;
        RECT 334.950 100.950 337.050 101.400 ;
        RECT 337.950 102.600 340.050 103.050 ;
        RECT 421.950 102.600 424.050 103.050 ;
        RECT 337.950 101.400 424.050 102.600 ;
        RECT 337.950 100.950 340.050 101.400 ;
        RECT 421.950 100.950 424.050 101.400 ;
        RECT 616.950 102.600 619.050 103.050 ;
        RECT 652.950 102.600 655.050 103.050 ;
        RECT 703.950 102.600 706.050 103.050 ;
        RECT 709.950 102.600 712.050 103.050 ;
        RECT 739.950 102.600 742.050 103.050 ;
        RECT 616.950 101.400 742.050 102.600 ;
        RECT 616.950 100.950 619.050 101.400 ;
        RECT 652.950 100.950 655.050 101.400 ;
        RECT 703.950 100.950 706.050 101.400 ;
        RECT 709.950 100.950 712.050 101.400 ;
        RECT 739.950 100.950 742.050 101.400 ;
        RECT 28.950 99.600 31.050 100.050 ;
        RECT 106.950 99.600 109.050 100.050 ;
        RECT 28.950 98.400 109.050 99.600 ;
        RECT 28.950 97.950 31.050 98.400 ;
        RECT 71.400 94.050 72.600 98.400 ;
        RECT 106.950 97.950 109.050 98.400 ;
        RECT 217.950 99.600 220.050 100.050 ;
        RECT 268.950 99.600 271.050 100.050 ;
        RECT 295.950 99.600 298.050 100.050 ;
        RECT 301.950 99.600 304.050 100.050 ;
        RECT 340.950 99.600 343.050 100.050 ;
        RECT 217.950 98.400 267.600 99.600 ;
        RECT 217.950 97.950 220.050 98.400 ;
        RECT 73.950 96.600 76.050 97.050 ;
        RECT 139.950 96.600 142.050 97.050 ;
        RECT 73.950 95.400 142.050 96.600 ;
        RECT 73.950 94.950 76.050 95.400 ;
        RECT 139.950 94.950 142.050 95.400 ;
        RECT 148.950 96.600 151.050 97.050 ;
        RECT 244.950 96.600 247.050 97.050 ;
        RECT 148.950 95.400 247.050 96.600 ;
        RECT 148.950 94.950 151.050 95.400 ;
        RECT 244.950 94.950 247.050 95.400 ;
        RECT 266.400 94.050 267.600 98.400 ;
        RECT 268.950 98.400 343.050 99.600 ;
        RECT 268.950 97.950 271.050 98.400 ;
        RECT 295.950 97.950 298.050 98.400 ;
        RECT 301.950 97.950 304.050 98.400 ;
        RECT 340.950 97.950 343.050 98.400 ;
        RECT 346.950 99.600 349.050 100.050 ;
        RECT 382.950 99.600 385.050 100.050 ;
        RECT 346.950 98.400 385.050 99.600 ;
        RECT 346.950 97.950 349.050 98.400 ;
        RECT 382.950 97.950 385.050 98.400 ;
        RECT 412.950 99.600 415.050 100.050 ;
        RECT 496.950 99.600 499.050 100.050 ;
        RECT 412.950 98.400 499.050 99.600 ;
        RECT 412.950 97.950 415.050 98.400 ;
        RECT 496.950 97.950 499.050 98.400 ;
        RECT 616.950 99.600 619.050 100.050 ;
        RECT 658.950 99.600 661.050 100.050 ;
        RECT 616.950 98.400 661.050 99.600 ;
        RECT 616.950 97.950 619.050 98.400 ;
        RECT 658.950 97.950 661.050 98.400 ;
        RECT 700.950 99.600 703.050 100.050 ;
        RECT 706.950 99.600 709.050 100.050 ;
        RECT 700.950 98.400 709.050 99.600 ;
        RECT 700.950 97.950 703.050 98.400 ;
        RECT 706.950 97.950 709.050 98.400 ;
        RECT 268.950 94.950 271.050 97.050 ;
        RECT 271.950 96.600 274.050 97.050 ;
        RECT 388.950 96.600 391.050 97.050 ;
        RECT 271.950 95.400 391.050 96.600 ;
        RECT 271.950 94.950 274.050 95.400 ;
        RECT 388.950 94.950 391.050 95.400 ;
        RECT 418.950 96.600 421.050 97.050 ;
        RECT 427.950 96.600 430.050 97.050 ;
        RECT 418.950 95.400 430.050 96.600 ;
        RECT 418.950 94.950 421.050 95.400 ;
        RECT 427.950 94.950 430.050 95.400 ;
        RECT 472.950 96.600 475.050 97.050 ;
        RECT 478.950 96.600 481.050 97.050 ;
        RECT 472.950 95.400 481.050 96.600 ;
        RECT 472.950 94.950 475.050 95.400 ;
        RECT 478.950 94.950 481.050 95.400 ;
        RECT 562.950 96.600 565.050 97.050 ;
        RECT 571.950 96.600 574.050 97.050 ;
        RECT 562.950 95.400 574.050 96.600 ;
        RECT 562.950 94.950 565.050 95.400 ;
        RECT 571.950 94.950 574.050 95.400 ;
        RECT 604.950 96.600 607.050 97.050 ;
        RECT 619.950 96.600 622.050 97.050 ;
        RECT 604.950 95.400 622.050 96.600 ;
        RECT 604.950 94.950 607.050 95.400 ;
        RECT 619.950 94.950 622.050 95.400 ;
        RECT 721.950 96.600 724.050 97.050 ;
        RECT 736.950 96.600 739.050 97.050 ;
        RECT 721.950 95.400 739.050 96.600 ;
        RECT 721.950 94.950 724.050 95.400 ;
        RECT 736.950 94.950 739.050 95.400 ;
        RECT 70.950 91.950 73.050 94.050 ;
        RECT 184.950 93.600 187.050 94.050 ;
        RECT 214.950 93.600 217.050 94.050 ;
        RECT 184.950 92.400 217.050 93.600 ;
        RECT 184.950 91.950 187.050 92.400 ;
        RECT 214.950 91.950 217.050 92.400 ;
        RECT 220.950 93.600 223.050 94.050 ;
        RECT 259.950 93.600 262.050 94.050 ;
        RECT 220.950 92.400 262.050 93.600 ;
        RECT 220.950 91.950 223.050 92.400 ;
        RECT 259.950 91.950 262.050 92.400 ;
        RECT 265.950 91.950 268.050 94.050 ;
        RECT 64.950 90.600 67.050 91.050 ;
        RECT 70.950 90.600 73.050 91.050 ;
        RECT 64.950 89.400 73.050 90.600 ;
        RECT 64.950 88.950 67.050 89.400 ;
        RECT 70.950 88.950 73.050 89.400 ;
        RECT 145.950 90.600 148.050 91.050 ;
        RECT 178.950 90.600 181.050 91.050 ;
        RECT 145.950 89.400 181.050 90.600 ;
        RECT 145.950 88.950 148.050 89.400 ;
        RECT 178.950 88.950 181.050 89.400 ;
        RECT 265.950 90.600 268.050 91.050 ;
        RECT 269.400 90.600 270.600 94.950 ;
        RECT 343.950 93.600 346.050 94.050 ;
        RECT 349.950 93.600 352.050 94.050 ;
        RECT 343.950 92.400 352.050 93.600 ;
        RECT 343.950 91.950 346.050 92.400 ;
        RECT 349.950 91.950 352.050 92.400 ;
        RECT 385.950 93.600 388.050 94.050 ;
        RECT 391.950 93.600 394.050 94.050 ;
        RECT 385.950 92.400 394.050 93.600 ;
        RECT 385.950 91.950 388.050 92.400 ;
        RECT 391.950 91.950 394.050 92.400 ;
        RECT 664.950 93.600 667.050 94.050 ;
        RECT 697.950 93.600 700.050 94.050 ;
        RECT 664.950 92.400 700.050 93.600 ;
        RECT 664.950 91.950 667.050 92.400 ;
        RECT 697.950 91.950 700.050 92.400 ;
        RECT 265.950 89.400 270.600 90.600 ;
        RECT 307.950 90.600 310.050 91.050 ;
        RECT 379.950 90.600 382.050 91.050 ;
        RECT 307.950 89.400 382.050 90.600 ;
        RECT 265.950 88.950 268.050 89.400 ;
        RECT 307.950 88.950 310.050 89.400 ;
        RECT 379.950 88.950 382.050 89.400 ;
        RECT 505.950 90.600 508.050 91.050 ;
        RECT 544.950 90.600 547.050 91.050 ;
        RECT 547.950 90.600 550.050 91.050 ;
        RECT 505.950 89.400 550.050 90.600 ;
        RECT 505.950 88.950 508.050 89.400 ;
        RECT 544.950 88.950 547.050 89.400 ;
        RECT 547.950 88.950 550.050 89.400 ;
        RECT 595.950 90.600 598.050 91.050 ;
        RECT 661.950 90.600 664.050 91.050 ;
        RECT 595.950 89.400 664.050 90.600 ;
        RECT 595.950 88.950 598.050 89.400 ;
        RECT 661.950 88.950 664.050 89.400 ;
        RECT 379.950 87.600 382.050 88.050 ;
        RECT 460.950 87.600 463.050 88.050 ;
        RECT 469.950 87.600 472.050 88.050 ;
        RECT 379.950 86.400 472.050 87.600 ;
        RECT 379.950 85.950 382.050 86.400 ;
        RECT 460.950 85.950 463.050 86.400 ;
        RECT 469.950 85.950 472.050 86.400 ;
        RECT 550.950 87.600 553.050 88.050 ;
        RECT 580.950 87.600 583.050 88.050 ;
        RECT 724.950 87.600 727.050 88.050 ;
        RECT 550.950 86.400 727.050 87.600 ;
        RECT 550.950 85.950 553.050 86.400 ;
        RECT 580.950 85.950 583.050 86.400 ;
        RECT 724.950 85.950 727.050 86.400 ;
        RECT 151.950 75.600 154.050 76.050 ;
        RECT 157.950 75.600 160.050 76.050 ;
        RECT 229.950 75.600 232.050 76.050 ;
        RECT 151.950 74.400 232.050 75.600 ;
        RECT 151.950 73.950 154.050 74.400 ;
        RECT 157.950 73.950 160.050 74.400 ;
        RECT 229.950 73.950 232.050 74.400 ;
        RECT 145.950 58.950 148.050 61.050 ;
        RECT 103.950 57.600 106.050 58.050 ;
        RECT 146.400 57.600 147.600 58.950 ;
        RECT 151.950 57.600 154.050 58.050 ;
        RECT 103.950 56.400 154.050 57.600 ;
        RECT 103.950 55.950 106.050 56.400 ;
        RECT 151.950 55.950 154.050 56.400 ;
        RECT 199.950 57.600 202.050 58.050 ;
        RECT 232.950 57.600 235.050 58.050 ;
        RECT 289.950 57.600 292.050 58.050 ;
        RECT 298.950 57.600 301.050 58.050 ;
        RECT 199.950 56.400 292.050 57.600 ;
        RECT 199.950 55.950 202.050 56.400 ;
        RECT 232.950 55.950 235.050 56.400 ;
        RECT 289.950 55.950 292.050 56.400 ;
        RECT 293.400 56.400 301.050 57.600 ;
        RECT 151.950 54.600 154.050 55.050 ;
        RECT 187.950 54.600 190.050 55.050 ;
        RECT 151.950 53.400 190.050 54.600 ;
        RECT 151.950 52.950 154.050 53.400 ;
        RECT 187.950 52.950 190.050 53.400 ;
        RECT 193.950 54.600 196.050 55.050 ;
        RECT 229.950 54.600 232.050 55.050 ;
        RECT 293.400 54.600 294.600 56.400 ;
        RECT 298.950 55.950 301.050 56.400 ;
        RECT 466.950 57.600 469.050 58.050 ;
        RECT 502.950 57.600 505.050 58.050 ;
        RECT 466.950 56.400 505.050 57.600 ;
        RECT 466.950 55.950 469.050 56.400 ;
        RECT 502.950 55.950 505.050 56.400 ;
        RECT 508.950 55.950 511.050 58.050 ;
        RECT 547.950 57.600 550.050 58.050 ;
        RECT 658.950 57.600 661.050 58.050 ;
        RECT 547.950 56.400 661.050 57.600 ;
        RECT 547.950 55.950 550.050 56.400 ;
        RECT 658.950 55.950 661.050 56.400 ;
        RECT 193.950 53.400 294.600 54.600 ;
        RECT 295.950 54.600 298.050 55.050 ;
        RECT 301.950 54.600 304.050 55.050 ;
        RECT 295.950 53.400 304.050 54.600 ;
        RECT 193.950 52.950 196.050 53.400 ;
        RECT 229.950 52.950 232.050 53.400 ;
        RECT 295.950 52.950 298.050 53.400 ;
        RECT 301.950 52.950 304.050 53.400 ;
        RECT 325.950 54.600 328.050 55.050 ;
        RECT 337.950 54.600 340.050 55.050 ;
        RECT 379.950 54.600 382.050 55.050 ;
        RECT 391.950 54.600 394.050 55.050 ;
        RECT 325.950 53.400 382.050 54.600 ;
        RECT 325.950 52.950 328.050 53.400 ;
        RECT 337.950 52.950 340.050 53.400 ;
        RECT 379.950 52.950 382.050 53.400 ;
        RECT 383.400 53.400 394.050 54.600 ;
        RECT 383.400 52.050 384.600 53.400 ;
        RECT 391.950 52.950 394.050 53.400 ;
        RECT 424.950 54.600 427.050 55.050 ;
        RECT 509.400 54.600 510.600 55.950 ;
        RECT 541.950 54.600 544.050 55.050 ;
        RECT 424.950 53.400 544.050 54.600 ;
        RECT 424.950 52.950 427.050 53.400 ;
        RECT 541.950 52.950 544.050 53.400 ;
        RECT 589.950 54.600 592.050 55.050 ;
        RECT 622.950 54.600 625.050 55.050 ;
        RECT 664.950 54.600 667.050 55.050 ;
        RECT 589.950 53.400 621.600 54.600 ;
        RECT 589.950 52.950 592.050 53.400 ;
        RECT 154.950 51.600 157.050 52.050 ;
        RECT 157.950 51.600 160.050 52.050 ;
        RECT 184.950 51.600 187.050 52.050 ;
        RECT 154.950 50.400 187.050 51.600 ;
        RECT 154.950 49.950 157.050 50.400 ;
        RECT 157.950 49.950 160.050 50.400 ;
        RECT 184.950 49.950 187.050 50.400 ;
        RECT 190.950 51.600 193.050 52.050 ;
        RECT 196.950 51.600 199.050 52.050 ;
        RECT 190.950 50.400 199.050 51.600 ;
        RECT 190.950 49.950 193.050 50.400 ;
        RECT 196.950 49.950 199.050 50.400 ;
        RECT 343.950 51.600 346.050 52.050 ;
        RECT 361.950 51.600 364.050 52.050 ;
        RECT 343.950 50.400 364.050 51.600 ;
        RECT 343.950 49.950 346.050 50.400 ;
        RECT 361.950 49.950 364.050 50.400 ;
        RECT 382.950 49.950 385.050 52.050 ;
        RECT 385.950 51.600 388.050 52.050 ;
        RECT 418.950 51.600 421.050 52.050 ;
        RECT 385.950 50.400 421.050 51.600 ;
        RECT 385.950 49.950 388.050 50.400 ;
        RECT 418.950 49.950 421.050 50.400 ;
        RECT 499.950 51.600 502.050 52.050 ;
        RECT 505.950 51.600 508.050 52.050 ;
        RECT 538.950 51.600 541.050 52.050 ;
        RECT 550.950 51.600 553.050 52.050 ;
        RECT 583.950 51.600 586.050 52.050 ;
        RECT 610.950 51.600 613.050 52.050 ;
        RECT 499.950 50.400 613.050 51.600 ;
        RECT 620.400 51.600 621.600 53.400 ;
        RECT 622.950 53.400 667.050 54.600 ;
        RECT 622.950 52.950 625.050 53.400 ;
        RECT 664.950 52.950 667.050 53.400 ;
        RECT 694.950 54.600 697.050 55.050 ;
        RECT 703.950 54.600 706.050 55.050 ;
        RECT 694.950 53.400 706.050 54.600 ;
        RECT 694.950 52.950 697.050 53.400 ;
        RECT 703.950 52.950 706.050 53.400 ;
        RECT 655.950 51.600 658.050 52.050 ;
        RECT 620.400 50.400 658.050 51.600 ;
        RECT 499.950 49.950 502.050 50.400 ;
        RECT 505.950 49.950 508.050 50.400 ;
        RECT 538.950 49.950 541.050 50.400 ;
        RECT 550.950 49.950 553.050 50.400 ;
        RECT 583.950 49.950 586.050 50.400 ;
        RECT 610.950 49.950 613.050 50.400 ;
        RECT 655.950 49.950 658.050 50.400 ;
        RECT 661.950 51.600 664.050 52.050 ;
        RECT 697.950 51.600 700.050 52.050 ;
        RECT 661.950 50.400 700.050 51.600 ;
        RECT 661.950 49.950 664.050 50.400 ;
        RECT 697.950 49.950 700.050 50.400 ;
        RECT 34.950 48.600 37.050 49.050 ;
        RECT 67.950 48.600 70.050 49.050 ;
        RECT 100.950 48.600 103.050 49.050 ;
        RECT 34.950 47.400 103.050 48.600 ;
        RECT 34.950 46.950 37.050 47.400 ;
        RECT 67.950 46.950 70.050 47.400 ;
        RECT 100.950 46.950 103.050 47.400 ;
        RECT 196.950 48.600 199.050 49.050 ;
        RECT 307.950 48.600 310.050 49.050 ;
        RECT 196.950 47.400 310.050 48.600 ;
        RECT 196.950 46.950 199.050 47.400 ;
        RECT 307.950 46.950 310.050 47.400 ;
        RECT 430.950 48.600 433.050 49.050 ;
        RECT 457.950 48.600 460.050 49.050 ;
        RECT 478.950 48.600 481.050 49.050 ;
        RECT 430.950 47.400 481.050 48.600 ;
        RECT 430.950 46.950 433.050 47.400 ;
        RECT 457.950 46.950 460.050 47.400 ;
        RECT 478.950 46.950 481.050 47.400 ;
        RECT 481.950 48.600 484.050 49.050 ;
        RECT 580.950 48.600 583.050 49.050 ;
        RECT 604.950 48.600 607.050 49.050 ;
        RECT 622.950 48.600 625.050 49.050 ;
        RECT 481.950 47.400 625.050 48.600 ;
        RECT 481.950 46.950 484.050 47.400 ;
        RECT 580.950 46.950 583.050 47.400 ;
        RECT 604.950 46.950 607.050 47.400 ;
        RECT 622.950 46.950 625.050 47.400 ;
        RECT 739.950 48.600 742.050 49.050 ;
        RECT 745.950 48.600 748.050 49.050 ;
        RECT 739.950 47.400 748.050 48.600 ;
        RECT 739.950 46.950 742.050 47.400 ;
        RECT 745.950 46.950 748.050 47.400 ;
        RECT 40.950 45.600 43.050 46.050 ;
        RECT 112.950 45.600 115.050 46.050 ;
        RECT 136.950 45.600 139.050 46.050 ;
        RECT 40.950 44.400 139.050 45.600 ;
        RECT 40.950 43.950 43.050 44.400 ;
        RECT 112.950 43.950 115.050 44.400 ;
        RECT 136.950 43.950 139.050 44.400 ;
        RECT 184.950 45.600 187.050 46.050 ;
        RECT 262.950 45.600 265.050 46.050 ;
        RECT 184.950 44.400 265.050 45.600 ;
        RECT 184.950 43.950 187.050 44.400 ;
        RECT 262.950 43.950 265.050 44.400 ;
        RECT 289.950 45.600 292.050 46.050 ;
        RECT 376.950 45.600 379.050 46.050 ;
        RECT 289.950 44.400 379.050 45.600 ;
        RECT 289.950 43.950 292.050 44.400 ;
        RECT 376.950 43.950 379.050 44.400 ;
        RECT 115.950 42.600 118.050 43.050 ;
        RECT 148.950 42.600 151.050 43.050 ;
        RECT 115.950 41.400 151.050 42.600 ;
        RECT 115.950 40.950 118.050 41.400 ;
        RECT 148.950 40.950 151.050 41.400 ;
        RECT 220.950 33.600 223.050 34.050 ;
        RECT 271.950 33.600 274.050 34.050 ;
        RECT 220.950 32.400 274.050 33.600 ;
        RECT 220.950 31.950 223.050 32.400 ;
        RECT 271.950 31.950 274.050 32.400 ;
        RECT 424.950 33.600 427.050 34.050 ;
        RECT 460.950 33.600 463.050 34.050 ;
        RECT 544.950 33.600 547.050 34.050 ;
        RECT 424.950 32.400 547.050 33.600 ;
        RECT 424.950 31.950 427.050 32.400 ;
        RECT 460.950 31.950 463.050 32.400 ;
        RECT 544.950 31.950 547.050 32.400 ;
        RECT 79.950 30.600 82.050 31.050 ;
        RECT 145.950 30.600 148.050 31.050 ;
        RECT 184.950 30.600 187.050 31.050 ;
        RECT 79.950 29.400 187.050 30.600 ;
        RECT 79.950 28.950 82.050 29.400 ;
        RECT 145.950 28.950 148.050 29.400 ;
        RECT 184.950 28.950 187.050 29.400 ;
        RECT 268.950 30.600 271.050 31.050 ;
        RECT 334.950 30.600 337.050 31.050 ;
        RECT 379.950 30.600 382.050 31.050 ;
        RECT 508.950 30.600 511.050 31.050 ;
        RECT 268.950 29.400 511.050 30.600 ;
        RECT 268.950 28.950 271.050 29.400 ;
        RECT 334.950 28.950 337.050 29.400 ;
        RECT 379.950 28.950 382.050 29.400 ;
        RECT 508.950 28.950 511.050 29.400 ;
        RECT 118.950 27.600 121.050 28.050 ;
        RECT 148.950 27.600 151.050 28.050 ;
        RECT 118.950 26.400 151.050 27.600 ;
        RECT 118.950 25.950 121.050 26.400 ;
        RECT 148.950 25.950 151.050 26.400 ;
        RECT 184.950 27.600 187.050 28.050 ;
        RECT 199.950 27.600 202.050 28.050 ;
        RECT 184.950 26.400 202.050 27.600 ;
        RECT 184.950 25.950 187.050 26.400 ;
        RECT 199.950 25.950 202.050 26.400 ;
        RECT 214.950 27.600 217.050 28.050 ;
        RECT 253.950 27.600 256.050 28.050 ;
        RECT 214.950 26.400 256.050 27.600 ;
        RECT 214.950 25.950 217.050 26.400 ;
        RECT 253.950 25.950 256.050 26.400 ;
        RECT 307.950 27.600 310.050 28.050 ;
        RECT 313.950 27.600 316.050 28.050 ;
        RECT 307.950 26.400 316.050 27.600 ;
        RECT 307.950 25.950 310.050 26.400 ;
        RECT 313.950 25.950 316.050 26.400 ;
        RECT 316.950 27.600 319.050 28.050 ;
        RECT 343.950 27.600 346.050 28.050 ;
        RECT 316.950 26.400 346.050 27.600 ;
        RECT 316.950 25.950 319.050 26.400 ;
        RECT 343.950 25.950 346.050 26.400 ;
        RECT 346.950 27.600 349.050 28.050 ;
        RECT 427.950 27.600 430.050 28.050 ;
        RECT 346.950 26.400 430.050 27.600 ;
        RECT 346.950 25.950 349.050 26.400 ;
        RECT 427.950 25.950 430.050 26.400 ;
        RECT 505.950 27.600 508.050 28.050 ;
        RECT 535.950 27.600 538.050 28.050 ;
        RECT 505.950 26.400 538.050 27.600 ;
        RECT 505.950 25.950 508.050 26.400 ;
        RECT 535.950 25.950 538.050 26.400 ;
        RECT 544.950 27.600 547.050 28.050 ;
        RECT 607.950 27.600 610.050 28.050 ;
        RECT 625.950 27.600 628.050 28.050 ;
        RECT 544.950 26.400 628.050 27.600 ;
        RECT 544.950 25.950 547.050 26.400 ;
        RECT 607.950 25.950 610.050 26.400 ;
        RECT 625.950 25.950 628.050 26.400 ;
        RECT 637.950 27.600 640.050 28.050 ;
        RECT 730.950 27.600 733.050 28.050 ;
        RECT 637.950 26.400 733.050 27.600 ;
        RECT 637.950 25.950 640.050 26.400 ;
        RECT 730.950 25.950 733.050 26.400 ;
        RECT 70.950 24.600 73.050 25.050 ;
        RECT 112.950 24.600 115.050 25.050 ;
        RECT 70.950 23.400 115.050 24.600 ;
        RECT 70.950 22.950 73.050 23.400 ;
        RECT 112.950 22.950 115.050 23.400 ;
        RECT 247.950 24.600 250.050 25.050 ;
        RECT 301.950 24.600 304.050 25.050 ;
        RECT 337.950 24.600 340.050 25.050 ;
        RECT 247.950 23.400 304.050 24.600 ;
        RECT 247.950 22.950 250.050 23.400 ;
        RECT 301.950 22.950 304.050 23.400 ;
        RECT 305.400 23.400 340.050 24.600 ;
        RECT 305.400 22.050 306.600 23.400 ;
        RECT 337.950 22.950 340.050 23.400 ;
        RECT 340.950 24.600 343.050 25.050 ;
        RECT 349.950 24.600 352.050 25.050 ;
        RECT 340.950 23.400 352.050 24.600 ;
        RECT 340.950 22.950 343.050 23.400 ;
        RECT 349.950 22.950 352.050 23.400 ;
        RECT 361.950 24.600 364.050 25.050 ;
        RECT 388.950 24.600 391.050 25.050 ;
        RECT 361.950 23.400 391.050 24.600 ;
        RECT 361.950 22.950 364.050 23.400 ;
        RECT 388.950 22.950 391.050 23.400 ;
        RECT 430.950 24.600 433.050 25.050 ;
        RECT 481.950 24.600 484.050 25.050 ;
        RECT 430.950 23.400 484.050 24.600 ;
        RECT 430.950 22.950 433.050 23.400 ;
        RECT 481.950 22.950 484.050 23.400 ;
        RECT 34.950 21.600 37.050 22.050 ;
        RECT 154.950 21.600 157.050 22.050 ;
        RECT 34.950 20.400 157.050 21.600 ;
        RECT 34.950 19.950 37.050 20.400 ;
        RECT 154.950 19.950 157.050 20.400 ;
        RECT 304.950 19.950 307.050 22.050 ;
        RECT 310.950 21.600 313.050 22.050 ;
        RECT 316.950 21.600 319.050 22.050 ;
        RECT 310.950 20.400 319.050 21.600 ;
        RECT 310.950 19.950 313.050 20.400 ;
        RECT 316.950 19.950 319.050 20.400 ;
        RECT 349.950 21.600 352.050 22.050 ;
        RECT 382.950 21.600 385.050 22.050 ;
        RECT 466.950 21.600 469.050 22.050 ;
        RECT 349.950 20.400 385.050 21.600 ;
        RECT 349.950 19.950 352.050 20.400 ;
        RECT 382.950 19.950 385.050 20.400 ;
        RECT 386.400 20.400 469.050 21.600 ;
        RECT 313.950 18.600 316.050 19.050 ;
        RECT 386.400 18.600 387.600 20.400 ;
        RECT 466.950 19.950 469.050 20.400 ;
        RECT 535.950 21.600 538.050 22.050 ;
        RECT 541.950 21.600 544.050 22.050 ;
        RECT 535.950 20.400 544.050 21.600 ;
        RECT 535.950 19.950 538.050 20.400 ;
        RECT 541.950 19.950 544.050 20.400 ;
        RECT 547.950 21.600 550.050 22.050 ;
        RECT 586.950 21.600 589.050 22.050 ;
        RECT 616.950 21.600 619.050 22.050 ;
        RECT 547.950 20.400 619.050 21.600 ;
        RECT 547.950 19.950 550.050 20.400 ;
        RECT 586.950 19.950 589.050 20.400 ;
        RECT 616.950 19.950 619.050 20.400 ;
        RECT 628.950 21.600 631.050 22.050 ;
        RECT 697.950 21.600 700.050 22.050 ;
        RECT 628.950 20.400 700.050 21.600 ;
        RECT 628.950 19.950 631.050 20.400 ;
        RECT 697.950 19.950 700.050 20.400 ;
        RECT 313.950 17.400 387.600 18.600 ;
        RECT 469.950 18.600 472.050 19.050 ;
        RECT 481.950 18.600 484.050 19.050 ;
        RECT 469.950 17.400 484.050 18.600 ;
        RECT 313.950 16.950 316.050 17.400 ;
        RECT 469.950 16.950 472.050 17.400 ;
        RECT 481.950 16.950 484.050 17.400 ;
        RECT 511.950 18.600 514.050 19.050 ;
        RECT 589.950 18.600 592.050 19.050 ;
        RECT 637.950 18.600 640.050 19.050 ;
        RECT 511.950 17.400 640.050 18.600 ;
        RECT 511.950 16.950 514.050 17.400 ;
        RECT 589.950 16.950 592.050 17.400 ;
        RECT 637.950 16.950 640.050 17.400 ;
        RECT 661.950 18.600 664.050 19.050 ;
        RECT 694.950 18.600 697.050 19.050 ;
        RECT 661.950 17.400 697.050 18.600 ;
        RECT 661.950 16.950 664.050 17.400 ;
        RECT 694.950 16.950 697.050 17.400 ;
        RECT 700.950 18.600 703.050 19.050 ;
        RECT 733.950 18.600 736.050 19.050 ;
        RECT 700.950 17.400 736.050 18.600 ;
        RECT 700.950 16.950 703.050 17.400 ;
        RECT 733.950 16.950 736.050 17.400 ;
  END
END phase_accumulator
END LIBRARY

