magic
tech scmos
magscale 1 6
timestamp 1569533753
<< checkpaint >>
rect -120 -120 2520 320
<< psubstratepdiff >>
rect 0 0 2400 200
<< metal1 >>
rect 0 0 2400 200
use CONT$4  CONT$4_0
timestamp 1569533753
transform 1 0 164 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_1
timestamp 1569533753
transform 1 0 128 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_2
timestamp 1569533753
transform 1 0 92 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_3
timestamp 1569533753
transform 1 0 236 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_4
timestamp 1569533753
transform 1 0 200 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_5
timestamp 1569533753
transform 1 0 164 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_6
timestamp 1569533753
transform 1 0 524 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_7
timestamp 1569533753
transform 1 0 488 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_8
timestamp 1569533753
transform 1 0 452 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_9
timestamp 1569533753
transform 1 0 416 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_10
timestamp 1569533753
transform 1 0 380 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_11
timestamp 1569533753
transform 1 0 344 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_12
timestamp 1569533753
transform 1 0 308 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_13
timestamp 1569533753
transform 1 0 272 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_14
timestamp 1569533753
transform 1 0 596 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_15
timestamp 1569533753
transform 1 0 560 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_16
timestamp 1569533753
transform 1 0 524 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_17
timestamp 1569533753
transform 1 0 488 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_18
timestamp 1569533753
transform 1 0 452 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_19
timestamp 1569533753
transform 1 0 416 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_20
timestamp 1569533753
transform 1 0 380 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_21
timestamp 1569533753
transform 1 0 344 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_22
timestamp 1569533753
transform 1 0 308 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_23
timestamp 1569533753
transform 1 0 272 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_24
timestamp 1569533753
transform 1 0 236 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_25
timestamp 1569533753
transform 1 0 200 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_26
timestamp 1569533753
transform 1 0 164 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_27
timestamp 1569533753
transform 1 0 128 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_28
timestamp 1569533753
transform 1 0 236 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_29
timestamp 1569533753
transform 1 0 200 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_30
timestamp 1569533753
transform 1 0 596 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_31
timestamp 1569533753
transform 1 0 596 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_32
timestamp 1569533753
transform 1 0 560 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_33
timestamp 1569533753
transform 1 0 524 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_34
timestamp 1569533753
transform 1 0 488 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_35
timestamp 1569533753
transform 1 0 452 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_36
timestamp 1569533753
transform 1 0 416 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_37
timestamp 1569533753
transform 1 0 380 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_38
timestamp 1569533753
transform 1 0 344 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_39
timestamp 1569533753
transform 1 0 596 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_40
timestamp 1569533753
transform 1 0 560 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_41
timestamp 1569533753
transform 1 0 524 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_42
timestamp 1569533753
transform 1 0 488 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_43
timestamp 1569533753
transform 1 0 452 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_44
timestamp 1569533753
transform 1 0 416 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_45
timestamp 1569533753
transform 1 0 380 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_46
timestamp 1569533753
transform 1 0 344 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_47
timestamp 1569533753
transform 1 0 308 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_48
timestamp 1569533753
transform 1 0 272 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_49
timestamp 1569533753
transform 1 0 236 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_50
timestamp 1569533753
transform 1 0 200 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_51
timestamp 1569533753
transform 1 0 164 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_52
timestamp 1569533753
transform 1 0 128 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_53
timestamp 1569533753
transform 1 0 92 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_54
timestamp 1569533753
transform 1 0 56 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_55
timestamp 1569533753
transform 1 0 92 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_56
timestamp 1569533753
transform 1 0 56 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_57
timestamp 1569533753
transform 1 0 56 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_58
timestamp 1569533753
transform 1 0 56 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_59
timestamp 1569533753
transform 1 0 308 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_60
timestamp 1569533753
transform 1 0 272 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_61
timestamp 1569533753
transform 1 0 236 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_62
timestamp 1569533753
transform 1 0 200 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_63
timestamp 1569533753
transform 1 0 164 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_64
timestamp 1569533753
transform 1 0 128 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_65
timestamp 1569533753
transform 1 0 92 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_66
timestamp 1569533753
transform 1 0 56 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_67
timestamp 1569533753
transform 1 0 128 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_68
timestamp 1569533753
transform 1 0 92 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_69
timestamp 1569533753
transform 1 0 560 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_70
timestamp 1569533753
transform 1 0 596 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_71
timestamp 1569533753
transform 1 0 560 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_72
timestamp 1569533753
transform 1 0 524 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_73
timestamp 1569533753
transform 1 0 488 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_74
timestamp 1569533753
transform 1 0 452 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_75
timestamp 1569533753
transform 1 0 416 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_76
timestamp 1569533753
transform 1 0 380 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_77
timestamp 1569533753
transform 1 0 344 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_78
timestamp 1569533753
transform 1 0 308 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_79
timestamp 1569533753
transform 1 0 272 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_80
timestamp 1569533753
transform 1 0 1172 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_81
timestamp 1569533753
transform 1 0 1136 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_82
timestamp 1569533753
transform 1 0 920 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_83
timestamp 1569533753
transform 1 0 884 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_84
timestamp 1569533753
transform 1 0 848 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_85
timestamp 1569533753
transform 1 0 812 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_86
timestamp 1569533753
transform 1 0 776 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_87
timestamp 1569533753
transform 1 0 740 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_88
timestamp 1569533753
transform 1 0 704 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_89
timestamp 1569533753
transform 1 0 668 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_90
timestamp 1569533753
transform 1 0 776 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_91
timestamp 1569533753
transform 1 0 1172 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_92
timestamp 1569533753
transform 1 0 1136 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_93
timestamp 1569533753
transform 1 0 920 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_94
timestamp 1569533753
transform 1 0 884 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_95
timestamp 1569533753
transform 1 0 848 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_96
timestamp 1569533753
transform 1 0 812 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_97
timestamp 1569533753
transform 1 0 776 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_98
timestamp 1569533753
transform 1 0 740 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_99
timestamp 1569533753
transform 1 0 704 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_100
timestamp 1569533753
transform 1 0 668 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_101
timestamp 1569533753
transform 1 0 740 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_102
timestamp 1569533753
transform 1 0 1172 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_103
timestamp 1569533753
transform 1 0 1136 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_104
timestamp 1569533753
transform 1 0 920 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_105
timestamp 1569533753
transform 1 0 884 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_106
timestamp 1569533753
transform 1 0 848 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_107
timestamp 1569533753
transform 1 0 812 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_108
timestamp 1569533753
transform 1 0 776 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_109
timestamp 1569533753
transform 1 0 740 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_110
timestamp 1569533753
transform 1 0 704 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_111
timestamp 1569533753
transform 1 0 668 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_112
timestamp 1569533753
transform 1 0 704 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_113
timestamp 1569533753
transform 1 0 1172 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_114
timestamp 1569533753
transform 1 0 1136 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_115
timestamp 1569533753
transform 1 0 920 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_116
timestamp 1569533753
transform 1 0 884 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_117
timestamp 1569533753
transform 1 0 848 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_118
timestamp 1569533753
transform 1 0 812 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_119
timestamp 1569533753
transform 1 0 776 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_120
timestamp 1569533753
transform 1 0 740 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_121
timestamp 1569533753
transform 1 0 704 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_122
timestamp 1569533753
transform 1 0 668 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_123
timestamp 1569533753
transform 1 0 668 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_124
timestamp 1569533753
transform 1 0 1172 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_125
timestamp 1569533753
transform 1 0 1136 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_126
timestamp 1569533753
transform 1 0 920 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_127
timestamp 1569533753
transform 1 0 884 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_128
timestamp 1569533753
transform 1 0 848 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_129
timestamp 1569533753
transform 1 0 812 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_130
timestamp 1569533753
transform 1 0 632 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_131
timestamp 1569533753
transform 1 0 632 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_132
timestamp 1569533753
transform 1 0 632 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_133
timestamp 1569533753
transform 1 0 632 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_134
timestamp 1569533753
transform 1 0 632 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_135
timestamp 1569533753
transform 1 0 1388 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_136
timestamp 1569533753
transform 1 0 1352 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_137
timestamp 1569533753
transform 1 0 1316 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_138
timestamp 1569533753
transform 1 0 1280 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_139
timestamp 1569533753
transform 1 0 1244 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_140
timestamp 1569533753
transform 1 0 1316 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_141
timestamp 1569533753
transform 1 0 1748 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_142
timestamp 1569533753
transform 1 0 1532 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_143
timestamp 1569533753
transform 1 0 1496 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_144
timestamp 1569533753
transform 1 0 1460 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_145
timestamp 1569533753
transform 1 0 1424 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_146
timestamp 1569533753
transform 1 0 1388 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_147
timestamp 1569533753
transform 1 0 1352 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_148
timestamp 1569533753
transform 1 0 1316 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_149
timestamp 1569533753
transform 1 0 1280 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_150
timestamp 1569533753
transform 1 0 1244 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_151
timestamp 1569533753
transform 1 0 1244 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_152
timestamp 1569533753
transform 1 0 1748 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_153
timestamp 1569533753
transform 1 0 1532 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_154
timestamp 1569533753
transform 1 0 1496 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_155
timestamp 1569533753
transform 1 0 1460 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_156
timestamp 1569533753
transform 1 0 1424 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_157
timestamp 1569533753
transform 1 0 1388 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_158
timestamp 1569533753
transform 1 0 1352 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_159
timestamp 1569533753
transform 1 0 1316 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_160
timestamp 1569533753
transform 1 0 1280 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_161
timestamp 1569533753
transform 1 0 1244 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_162
timestamp 1569533753
transform 1 0 1352 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_163
timestamp 1569533753
transform 1 0 1532 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_164
timestamp 1569533753
transform 1 0 1496 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_165
timestamp 1569533753
transform 1 0 1460 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_166
timestamp 1569533753
transform 1 0 1424 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_167
timestamp 1569533753
transform 1 0 1388 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_168
timestamp 1569533753
transform 1 0 1748 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_169
timestamp 1569533753
transform 1 0 1748 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_170
timestamp 1569533753
transform 1 0 1532 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_171
timestamp 1569533753
transform 1 0 1496 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_172
timestamp 1569533753
transform 1 0 1460 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_173
timestamp 1569533753
transform 1 0 1424 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_174
timestamp 1569533753
transform 1 0 1388 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_175
timestamp 1569533753
transform 1 0 1352 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_176
timestamp 1569533753
transform 1 0 1316 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_177
timestamp 1569533753
transform 1 0 1280 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_178
timestamp 1569533753
transform 1 0 1244 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_179
timestamp 1569533753
transform 1 0 1280 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_180
timestamp 1569533753
transform 1 0 1748 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_181
timestamp 1569533753
transform 1 0 1532 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_182
timestamp 1569533753
transform 1 0 1496 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_183
timestamp 1569533753
transform 1 0 1460 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_184
timestamp 1569533753
transform 1 0 1424 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_185
timestamp 1569533753
transform 1 0 2360 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_186
timestamp 1569533753
transform 1 0 2324 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_187
timestamp 1569533753
transform 1 0 2288 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_188
timestamp 1569533753
transform 1 0 2252 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_189
timestamp 1569533753
transform 1 0 2216 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_190
timestamp 1569533753
transform 1 0 2180 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_191
timestamp 1569533753
transform 1 0 2144 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_192
timestamp 1569533753
transform 1 0 2108 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_193
timestamp 1569533753
transform 1 0 2072 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_194
timestamp 1569533753
transform 1 0 2036 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_195
timestamp 1569533753
transform 1 0 2000 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_196
timestamp 1569533753
transform 1 0 1964 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_197
timestamp 1569533753
transform 1 0 1928 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_198
timestamp 1569533753
transform 1 0 1892 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_199
timestamp 1569533753
transform 1 0 1856 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_200
timestamp 1569533753
transform 1 0 1820 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_201
timestamp 1569533753
transform 1 0 1928 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_202
timestamp 1569533753
transform 1 0 2360 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_203
timestamp 1569533753
transform 1 0 2324 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_204
timestamp 1569533753
transform 1 0 2288 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_205
timestamp 1569533753
transform 1 0 2252 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_206
timestamp 1569533753
transform 1 0 2216 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_207
timestamp 1569533753
transform 1 0 2180 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_208
timestamp 1569533753
transform 1 0 2144 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_209
timestamp 1569533753
transform 1 0 2108 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_210
timestamp 1569533753
transform 1 0 2072 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_211
timestamp 1569533753
transform 1 0 2036 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_212
timestamp 1569533753
transform 1 0 2000 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_213
timestamp 1569533753
transform 1 0 1964 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_214
timestamp 1569533753
transform 1 0 1928 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_215
timestamp 1569533753
transform 1 0 1892 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_216
timestamp 1569533753
transform 1 0 1856 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_217
timestamp 1569533753
transform 1 0 1820 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_218
timestamp 1569533753
transform 1 0 1892 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_219
timestamp 1569533753
transform 1 0 2360 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_220
timestamp 1569533753
transform 1 0 2324 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_221
timestamp 1569533753
transform 1 0 2288 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_222
timestamp 1569533753
transform 1 0 2252 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_223
timestamp 1569533753
transform 1 0 2216 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_224
timestamp 1569533753
transform 1 0 2180 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_225
timestamp 1569533753
transform 1 0 2144 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_226
timestamp 1569533753
transform 1 0 2108 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_227
timestamp 1569533753
transform 1 0 2072 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_228
timestamp 1569533753
transform 1 0 2036 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_229
timestamp 1569533753
transform 1 0 2000 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_230
timestamp 1569533753
transform 1 0 1964 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_231
timestamp 1569533753
transform 1 0 1928 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_232
timestamp 1569533753
transform 1 0 1892 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_233
timestamp 1569533753
transform 1 0 1856 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_234
timestamp 1569533753
transform 1 0 1820 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_235
timestamp 1569533753
transform 1 0 1856 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_236
timestamp 1569533753
transform 1 0 2360 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_237
timestamp 1569533753
transform 1 0 2324 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_238
timestamp 1569533753
transform 1 0 2288 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_239
timestamp 1569533753
transform 1 0 2252 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_240
timestamp 1569533753
transform 1 0 2216 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_241
timestamp 1569533753
transform 1 0 2180 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_242
timestamp 1569533753
transform 1 0 2144 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_243
timestamp 1569533753
transform 1 0 2108 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_244
timestamp 1569533753
transform 1 0 2072 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_245
timestamp 1569533753
transform 1 0 2036 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_246
timestamp 1569533753
transform 1 0 2000 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_247
timestamp 1569533753
transform 1 0 1964 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_248
timestamp 1569533753
transform 1 0 1928 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_249
timestamp 1569533753
transform 1 0 1892 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_250
timestamp 1569533753
transform 1 0 1856 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_251
timestamp 1569533753
transform 1 0 1820 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_252
timestamp 1569533753
transform 1 0 1820 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_253
timestamp 1569533753
transform 1 0 2360 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_254
timestamp 1569533753
transform 1 0 2324 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_255
timestamp 1569533753
transform 1 0 2288 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_256
timestamp 1569533753
transform 1 0 2252 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_257
timestamp 1569533753
transform 1 0 2216 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_258
timestamp 1569533753
transform 1 0 2180 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_259
timestamp 1569533753
transform 1 0 2144 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_260
timestamp 1569533753
transform 1 0 2108 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_261
timestamp 1569533753
transform 1 0 2072 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_262
timestamp 1569533753
transform 1 0 2036 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_263
timestamp 1569533753
transform 1 0 2000 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_264
timestamp 1569533753
transform 1 0 1964 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_265
timestamp 1569533753
transform 1 0 1784 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_266
timestamp 1569533753
transform 1 0 1784 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_267
timestamp 1569533753
transform 1 0 1784 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_268
timestamp 1569533753
transform 1 0 1784 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_269
timestamp 1569533753
transform 1 0 1784 0 1 27
box -6 -6 6 6
use CONT$4  CONT$4_270
timestamp 1569533753
transform 1 0 1208 0 1 171
box -6 -6 6 6
use CONT$4  CONT$4_271
timestamp 1569533753
transform 1 0 1208 0 1 135
box -6 -6 6 6
use CONT$4  CONT$4_272
timestamp 1569533753
transform 1 0 1208 0 1 99
box -6 -6 6 6
use CONT$4  CONT$4_273
timestamp 1569533753
transform 1 0 1208 0 1 63
box -6 -6 6 6
use CONT$4  CONT$4_274
timestamp 1569533753
transform 1 0 1208 0 1 27
box -6 -6 6 6
<< end >>
