/* Verilog module written by vlogFanout (qflow) */
/* With clock tree generation and fanout reduction */
/* and gate resizing */

module DDFS(
    output [11:0] Dout,
    input En,
    input [19:0] FCW,
    output Vld,
    input clk,
    input selXY
);

wire _4972_ ;
wire _4552_ ;
wire _4132_ ;
wire _5757_ ;
wire _5337_ ;
wire _1677_ ;
wire _1257_ ;
wire _5090_ ;
wire _588_ ;
wire _168_ ;
wire _3823_ ;
wire _3403_ ;
wire _6295_ ;
wire _4608_ ;
wire _4781_ ;
wire _4361_ ;
wire _800_ ;
wire _5986_ ;
wire _5566_ ;
wire _5146_ ;
wire _60_ ;
wire _1486_ ;
wire _1066_ ;
wire _397_ ;
wire _3632_ ;
wire _3212_ ;
wire _4837_ ;
wire _4417_ ;
wire _4590_ ;
wire _4170_ ;
wire _2903_ ;
wire _5795_ ;
wire _5375_ ;
wire _1295_ ;
wire _3861_ ;
wire _3441_ ;
wire _3021_ ;
wire _4646_ ;
wire _4226_ ;
wire \genblk1[0].u_ce.Vld_bF$buf4  ;
wire _2712_ ;
wire _5184_ ;
wire _3917_ ;
wire [1:0] \a[5]  ;
wire _3670_ ;
wire _3250_ ;
wire _4875_ ;
wire _4455_ ;
wire _4035_ ;
wire _2941_ ;
wire _2521_ ;
wire _2101_ ;
wire _3726_ ;
wire _3306_ ;
wire _6198_ ;
wire _4684_ ;
wire _4264_ ;
wire _703_ ;
wire _5889_ ;
wire _5469_ ;
wire _5049_ ;
wire _1389_ ;
wire _2750_ ;
wire _2330_ ;
wire _3955_ ;
wire _3535_ ;
wire _3115_ ;
wire \genblk1[2].u_ce.Vld_bF$buf0  ;
wire [1:0] \genblk1[2].u_ce.Y_  ;
wire _19_ ;
wire _1601_ ;
wire _4493_ ;
wire _4073_ ;
wire _932_ ;
wire _512_ ;
wire _2806_ ;
wire _5698_ ;
wire _5278_ ;
wire _1198_ ;
wire _3764_ ;
wire _3344_ ;
wire _4969_ ;
wire _4549_ ;
wire _4129_ ;
wire _5910_ ;
wire _1830_ ;
wire _1410_ ;
wire _741_ ;
wire _321_ ;
wire _2615_ ;
wire _5087_ ;
wire _3993_ ;
wire _3573_ ;
wire _3153_ ;
wire _4778_ ;
wire _4358_ ;
wire _57_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _2844_ ;
wire [1:0] \genblk1[5].u_ce.Yin0  ;
wire _2424_ ;
wire _2004_ ;
wire _3629_ ;
wire _3209_ ;
wire _3382_ ;
wire _4587_ ;
wire _4167_ ;
wire _606_ ;
wire _6313_ ;
wire _2653_ ;
wire _2233_ ;
wire _3858_ ;
wire _3438_ ;
wire _3018_ ;
wire _3191_ ;
wire _1924_ ;
wire _1504_ ;
wire _4396_ ;
wire _835_ ;
wire _415_ ;
wire _2709_ ;
wire _95_ ;
wire _6122_ ;
wire _2882_ ;
wire _2462_ ;
wire _2042_ ;
wire _3667_ ;
wire _3247_ ;
wire _5813_ ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _2938_ ;
wire _2518_ ;
wire _2691_ ;
wire _2271_ ;
wire _3896_ ;
wire _3476_ ;
wire _3056_ ;
wire _5622_ ;
wire _5202_ ;
wire _1962_ ;
wire _1542_ ;
wire \genblk1[4].u_ce.Ain12b_11_bF$buf1  ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _2747_ ;
wire _2327_ ;
wire _6160_ ;
wire _2080_ ;
wire _3285_ ;
wire _5851_ ;
wire _5431_ ;
wire _5011_ ;
wire _929_ ;
wire _509_ ;
wire _6216_ ;
wire _1771_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _2976_ ;
wire _2556_ ;
wire _2136_ ;
wire _4702_ ;
wire _5907_ ;
wire _3094_ ;
wire \genblk1[1].u_ce.LoadCtl_0_bF$buf2  ;
wire _1827_ ;
wire _1407_ ;
wire _4299_ ;
wire _5660_ ;
wire _5240_ ;
wire _738_ ;
wire _318_ ;
wire _6025_ ;
wire _1580_ ;
wire _1160_ ;
wire _491_ ;
wire _2785_ ;
wire _2365_ ;
wire _4931_ ;
wire _4511_ ;
wire _5716_ ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _6254_ ;
wire _2594_ ;
wire _2174_ ;
wire _3799_ ;
wire _3379_ ;
wire _4740_ ;
wire _4320_ ;
wire _5945_ ;
wire _5525_ ;
wire _5105_ ;
wire _1865_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _6063_ ;
wire _3188_ ;
wire _5754_ ;
wire _5334_ ;
wire _6119_ ;
wire _1674_ ;
wire _1254_ ;
wire [1:0] \genblk1[2].u_ce.Xin1  ;
wire _585_ ;
wire _165_ ;
wire _2879_ ;
wire _2459_ ;
wire _2039_ ;
wire _3820_ ;
wire _3400_ ;
wire _6292_ ;
wire _4605_ ;
wire _5983_ ;
wire _5563_ ;
wire _5143_ ;
wire [11:0] _6348_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _2688_ ;
wire _2268_ ;
wire _4834_ ;
wire _4414_ ;
wire _5619_ ;
wire _1959_ ;
wire _1539_ ;
wire _1119_ ;
wire _2900_ ;
wire _5792_ ;
wire _5372_ ;
wire _6157_ ;
wire _1292_ ;
wire _2497_ ;
wire _2077_ ;
wire _4643_ ;
wire _4223_ ;
wire _5848_ ;
wire _5428_ ;
wire _5008_ ;
wire \genblk1[0].u_ce.Vld_bF$buf1  ;
wire _1768_ ;
wire _1348_ ;
wire _5181_ ;
wire _679_ ;
wire _259_ ;
wire _3914_ ;
wire _4872_ ;
wire _4452_ ;
wire _4032_ ;
wire _5657_ ;
wire _5237_ ;
wire _1997_ ;
wire _1577_ ;
wire _1157_ ;
wire _488_ ;
wire _3723_ ;
wire _3303_ ;
wire _6195_ ;
wire _4928_ ;
wire _4508_ ;
wire _4681_ ;
wire _4261_ ;
wire _700_ ;
wire _5886_ ;
wire _5466_ ;
wire _5046_ ;
wire _1386_ ;
wire _297_ ;
wire _3952_ ;
wire _3532_ ;
wire _3112_ ;
wire _4737_ ;
wire _4317_ ;
wire _16_ ;
wire _4490_ ;
wire _4070_ ;
wire _2803_ ;
wire _5695_ ;
wire _5275_ ;
wire _1195_ ;
wire [11:0] \u_pa.Atmp  ;
wire _3761_ ;
wire _3341_ ;
wire _4966_ ;
wire _4546_ ;
wire _4126_ ;
wire _3655__bF$buf0 ;
wire _3655__bF$buf1 ;
wire _3655__bF$buf2 ;
wire _3655__bF$buf3 ;
wire _2612_ ;
wire _5084_ ;
wire _3817_ ;
wire _6289_ ;
wire _3990_ ;
wire _3570_ ;
wire _3150_ ;
wire _4775_ ;
wire _4355_ ;
wire _54_ ;
wire _2841_ ;
wire _2421_ ;
wire _2001_ ;
wire _3626_ ;
wire _3206_ ;
wire _6098_ ;
wire _4584_ ;
wire _4164_ ;
wire _603_ ;
wire _5789_ ;
wire _5369_ ;
wire _6310_ ;
wire _1289_ ;
wire _2650_ ;
wire _2230_ ;
wire \u_ot.ISout_bF$buf2  ;
wire \genblk1[2].u_ce.Ain12b_11_bF$buf4  ;
wire _3855_ ;
wire _3435_ ;
wire _3015_ ;
wire _1921_ ;
wire _1501_ ;
wire _4393_ ;
wire _832_ ;
wire _412_ ;
wire _2706_ ;
wire _5598_ ;
wire _5178_ ;
wire _92_ ;
wire _1098_ ;
wire _3664_ ;
wire _3244_ ;
wire _4869_ ;
wire _4449_ ;
wire _4029_ ;
wire _5810_ ;
wire _1730_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _2935_ ;
wire _2515_ ;
wire _4480__bF$buf0 ;
wire _4480__bF$buf1 ;
wire _4480__bF$buf2 ;
wire _4480__bF$buf3 ;
wire _4480__bF$buf4 ;
wire _3893_ ;
wire _3473_ ;
wire _3053_ ;
wire _4678_ ;
wire _4258_ ;
wire _870_ ;
wire _450_ ;
wire _2744_ ;
wire _2324_ ;
wire _3949_ ;
wire _3529_ ;
wire _3109_ ;
wire _3282_ ;
wire _4487_ ;
wire _4067_ ;
wire _926_ ;
wire _506_ ;
wire _6213_ ;
wire _2973_ ;
wire _2553_ ;
wire _2133_ ;
wire _3758_ ;
wire _3338_ ;
wire \genblk1[2].u_ce.ISout  ;
wire _5904_ ;
wire _3091_ ;
wire _1824_ ;
wire _1404_ ;
wire _4296_ ;
wire _735_ ;
wire _315_ ;
wire _2609_ ;
wire _6022_ ;
wire _2782_ ;
wire _2362_ ;
wire _3987_ ;
wire _3567_ ;
wire _3147_ ;
wire _5713_ ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire _2838_ ;
wire _2418_ ;
wire _6251_ ;
wire _2591_ ;
wire _2171_ ;
wire _3796_ ;
wire _3376_ ;
wire [11:0] \genblk1[5].u_ce.Xcalc  ;
wire _5942_ ;
wire _5522_ ;
wire _5102_ ;
wire _6307_ ;
wire _1862_ ;
wire _1442_ ;
wire _1022_ ;
wire _773_ ;
wire _353_ ;
wire _2647_ ;
wire _2227_ ;
wire _6060_ ;
wire [6:0] \genblk1[5].u_ce.ISpipe  ;
wire _3185_ ;
wire _1918_ ;
wire _5751_ ;
wire _5331_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _6116_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _2876_ ;
wire _2456_ ;
wire _2036_ ;
wire _4602_ ;
wire _5807_ ;
wire _1727_ ;
wire _1307_ ;
wire _4199_ ;
wire _5980_ ;
wire _5560_ ;
wire _5140_ ;
wire _638_ ;
wire _218_ ;
wire _6345_ ;
wire _1480_ ;
wire _1060_ ;
wire _1030__bF$buf0 ;
wire _391_ ;
wire _1030__bF$buf1 ;
wire _1030__bF$buf2 ;
wire _1030__bF$buf3 ;
wire _1030__bF$buf4 ;
wire _2685_ ;
wire _2265_ ;
wire _4831_ ;
wire _4411_ ;
wire _5616_ ;
wire _1956_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _6154_ ;
wire _2494_ ;
wire _2074_ ;
wire _3699_ ;
wire _3279_ ;
wire _4640_ ;
wire _4220_ ;
wire [11:0] _5845_ ;
wire _5425_ ;
wire _5005_ ;
wire _1765_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _3911_ ;
wire _3088_ ;
wire _5654_ ;
wire _5234_ ;
wire _6019_ ;
wire _1994_ ;
wire _1574_ ;
wire _1154_ ;
wire _485_ ;
wire _2779_ ;
wire _2359_ ;
wire _3720_ ;
wire _3300_ ;
wire _6192_ ;
wire \genblk1[6].u_ce.LoadCtl_0_bF$buf2  ;
wire _4925_ ;
wire _4505_ ;
wire \genblk1[5].u_ce.Vld_bF$buf2  ;
wire _5883_ ;
wire _5463_ ;
wire _5043_ ;
wire _6248_ ;
wire _1383_ ;
wire _294_ ;
wire _2588_ ;
wire _2168_ ;
wire _4734_ ;
wire _4314_ ;
wire _5939_ ;
wire _5519_ ;
wire _13_ ;
wire _1859_ ;
wire _1439_ ;
wire _1019_ ;
wire _2800_ ;
wire _5692_ ;
wire _5272_ ;
wire _6057_ ;
wire _1192_ ;
wire _2397_ ;
wire _4963_ ;
wire _4543_ ;
wire _4123_ ;
wire _5748_ ;
wire _5328_ ;
wire _1668_ ;
wire _1248_ ;
wire _5081_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _3814_ ;
wire _6286_ ;
wire _4772_ ;
wire _4352_ ;
wire _2789__bF$buf0 ;
wire _2789__bF$buf1 ;
wire _2789__bF$buf2 ;
wire _2789__bF$buf3 ;
wire _5977_ ;
wire _5557_ ;
wire _5137_ ;
wire _51_ ;
wire _1897_ ;
wire _1477_ ;
wire _1057_ ;
wire _388_ ;
wire _3623_ ;
wire _3203_ ;
wire _6095_ ;
wire _4828_ ;
wire _4408_ ;
wire _4581_ ;
wire _4161_ ;
wire _600_ ;
wire _5786_ ;
wire _5366_ ;
wire _1286_ ;
wire _197_ ;
wire \genblk1[2].u_ce.Ain12b_11_bF$buf1  ;
wire _3852_ ;
wire _3432_ ;
wire _3012_ ;
wire _4637_ ;
wire _4217_ ;
wire _4390_ ;
wire _2703_ ;
wire _5595_ ;
wire _5175_ ;
wire _3908_ ;
wire _1095_ ;
wire _3661_ ;
wire _3241_ ;
wire _4866_ ;
wire _4446_ ;
wire _4026_ ;
wire _2932_ ;
wire _2512_ ;
wire _3717_ ;
wire _6189_ ;
wire _3890_ ;
wire _3470_ ;
wire _3050_ ;
wire _4675_ ;
wire _4255_ ;
wire _2741_ ;
wire _2321_ ;
wire _3946_ ;
wire _3526_ ;
wire _3106_ ;
wire _7_ ;
wire [11:0] \u_ot.Xcalc  ;
wire _4484_ ;
wire _4064_ ;
wire _923_ ;
wire _503_ ;
wire _5689_ ;
wire _5269_ ;
wire _6210_ ;
wire [1:0] \genblk1[0].u_ce.Ain1  ;
wire _1189_ ;
wire _2970_ ;
wire _2550_ ;
wire _2130_ ;
wire [1:0] \genblk1[3].u_ce.Y_  ;
wire _3755_ ;
wire _3335_ ;
wire _5901_ ;
wire _1821_ ;
wire _1401_ ;
wire _4293_ ;
wire _732_ ;
wire _312_ ;
wire _2606_ ;
wire _5498_ ;
wire _5078_ ;
wire _3984_ ;
wire _3564_ ;
wire _3144_ ;
wire _4769_ ;
wire _4349_ ;
wire _5710_ ;
wire _48_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _2835_ ;
wire _2415_ ;
wire _3793_ ;
wire _3373_ ;
wire _4998_ ;
wire _4578_ ;
wire _4158_ ;
wire \genblk1[4].u_ce.LoadCtl_0_bF$buf3  ;
wire _6304_ ;
wire _770_ ;
wire _350_ ;
wire _2644_ ;
wire _2224_ ;
wire _3849_ ;
wire _3429_ ;
wire _3009_ ;
wire _3182_ ;
wire _1915_ ;
wire _4387_ ;
wire [11:0] \genblk1[0].u_ce.Yin12b  ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _6113_ ;
wire [1:0] \genblk1[1].u_ce.Xin0  ;
wire _2873_ ;
wire _2453_ ;
wire _2033_ ;
wire _3658_ ;
wire _3238_ ;
wire _5804_ ;
wire _1724_ ;
wire _1304_ ;
wire _4196_ ;
wire _635_ ;
wire _215_ ;
wire _2929_ ;
wire _2509_ ;
wire _6342_ ;
wire _2682_ ;
wire _2262_ ;
wire _158__bF$buf0 ;
wire _158__bF$buf1 ;
wire _158__bF$buf2 ;
wire _158__bF$buf3 ;
wire _158__bF$buf4 ;
wire _3887_ ;
wire _3467_ ;
wire _3047_ ;
wire _5613_ ;
wire _1953_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _2738_ ;
wire _2318_ ;
wire _6151_ ;
wire _2491_ ;
wire _2071_ ;
wire _3696_ ;
wire _3276_ ;
wire _5842_ ;
wire _5422_ ;
wire _5002_ ;
wire _6207_ ;
wire _1762_ ;
wire _1342_ ;
wire _673_ ;
wire _253_ ;
wire _2967_ ;
wire _2547_ ;
wire _2127_ ;
wire _3085_ ;
wire _1818_ ;
wire _5651_ ;
wire _5231_ ;
wire _729_ ;
wire _309_ ;
wire [11:0] \genblk1[2].u_ce.Yin12b  ;
wire _6016_ ;
wire _1991_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _2776_ ;
wire _2356_ ;
wire _4922_ ;
wire _4502_ ;
wire _5707_ ;
wire _1627_ ;
wire _1207_ ;
wire _4099_ ;
wire _5880_ ;
wire _5460_ ;
wire _5040_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _6245_ ;
wire _1380_ ;
wire _291_ ;
wire _2585_ ;
wire _2165_ ;
wire _4731_ ;
wire _4311_ ;
wire _5936_ ;
wire _5516_ ;
wire _10_ ;
wire \genblk1[2].u_ce.Vld  ;
wire _1856_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _6054_ ;
wire _2394_ ;
wire _3599_ ;
wire _3179_ ;
wire _4960_ ;
wire \genblk1[0].u_ce.Ain12b_11_bF$buf4  ;
wire _4540_ ;
wire _4120_ ;
wire _5745_ ;
wire _5325_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _3811_ ;
wire _6283_ ;
wire _5974_ ;
wire _5554_ ;
wire _5134_ ;
wire _6339_ ;
wire _1894_ ;
wire [11:0] \genblk1[4].u_ce.Yin12b  ;
wire _1474_ ;
wire _1054_ ;
wire _385_ ;
wire [1:0] \a[0]  ;
wire _2679_ ;
wire _2259_ ;
wire [1:0] \genblk1[3].u_ce.Yin1  ;
wire _3620_ ;
wire _3200_ ;
wire _6092_ ;
wire _4825_ ;
wire _4405_ ;
wire _5783_ ;
wire _5363_ ;
wire _6148_ ;
wire _1283_ ;
wire _194_ ;
wire _2488_ ;
wire _2068_ ;
wire _4634_ ;
wire _4214_ ;
wire _5839_ ;
wire _5419_ ;
wire _1759_ ;
wire _1339_ ;
wire _2700_ ;
wire _5592_ ;
wire _5172_ ;
wire _3905_ ;
wire _1092_ ;
wire _2297_ ;
wire _4863_ ;
wire _4443_ ;
wire _4023_ ;
wire _5648_ ;
wire _5228_ ;
wire _1988_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire _3714_ ;
wire _6186_ ;
wire _4919_ ;
wire _4672_ ;
wire _4252_ ;
wire [11:0] \u_ot.Yin12b  ;
wire _5877_ ;
wire _5457_ ;
wire _5037_ ;
wire _1797_ ;
wire _1377_ ;
wire [11:0] \genblk1[6].u_ce.Yin12b  ;
wire _288_ ;
wire _3943_ ;
wire _3523_ ;
wire _3103_ ;
wire _4_ ;
wire _4728_ ;
wire _4308_ ;
wire _4481_ ;
wire _4061_ ;
wire _920_ ;
wire _500_ ;
wire _5686_ ;
wire _5266_ ;
wire _1186_ ;
wire _3752_ ;
wire _3332_ ;
wire _4957_ ;
wire _4537_ ;
wire _4117_ ;
wire _4290_ ;
wire _2603_ ;
wire _5495_ ;
wire _5075_ ;
wire _3808_ ;
wire _3981_ ;
wire _3561_ ;
wire _3141_ ;
wire _4766_ ;
wire _4346_ ;
wire _45_ ;
wire _2832_ ;
wire _2412_ ;
wire _1896__bF$buf0 ;
wire _1896__bF$buf1 ;
wire _1896__bF$buf2 ;
wire _1896__bF$buf3 ;
wire _1896__bF$buf4 ;
wire _3617_ ;
wire _6089_ ;
wire _3790_ ;
wire _3370_ ;
wire _4995_ ;
wire _4575_ ;
wire _4155_ ;
wire \genblk1[4].u_ce.LoadCtl_0_bF$buf0  ;
wire _6301_ ;
wire _2641_ ;
wire _2221_ ;
wire _3846_ ;
wire _3426_ ;
wire _3006_ ;
wire _1912_ ;
wire _4384_ ;
wire _823_ ;
wire _403_ ;
wire _5589_ ;
wire _5169_ ;
wire _83_ ;
wire _6110_ ;
wire _1089_ ;
wire _2870_ ;
wire _2450_ ;
wire _2030_ ;
wire _3655_ ;
wire _3235_ ;
wire _5801_ ;
wire _1721_ ;
wire _1301_ ;
wire _4193_ ;
wire _632_ ;
wire _212_ ;
wire _2926_ ;
wire _2506_ ;
wire _5398_ ;
wire _1923__bF$buf0 ;
wire _1923__bF$buf1 ;
wire _1923__bF$buf2 ;
wire _1923__bF$buf3 ;
wire _3884_ ;
wire _3464_ ;
wire _3044_ ;
wire _4669_ ;
wire _4249_ ;
wire _5610_ ;
wire _1950_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _2735_ ;
wire _2315_ ;
wire _3693_ ;
wire _3273_ ;
wire _4898_ ;
wire _4478_ ;
wire _4058_ ;
wire _917_ ;
wire _6204_ ;
wire _670_ ;
wire _250_ ;
wire _2964_ ;
wire _2544_ ;
wire _2124_ ;
wire _3749_ ;
wire _3329_ ;
wire _3082_ ;
wire _1815_ ;
wire _4287_ ;
wire _726_ ;
wire _306_ ;
wire _6013_ ;
wire _2773_ ;
wire _2353_ ;
wire _3978_ ;
wire _3558_ ;
wire _3138_ ;
wire _5704_ ;
wire \genblk1[3].u_ce.Vld_bF$buf2  ;
wire _1624_ ;
wire _1204_ ;
wire _4096_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _2829_ ;
wire _2409_ ;
wire _6242_ ;
wire _2582_ ;
wire _2162_ ;
wire _3787_ ;
wire _3367_ ;
wire _5933_ ;
wire _5513_ ;
wire _1853_ ;
wire _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _2638_ ;
wire _2218_ ;
wire _6051_ ;
wire _2391_ ;
wire _3596_ ;
wire _3176_ ;
wire \genblk1[0].u_ce.Ain12b_11_bF$buf1  ;
wire _1909_ ;
wire _5742_ ;
wire _5322_ ;
wire _6107_ ;
wire _1662_ ;
wire _1242_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _2867_ ;
wire _2447_ ;
wire _2027_ ;
wire _6280_ ;
wire _1718_ ;
wire _5971_ ;
wire _5551_ ;
wire _5131_ ;
wire _629_ ;
wire _209_ ;
wire _6336_ ;
wire _1891_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _2676_ ;
wire _2256_ ;
wire clk_bF$buf50 ;
wire clk_bF$buf51 ;
wire clk_bF$buf52 ;
wire clk_bF$buf53 ;
wire clk_bF$buf54 ;
wire clk_bF$buf55 ;
wire clk_bF$buf56 ;
wire clk_bF$buf57 ;
wire clk_bF$buf58 ;
wire clk_bF$buf59 ;
wire _4822_ ;
wire _4402_ ;
wire _5607_ ;
wire _1947_ ;
wire _1527_ ;
wire _1107_ ;
wire _5780_ ;
wire _5360_ ;
wire _858_ ;
wire _438_ ;
wire _6145_ ;
wire _1280_ ;
wire _191_ ;
wire _2485_ ;
wire _2065_ ;
wire _4631_ ;
wire _4211_ ;
wire _5836_ ;
wire _5416_ ;
wire _1756_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _3902_ ;
wire _2294_ ;
wire _3499_ ;
wire _3079_ ;
wire _4860_ ;
wire _4440_ ;
wire _4020_ ;
wire [11:0] \genblk1[2].u_ce.Xcalc  ;
wire _5645_ ;
wire _5225_ ;
wire _1985_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire [6:0] \genblk1[1].u_ce.LoadCtl  ;
wire _476_ ;
wire _3711_ ;
wire \genblk1[5].u_ce.Ain12b_11_bF$buf2  ;
wire _6183_ ;
wire _4916_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire clk_bF$buf9 ;
wire _5874_ ;
wire _5454_ ;
wire _5034_ ;
wire _6239_ ;
wire _1794_ ;
wire _1374_ ;
wire _285_ ;
wire _2999_ ;
wire _2579_ ;
wire _2159_ ;
wire _3940_ ;
wire _3520_ ;
wire _3100_ ;
wire _1_ ;
wire _4725_ ;
wire _4305_ ;
wire [1:0] \genblk1[6].u_ce.Xin1  ;
wire _5683_ ;
wire _5263_ ;
wire \genblk1[2].u_ce.LoadCtl_0_bF$buf3  ;
wire _6048_ ;
wire _1183_ ;
wire _2388_ ;
wire _5303__bF$buf0 ;
wire _5303__bF$buf1 ;
wire _5303__bF$buf2 ;
wire _5303__bF$buf3 ;
wire _4954_ ;
wire _4534_ ;
wire _4114_ ;
wire _5739_ ;
wire _5319_ ;
wire _1659_ ;
wire _1239_ ;
wire _2600_ ;
wire _5492_ ;
wire _5072_ ;
wire _3805_ ;
wire _6277_ ;
wire _2197_ ;
wire _4763_ ;
wire _4343_ ;
wire _5968_ ;
wire _5548_ ;
wire _5128_ ;
wire _42_ ;
wire _1888_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _3614_ ;
wire _6086_ ;
wire _4819_ ;
wire _4992_ ;
wire _4572_ ;
wire _4152_ ;
wire _5777_ ;
wire _5357_ ;
wire _1697_ ;
wire _1277_ ;
wire _188_ ;
wire _3843_ ;
wire _3423_ ;
wire _3003_ ;
wire _4628_ ;
wire _4208_ ;
wire _4381_ ;
wire _820_ ;
wire _400_ ;
wire _5586_ ;
wire _5166_ ;
wire _80_ ;
wire _1086_ ;
wire _3652_ ;
wire _3232_ ;
wire _4857_ ;
wire _4437_ ;
wire _4017_ ;
wire _4190_ ;
wire _2923_ ;
wire _2503_ ;
wire _5395_ ;
wire _3708_ ;
wire _3881_ ;
wire _3461_ ;
wire _3041_ ;
wire _4666_ ;
wire _4246_ ;
wire _2732_ ;
wire _2312_ ;
wire \genblk1[1].u_ce.Vld_bF$buf3  ;
wire _3937_ ;
wire _3517_ ;
wire _3690_ ;
wire _3270_ ;
wire _4895_ ;
wire _4475_ ;
wire _4055_ ;
wire _914_ ;
wire _6201_ ;
wire _2961_ ;
wire _2541_ ;
wire _2121_ ;
wire _3746_ ;
wire _3326_ ;
wire _1812_ ;
wire _4284_ ;
wire [1:0] \genblk1[4].u_ce.Y_  ;
wire _723_ ;
wire _303_ ;
wire _5489_ ;
wire _5069_ ;
wire _6010_ ;
wire _2770_ ;
wire _2350_ ;
wire _3975_ ;
wire _3555_ ;
wire _3135_ ;
wire _5701_ ;
wire _39_ ;
wire _1621_ ;
wire _1201_ ;
wire _4093_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _2826_ ;
wire _2406_ ;
wire _5298_ ;
wire _3784_ ;
wire _3364_ ;
wire _4989_ ;
wire _4569_ ;
wire _4149_ ;
wire _5930_ ;
wire _5510_ ;
wire _1850_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire _2635_ ;
wire _2215_ ;
wire clk ;
wire _3593_ ;
wire _3173_ ;
wire _1906_ ;
wire _4798_ ;
wire _4378_ ;
wire _817_ ;
wire _77_ ;
wire _6104_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _2864_ ;
wire _2444_ ;
wire _2024_ ;
wire \genblk1[6].u_ce.ISout  ;
wire _3649_ ;
wire _3229_ ;
wire _1715_ ;
wire _4187_ ;
wire _626_ ;
wire _206_ ;
wire _6333_ ;
wire _2673_ ;
wire _2253_ ;
wire clk_bF$buf20 ;
wire clk_bF$buf21 ;
wire clk_bF$buf22 ;
wire clk_bF$buf23 ;
wire clk_bF$buf24 ;
wire clk_bF$buf25 ;
wire clk_bF$buf26 ;
wire clk_bF$buf27 ;
wire [1:0] \genblk1[2].u_ce.Yin0  ;
wire clk_bF$buf28 ;
wire clk_bF$buf29 ;
wire _3878_ ;
wire _3458_ ;
wire _3038_ ;
wire _5604_ ;
wire _1944_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _2729_ ;
wire _2309_ ;
wire _6142_ ;
wire _2482_ ;
wire _2062_ ;
wire _3687_ ;
wire _3267_ ;
wire _5833_ ;
wire _5413_ ;
wire _1753_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _2958_ ;
wire _2538_ ;
wire _2118_ ;
wire _2291_ ;
wire _3496_ ;
wire _3076_ ;
wire _1809_ ;
wire _5642_ ;
wire _5222_ ;
wire _6007_ ;
wire _1982_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _2767_ ;
wire _2347_ ;
wire _6180_ ;
wire [6:0] \u_pa.RdyCtl  ;
wire _4913_ ;
wire _1618_ ;
wire _5871_ ;
wire _5451_ ;
wire _5031_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _6236_ ;
wire _1791_ ;
wire _1371_ ;
wire _282_ ;
wire _2996_ ;
wire _2576_ ;
wire _2156_ ;
wire _4722_ ;
wire _4302_ ;
wire _5927_ ;
wire _5507_ ;
wire _1847_ ;
wire _1427_ ;
wire _1007_ ;
wire _5680_ ;
wire _5260_ ;
wire _758_ ;
wire _338_ ;
wire \genblk1[2].u_ce.LoadCtl_0_bF$buf0  ;
wire _6045_ ;
wire _1180_ ;
wire _2385_ ;
wire selXY_bF$buf0 ;
wire selXY_bF$buf1 ;
wire selXY_bF$buf2 ;
wire selXY_bF$buf3 ;
wire _4951_ ;
wire _4531_ ;
wire _4111_ ;
wire _5736_ ;
wire _5316_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _3802_ ;
wire _6274_ ;
wire _2194_ ;
wire _3399_ ;
wire _4760_ ;
wire _4340_ ;
wire _5965_ ;
wire _5545_ ;
wire _5125_ ;
wire _1885_ ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire _376_ ;
wire _3611_ ;
wire _6083_ ;
wire _4816_ ;
wire _5774_ ;
wire _5354_ ;
wire _6139_ ;
wire _1694_ ;
wire _1274_ ;
wire _1985__bF$buf0 ;
wire _1985__bF$buf1 ;
wire _1985__bF$buf2 ;
wire _1985__bF$buf3 ;
wire _1985__bF$buf4 ;
wire _1985__bF$buf5 ;
wire _185_ ;
wire _2899_ ;
wire _2479_ ;
wire _2059_ ;
wire _3840_ ;
wire _3420_ ;
wire _3000_ ;
wire selXY ;
wire _4625_ ;
wire _4205_ ;
wire _5583_ ;
wire _5163_ ;
wire _1083_ ;
wire _2288_ ;
wire _4854_ ;
wire _4434_ ;
wire _4014_ ;
wire _5639_ ;
wire _5219_ ;
wire _1979_ ;
wire _1559_ ;
wire _1139_ ;
wire _2920_ ;
wire _2500_ ;
wire _5392_ ;
wire _3705_ ;
wire _6177_ ;
wire _2097_ ;
wire _4663_ ;
wire _4243_ ;
wire _5868_ ;
wire _5448_ ;
wire _5028_ ;
wire _1788_ ;
wire _1368_ ;
wire \genblk1[1].u_ce.Vld_bF$buf0  ;
wire _699_ ;
wire _279_ ;
wire _3934_ ;
wire _3514_ ;
wire _4719_ ;
wire _4892_ ;
wire _4472_ ;
wire _4052_ ;
wire [6:0] \genblk1[0].u_ce.ISpipe  ;
wire _911_ ;
wire _5677_ ;
wire _5257_ ;
wire _1597_ ;
wire _1177_ ;
wire _3743_ ;
wire _3323_ ;
wire _4948_ ;
wire _4528_ ;
wire _4108_ ;
wire _4281_ ;
wire _720_ ;
wire _300_ ;
wire _5486_ ;
wire _5066_ ;
wire _3972_ ;
wire _3552_ ;
wire _3132_ ;
wire _4757_ ;
wire _4337_ ;
wire _36_ ;
wire _4090_ ;
wire _2823_ ;
wire _2403_ ;
wire _5295_ ;
wire _3608_ ;
wire _3781_ ;
wire _3361_ ;
wire _4986_ ;
wire _4566_ ;
wire _4146_ ;
wire _2632_ ;
wire _2212_ ;
wire _3837_ ;
wire _3417_ ;
wire _3590_ ;
wire _3170_ ;
wire _1903_ ;
wire _4795_ ;
wire _4375_ ;
wire _814_ ;
wire [6:0] \genblk1[2].u_ce.ISpipe  ;
wire _74_ ;
wire _6101_ ;
wire _2861_ ;
wire _2441_ ;
wire _2021_ ;
wire _3646_ ;
wire _3226_ ;
wire _1712_ ;
wire _4184_ ;
wire _623_ ;
wire _203_ ;
wire _2917_ ;
wire _5389_ ;
wire _6330_ ;
wire _2670_ ;
wire _2250_ ;
wire _3875_ ;
wire _3455_ ;
wire _3035_ ;
wire \genblk1[3].u_ce.Ain12b_11_bF$buf2  ;
wire _5601_ ;
wire [1:0] \genblk1[4].u_ce.Ain1  ;
wire _1941_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _2726_ ;
wire _2306_ ;
wire _5198_ ;
wire _3684_ ;
wire _3264_ ;
wire _4889_ ;
wire _4469_ ;
wire _4049_ ;
wire _5830_ ;
wire _5410_ ;
wire _908_ ;
wire _1750_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire [11:0] \genblk1[4].u_ce.Ycalc  ;
wire _2955_ ;
wire _2535_ ;
wire _2115_ ;
wire \genblk1[0].u_ce.LoadCtl_0_bF$buf3  ;
wire _3493_ ;
wire _3073_ ;
wire _1806_ ;
wire _4698_ ;
wire _4278_ ;
wire _717_ ;
wire _6004_ ;
wire [6:0] \genblk1[4].u_ce.ISpipe  ;
wire _890_ ;
wire _470_ ;
wire _2764_ ;
wire _2344_ ;
wire _3969_ ;
wire _3549_ ;
wire _3129_ ;
wire _4910_ ;
wire _1615_ ;
wire _4087_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _6233_ ;
wire _2993_ ;
wire _2573_ ;
wire _2153_ ;
wire _3778_ ;
wire _3358_ ;
wire _5924_ ;
wire _5504_ ;
wire _1844_ ;
wire [1:0] \genblk1[5].u_ce.Xin0  ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire _2629_ ;
wire _2209_ ;
wire _6042_ ;
wire _2382_ ;
wire _3587_ ;
wire _3167_ ;
wire _5733_ ;
wire _5313_ ;
wire _1653_ ;
wire _1233_ ;
wire [11:0] \genblk1[5].u_ce.Acalc  ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _2858_ ;
wire _2438_ ;
wire _2018_ ;
wire _6271_ ;
wire _2191_ ;
wire _3396_ ;
wire _1709_ ;
wire _5962_ ;
wire _5542_ ;
wire _5122_ ;
wire _6327_ ;
wire _1882_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire [6:0] \genblk1[6].u_ce.ISpipe  ;
wire _2667_ ;
wire _2247_ ;
wire _6080_ ;
wire _4813_ ;
wire _1938_ ;
wire _1518_ ;
wire _5771_ ;
wire _5351_ ;
wire _849_ ;
wire _429_ ;
wire _6136_ ;
wire _1691_ ;
wire _1271_ ;
wire _182_ ;
wire _2896_ ;
wire _2476_ ;
wire _2056_ ;
wire _4622_ ;
wire _4202_ ;
wire _5827_ ;
wire _5407_ ;
wire _1747_ ;
wire _1327_ ;
wire _5580_ ;
wire _5160_ ;
wire _658_ ;
wire _238_ ;
wire _1080_ ;
wire _2285_ ;
wire _4851_ ;
wire _4431_ ;
wire _4011_ ;
wire _5636_ ;
wire _5216_ ;
wire _1976_ ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _3702_ ;
wire _6174_ ;
wire _4907_ ;
wire _2094_ ;
wire _3299_ ;
wire _4660_ ;
wire _4240_ ;
wire _5865_ ;
wire _5445_ ;
wire _5025_ ;
wire _1785_ ;
wire _1365_ ;
wire _696_ ;
wire _276_ ;
wire _3931_ ;
wire _3511_ ;
wire _4716_ ;
wire \genblk1[0].u_ce.Vld  ;
wire _5674_ ;
wire _5254_ ;
wire _6039_ ;
wire _1594_ ;
wire _1174_ ;
wire _2799_ ;
wire _2379_ ;
wire _3740_ ;
wire _3320_ ;
wire _4945_ ;
wire _4525_ ;
wire _4105_ ;
wire _5483_ ;
wire _5063_ ;
wire _6268_ ;
wire _2188_ ;
wire _4754_ ;
wire _4334_ ;
wire _5959_ ;
wire _5539_ ;
wire _5119_ ;
wire _33_ ;
wire _1879_ ;
wire _1459_ ;
wire _1039_ ;
wire _2820_ ;
wire _2400_ ;
wire _5292_ ;
wire _3605_ ;
wire _6077_ ;
wire _4983_ ;
wire _4563_ ;
wire _4143_ ;
wire _5768_ ;
wire _5348_ ;
wire _1688_ ;
wire _1268_ ;
wire _599_ ;
wire _179_ ;
wire _3834_ ;
wire _3414_ ;
wire _4619_ ;
wire _1900_ ;
wire _4792_ ;
wire _4372_ ;
wire _811_ ;
wire _5997_ ;
wire _5577_ ;
wire _5157_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _4507__bF$buf0 ;
wire _4507__bF$buf1 ;
wire _4507__bF$buf2 ;
wire _4507__bF$buf3 ;
wire _3643_ ;
wire _3223_ ;
wire [1:0] \u_ot.Yin1  ;
wire _4848_ ;
wire _4428_ ;
wire _4008_ ;
wire _4181_ ;
wire _620_ ;
wire _200_ ;
wire _2914_ ;
wire _5386_ ;
wire _3872_ ;
wire _3452_ ;
wire _3032_ ;
wire _4657_ ;
wire _4237_ ;
wire _2723_ ;
wire _2303_ ;
wire _5195_ ;
wire _3928_ ;
wire _3508_ ;
wire _3681_ ;
wire _3261_ ;
wire _4886_ ;
wire _4466_ ;
wire _4046_ ;
wire _905_ ;
wire _2952_ ;
wire _2532_ ;
wire _2112_ ;
wire _3737_ ;
wire _3317_ ;
wire \genblk1[0].u_ce.LoadCtl_0_bF$buf0  ;
wire _3490_ ;
wire _3070_ ;
wire _1803_ ;
wire _4695_ ;
wire _4275_ ;
wire _714_ ;
wire _6001_ ;
wire _2761_ ;
wire _2341_ ;
wire _3966_ ;
wire _3546_ ;
wire _3126_ ;
wire [1:0] \genblk1[5].u_ce.Y_  ;
wire _1612_ ;
wire _4084_ ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _2817_ ;
wire _5289_ ;
wire _6230_ ;
wire _2990_ ;
wire _2570_ ;
wire _2150_ ;
wire _3775_ ;
wire _3355_ ;
wire _5921_ ;
wire _5501_ ;
wire _1841_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire _2626_ ;
wire _2206_ ;
wire _5098_ ;
wire _3584_ ;
wire _3164_ ;
wire _4789_ ;
wire _4369_ ;
wire _5730_ ;
wire _5310_ ;
wire _808_ ;
wire _68_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _2855_ ;
wire _2435_ ;
wire _2015_ ;
wire _3393_ ;
wire _1706_ ;
wire _4598_ ;
wire _4178_ ;
wire _617_ ;
wire _6324_ ;
wire _790_ ;
wire _370_ ;
wire _2664_ ;
wire _2244_ ;
wire [11:0] \genblk1[1].u_ce.Yin12b  ;
wire _3869_ ;
wire _3449_ ;
wire _3029_ ;
wire _4810_ ;
wire _1935_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _6133_ ;
wire _2893_ ;
wire _2473_ ;
wire _2053_ ;
wire _3678_ ;
wire _3258_ ;
wire _5824_ ;
wire _5404_ ;
wire _1744_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _2949_ ;
wire _2529_ ;
wire _2109_ ;
wire _2282_ ;
wire _3487_ ;
wire _3067_ ;
wire _5633_ ;
wire _5213_ ;
wire _1973_ ;
wire _1553_ ;
wire _1133_ ;
wire \genblk1[5].u_ce.LoadCtl_0_bF$buf3  ;
wire _884_ ;
wire _464_ ;
wire _2758_ ;
wire _2338_ ;
wire \genblk1[4].u_ce.Vld_bF$buf2  ;
wire _6171_ ;
wire _4904_ ;
wire _2091_ ;
wire _3296_ ;
wire _1609_ ;
wire _5862_ ;
wire _5442_ ;
wire _5022_ ;
wire _6227_ ;
wire _1782_ ;
wire _1362_ ;
wire _693_ ;
wire _273_ ;
wire _2987_ ;
wire _2567_ ;
wire _2147_ ;
wire \genblk1[3].u_ce.ISout  ;
wire _4713_ ;
wire _5918_ ;
wire _1838_ ;
wire _1418_ ;
wire _5671_ ;
wire _5251_ ;
wire _749_ ;
wire _329_ ;
wire _6036_ ;
wire _1591_ ;
wire _1171_ ;
wire _2796_ ;
wire _2376_ ;
wire _4942_ ;
wire _4522_ ;
wire _4102_ ;
wire _5727_ ;
wire _5307_ ;
wire _1647_ ;
wire _1227_ ;
wire _5480_ ;
wire _5060_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _6265_ ;
wire _2185_ ;
wire [11:0] \genblk1[6].u_ce.Xcalc  ;
wire _4751_ ;
wire _4331_ ;
wire _5956_ ;
wire _5536_ ;
wire _5116_ ;
wire _30_ ;
wire En ;
wire _1876_ ;
wire _1456_ ;
wire _1036_ ;
wire _787_ ;
wire _367_ ;
wire _3602_ ;
wire _6074_ ;
wire _4807_ ;
wire _3199_ ;
wire _4980_ ;
wire _4560_ ;
wire _4140_ ;
wire _5765_ ;
wire _5345_ ;
wire \genblk1[1].u_ce.Ain12b_11_bF$buf2  ;
wire _1685_ ;
wire _1265_ ;
wire _596_ ;
wire _176_ ;
wire _3831_ ;
wire _3411_ ;
wire _4616_ ;
wire _5994_ ;
wire _5574_ ;
wire _5154_ ;
wire _1494_ ;
wire _1074_ ;
wire [1:0] \a[2]  ;
wire _2699_ ;
wire _2279_ ;
wire _3640_ ;
wire _3220_ ;
wire _4845_ ;
wire _4425_ ;
wire _4005_ ;
wire _2911_ ;
wire \genblk1[5].u_ce.Vld  ;
wire _5383_ ;
wire _6168_ ;
wire clk_hier0_bF$buf0 ;
wire clk_hier0_bF$buf1 ;
wire clk_hier0_bF$buf2 ;
wire clk_hier0_bF$buf3 ;
wire clk_hier0_bF$buf4 ;
wire clk_hier0_bF$buf5 ;
wire clk_hier0_bF$buf6 ;
wire clk_hier0_bF$buf7 ;
wire _2088_ ;
wire [1:0] \genblk1[0].u_ce.Yin1  ;
wire _4654_ ;
wire _4234_ ;
wire _5859_ ;
wire _5439_ ;
wire _5019_ ;
wire [1:0] \genblk1[3].u_ce.Ain0  ;
wire _1779_ ;
wire _1359_ ;
wire _2720_ ;
wire _2300_ ;
wire _5192_ ;
wire _3925_ ;
wire _3505_ ;
wire _4883_ ;
wire _4463_ ;
wire _4043_ ;
wire _902_ ;
wire _5668_ ;
wire _5248_ ;
wire _1588_ ;
wire _1168_ ;
wire [1:0] \genblk1[0].u_ce.X_  ;
wire _499_ ;
wire _3734_ ;
wire _3314_ ;
wire _4939_ ;
wire _4519_ ;
wire \genblk1[6].u_ce.Ain12b_11_bF$buf3  ;
wire _1800_ ;
wire _4692_ ;
wire _4272_ ;
wire _711_ ;
wire _5897_ ;
wire _5477_ ;
wire _5057_ ;
wire _1397_ ;
wire _3963_ ;
wire _3543_ ;
wire _3123_ ;
wire _4748_ ;
wire _4328_ ;
wire _27_ ;
wire _4081_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire _2814_ ;
wire _5286_ ;
wire \genblk1[3].u_ce.LoadCtl_0_bF$buf4  ;
wire _3772_ ;
wire _3352_ ;
wire _4977_ ;
wire _4557_ ;
wire _4137_ ;
wire _2623_ ;
wire _2203_ ;
wire _5095_ ;
wire _3828_ ;
wire _3408_ ;
wire _3581_ ;
wire _3161_ ;
wire _4786_ ;
wire _4366_ ;
wire _805_ ;
wire _65_ ;
wire _2852_ ;
wire _2432_ ;
wire _2012_ ;
wire _3637_ ;
wire _3217_ ;
wire _3390_ ;
wire _1703_ ;
wire _4595_ ;
wire _4175_ ;
wire _614_ ;
wire _2908_ ;
wire _6321_ ;
wire _2661_ ;
wire _2241_ ;
wire _3866_ ;
wire _3446_ ;
wire _3026_ ;
wire _1932_ ;
wire _1512_ ;
wire _843_ ;
wire _423_ ;
wire _2717_ ;
wire _5189_ ;
wire _6130_ ;
wire _2890_ ;
wire _2470_ ;
wire _2050_ ;
wire _3675_ ;
wire _3255_ ;
wire _5821_ ;
wire _5401_ ;
wire _1741_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _2946_ ;
wire _2526_ ;
wire _2106_ ;
wire _3484_ ;
wire _3064_ ;
wire _4689_ ;
wire _4269_ ;
wire _5630_ ;
wire _5210_ ;
wire _708_ ;
wire _1970_ ;
wire _1550_ ;
wire _1130_ ;
wire \genblk1[5].u_ce.LoadCtl_0_bF$buf0  ;
wire _881_ ;
wire _461_ ;
wire _2755_ ;
wire _2335_ ;
wire _4901_ ;
wire _3293_ ;
wire _1606_ ;
wire _4498_ ;
wire _4078_ ;
wire _937_ ;
wire _517_ ;
wire _6224_ ;
wire [6:0] \genblk1[3].u_ce.LoadCtl  ;
wire _690_ ;
wire _270_ ;
wire _2984_ ;
wire _2564_ ;
wire _2144_ ;
wire _3769_ ;
wire _3349_ ;
wire _4710_ ;
wire _5915_ ;
wire _1835_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _6033_ ;
wire _2793_ ;
wire _2373_ ;
wire _3998_ ;
wire _3578_ ;
wire _3158_ ;
wire _5724_ ;
wire _5304_ ;
wire _1644_ ;
wire _1224_ ;
wire [1:0] \genblk1[6].u_ce.Yin0  ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire _2849_ ;
wire _2429_ ;
wire _2009_ ;
wire _6262_ ;
wire _2182_ ;
wire _3387_ ;
wire _5953_ ;
wire _5533_ ;
wire _5113_ ;
wire _6318_ ;
wire _1873_ ;
wire _1453_ ;
wire _1033_ ;
wire [11:0] \genblk1[1].u_ce.Ycalc  ;
wire _784_ ;
wire _364_ ;
wire _2658_ ;
wire _2238_ ;
wire _6071_ ;
wire _4804_ ;
wire _3196_ ;
wire _1929_ ;
wire _1509_ ;
wire _5762_ ;
wire _5342_ ;
wire _6127_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _2887_ ;
wire _2467_ ;
wire _2047_ ;
wire _4613_ ;
wire _5818_ ;
wire _1738_ ;
wire _1318_ ;
wire _5991_ ;
wire _5571_ ;
wire _5151_ ;
wire _649_ ;
wire _229_ ;
wire _1491_ ;
wire _1071_ ;
wire _2696_ ;
wire _2276_ ;
wire _4842_ ;
wire _4422_ ;
wire _4002_ ;
wire _5627_ ;
wire _5207_ ;
wire _1967_ ;
wire _1547_ ;
wire _1127_ ;
wire _5380_ ;
wire _878_ ;
wire _458_ ;
wire _6165_ ;
wire _2085_ ;
wire _4651_ ;
wire _4231_ ;
wire _5856_ ;
wire _5436_ ;
wire _5016_ ;
wire _1776_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _3922_ ;
wire _3502_ ;
wire _4707_ ;
wire _3099_ ;
wire _4880_ ;
wire _4460_ ;
wire _4040_ ;
wire _5665_ ;
wire _5245_ ;
wire _1585_ ;
wire _1165_ ;
wire _496_ ;
wire _3731_ ;
wire _3311_ ;
wire _4936_ ;
wire _4516_ ;
wire \genblk1[6].u_ce.Ain12b_11_bF$buf0  ;
wire _5894_ ;
wire _5474_ ;
wire _5054_ ;
wire _6259_ ;
wire _1394_ ;
wire _2599_ ;
wire _2179_ ;
wire _3960_ ;
wire _3540_ ;
wire _3120_ ;
wire _4745_ ;
wire _4325_ ;
wire _24_ ;
wire _1119__bF$buf0 ;
wire _1119__bF$buf1 ;
wire _1119__bF$buf2 ;
wire _1119__bF$buf3 ;
wire _1119__bF$buf4 ;
wire _1119__bF$buf5 ;
wire _2811_ ;
wire _5283_ ;
wire _6068_ ;
wire \genblk1[3].u_ce.LoadCtl_0_bF$buf1  ;
wire _4974_ ;
wire _4554_ ;
wire _4134_ ;
wire _5759_ ;
wire _5339_ ;
wire _1679_ ;
wire _1259_ ;
wire [1:0] \genblk1[3].u_ce.Xin1  ;
wire _2620_ ;
wire _2200_ ;
wire _5092_ ;
wire _3825_ ;
wire _3405_ ;
wire _6297_ ;
wire _4783_ ;
wire _4363_ ;
wire _802_ ;
wire _5988_ ;
wire _5568_ ;
wire _5148_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _399_ ;
wire _3634_ ;
wire _3214_ ;
wire _4839_ ;
wire _4419_ ;
wire _1700_ ;
wire _4592_ ;
wire _4172_ ;
wire _611_ ;
wire _2905_ ;
wire _5797_ ;
wire _5377_ ;
wire _1297_ ;
wire _3863_ ;
wire _3443_ ;
wire _3023_ ;
wire _4648_ ;
wire _4228_ ;
wire _840_ ;
wire _420_ ;
wire _2714_ ;
wire _5186_ ;
wire _3919_ ;
wire _3672_ ;
wire _3252_ ;
wire _4877_ ;
wire _4457_ ;
wire _4037_ ;
wire _2943_ ;
wire _2523_ ;
wire _2103_ ;
wire _3728_ ;
wire _3308_ ;
wire _3481_ ;
wire _3061_ ;
wire _4686_ ;
wire _4266_ ;
wire _705_ ;
wire _2752_ ;
wire _2332_ ;
wire _3957_ ;
wire _3537_ ;
wire _3117_ ;
wire \genblk1[2].u_ce.Vld_bF$buf2  ;
wire _3290_ ;
wire _1603_ ;
wire _4495_ ;
wire _4075_ ;
wire [11:0] \genblk1[6].u_ce.Ain12b  ;
wire _934_ ;
wire _514_ ;
wire _2808_ ;
wire _6221_ ;
wire [1:0] \genblk1[6].u_ce.Y_  ;
wire _2981_ ;
wire _2561_ ;
wire _2141_ ;
wire _3766_ ;
wire _3346_ ;
wire _5912_ ;
wire _1832_ ;
wire _1412_ ;
wire _743_ ;
wire _323_ ;
wire _2617_ ;
wire _5089_ ;
wire _6030_ ;
wire _2790_ ;
wire _2370_ ;
wire _3995_ ;
wire _3575_ ;
wire _3155_ ;
wire _5721_ ;
wire _5301_ ;
wire _59_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _2846_ ;
wire _2426_ ;
wire _2006_ ;
wire _3384_ ;
wire _4589_ ;
wire _4169_ ;
wire _5950_ ;
wire _5530_ ;
wire _5110_ ;
wire _608_ ;
wire _6315_ ;
wire _1870_ ;
wire _1450_ ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _2655_ ;
wire _2235_ ;
wire _4801_ ;
wire _3193_ ;
wire _1926_ ;
wire _1506_ ;
wire _4398_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _6124_ ;
wire _590_ ;
wire _170_ ;
wire _2884_ ;
wire _2464_ ;
wire _2044_ ;
wire _3669_ ;
wire _3249_ ;
wire _4610_ ;
wire _5815_ ;
wire _1735_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire _2693_ ;
wire _2273_ ;
wire _3898_ ;
wire _3478_ ;
wire _3058_ ;
wire _5624_ ;
wire _5204_ ;
wire _1964_ ;
wire _1544_ ;
wire \genblk1[4].u_ce.Ain12b_11_bF$buf3  ;
wire _1124_ ;
wire _875_ ;
wire _455_ ;
wire _2749_ ;
wire _2329_ ;
wire _6162_ ;
wire _2082_ ;
wire _3287_ ;
wire _5853_ ;
wire _5433_ ;
wire _5013_ ;
wire _6218_ ;
wire _1773_ ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _2978_ ;
wire _2558_ ;
wire _2138_ ;
wire _4704_ ;
wire [11:0] Dout ;
wire _5909_ ;
wire _3096_ ;
wire \genblk1[1].u_ce.LoadCtl_0_bF$buf4  ;
wire _1829_ ;
wire _1409_ ;
wire _5662_ ;
wire _5242_ ;
wire _6027_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _2787_ ;
wire _2367_ ;
wire _4933_ ;
wire _4513_ ;
wire _5718_ ;
wire _1638_ ;
wire _1218_ ;
wire _5891_ ;
wire _5471_ ;
wire _5051_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _6256_ ;
wire _1391_ ;
wire _2596_ ;
wire _2176_ ;
wire _4742_ ;
wire _4322_ ;
wire _5947_ ;
wire _5527_ ;
wire _5107_ ;
wire _21_ ;
wire _1867_ ;
wire _1447_ ;
wire _1027_ ;
wire _5280_ ;
wire _778_ ;
wire _358_ ;
wire _6065_ ;
wire _4971_ ;
wire _4551_ ;
wire _4131_ ;
wire _5756_ ;
wire _5336_ ;
wire _1676_ ;
wire _1256_ ;
wire _587_ ;
wire _167_ ;
wire _3822_ ;
wire _3402_ ;
wire _6294_ ;
wire _4607_ ;
wire _4780_ ;
wire _4360_ ;
wire _5985_ ;
wire _5565_ ;
wire _5145_ ;
wire _1485_ ;
wire _1065_ ;
wire \genblk1[0].u_ce.ISout  ;
wire _396_ ;
wire _3631_ ;
wire _3211_ ;
wire _4836_ ;
wire _4416_ ;
wire _2902_ ;
wire _5794_ ;
wire _5374_ ;
wire _6159_ ;
wire _1294_ ;
wire _2499_ ;
wire _2079_ ;
wire _3860_ ;
wire _3440_ ;
wire _3020_ ;
wire _4645_ ;
wire _4225_ ;
wire \genblk1[0].u_ce.Vld_bF$buf3  ;
wire _2711_ ;
wire _5183_ ;
wire _3916_ ;
wire [11:0] \genblk1[3].u_ce.Xcalc  ;
wire _4874_ ;
wire _4454_ ;
wire _4034_ ;
wire _5659_ ;
wire _5239_ ;
wire _1999_ ;
wire _1579_ ;
wire _1159_ ;
wire _2940_ ;
wire _2520_ ;
wire _2100_ ;
wire _3725_ ;
wire _3305_ ;
wire _6197_ ;
wire _4683_ ;
wire _4263_ ;
wire _702_ ;
wire [1:0] \genblk1[1].u_ce.X_  ;
wire _5888_ ;
wire _5468_ ;
wire _5048_ ;
wire _1388_ ;
wire _299_ ;
wire _3954_ ;
wire _3534_ ;
wire _3114_ ;
wire [6:0] \genblk1[1].u_ce.ISpipe  ;
wire _4739_ ;
wire _4319_ ;
wire _1890__bF$buf0 ;
wire _1890__bF$buf1 ;
wire _1890__bF$buf2 ;
wire _1890__bF$buf3 ;
wire _1890__bF$buf4 ;
wire _18_ ;
wire _1600_ ;
wire _4492_ ;
wire _4072_ ;
wire _931_ ;
wire _511_ ;
wire _2805_ ;
wire _5697_ ;
wire _5277_ ;
wire _1197_ ;
wire _3763_ ;
wire _3343_ ;
wire _4968_ ;
wire _4548_ ;
wire _4128_ ;
wire _740_ ;
wire _320_ ;
wire _2614_ ;
wire _5086_ ;
wire _3819_ ;
wire _3992_ ;
wire _3572_ ;
wire _3152_ ;
wire _4777_ ;
wire _4357_ ;
wire _56_ ;
wire _2843_ ;
wire _2423_ ;
wire _2003_ ;
wire _3628_ ;
wire _3208_ ;
wire _3381_ ;
wire _4586_ ;
wire _4166_ ;
wire _605_ ;
wire _6312_ ;
wire _2652_ ;
wire _2232_ ;
wire \u_ot.ISout_bF$buf4  ;
wire _3857_ ;
wire _3437_ ;
wire _3017_ ;
wire [6:0] \genblk1[3].u_ce.ISpipe  ;
wire _3190_ ;
wire _1923_ ;
wire _1503_ ;
wire _4395_ ;
wire _834_ ;
wire _414_ ;
wire _2708_ ;
wire _94_ ;
wire _6121_ ;
wire _2881_ ;
wire _2461_ ;
wire _2041_ ;
wire _3666_ ;
wire _3246_ ;
wire _5812_ ;
wire _1732_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _2937_ ;
wire _2517_ ;
wire _2690_ ;
wire _2270_ ;
wire _3895_ ;
wire _3475_ ;
wire _3055_ ;
wire _5621_ ;
wire _5201_ ;
wire _1961_ ;
wire _1541_ ;
wire \genblk1[4].u_ce.Ain12b_11_bF$buf0  ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _2746_ ;
wire _2326_ ;
wire _3284_ ;
wire _4489_ ;
wire _4069_ ;
wire _5850_ ;
wire _5430_ ;
wire _5010_ ;
wire _928_ ;
wire _508_ ;
wire _6215_ ;
wire [1:0] \genblk1[1].u_ce.Ain1  ;
wire _1770_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _2975_ ;
wire _2555_ ;
wire _2135_ ;
wire _4701_ ;
wire _5906_ ;
wire _3093_ ;
wire \genblk1[1].u_ce.LoadCtl_0_bF$buf1  ;
wire _1826_ ;
wire _1406_ ;
wire _4298_ ;
wire _737_ ;
wire _317_ ;
wire _6024_ ;
wire _490_ ;
wire _2784_ ;
wire _2364_ ;
wire _3989_ ;
wire _3569_ ;
wire _3149_ ;
wire _4930_ ;
wire _4510_ ;
wire _5715_ ;
wire _1635_ ;
wire _1215_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _6253_ ;
wire _2593_ ;
wire _2173_ ;
wire _3798_ ;
wire _3378_ ;
wire _5944_ ;
wire _5524_ ;
wire _5104_ ;
wire _6309_ ;
wire _1864_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _2649_ ;
wire _2229_ ;
wire _6062_ ;
wire _3187_ ;
wire _5753_ ;
wire _5333_ ;
wire _6118_ ;
wire _1673_ ;
wire _1253_ ;
wire [1:0] \genblk1[2].u_ce.Xin0  ;
wire _584_ ;
wire _164_ ;
wire _2878_ ;
wire _2458_ ;
wire _2038_ ;
wire _6291_ ;
wire _4604_ ;
wire _5809_ ;
wire _5270__bF$buf0 ;
wire _5270__bF$buf1 ;
wire _5270__bF$buf2 ;
wire _5270__bF$buf3 ;
wire _1729_ ;
wire _1309_ ;
wire _5982_ ;
wire _5562_ ;
wire _5142_ ;
wire _6347_ ;
wire _1482_ ;
wire _1062_ ;
wire _393_ ;
wire _2687_ ;
wire _2267_ ;
wire _4833_ ;
wire _4413_ ;
wire _5618_ ;
wire _1958_ ;
wire _1538_ ;
wire _1118_ ;
wire _5791_ ;
wire _5371_ ;
wire _869_ ;
wire _449_ ;
wire _6156_ ;
wire _1291_ ;
wire _2496_ ;
wire _2076_ ;
wire _4642_ ;
wire _4222_ ;
wire _5847_ ;
wire _5427_ ;
wire _5007_ ;
wire \genblk1[0].u_ce.Vld_bF$buf0  ;
wire _1767_ ;
wire _1347_ ;
wire _5180_ ;
wire _678_ ;
wire _258_ ;
wire _3913_ ;
wire _4871_ ;
wire _4451_ ;
wire _4031_ ;
wire _5656_ ;
wire _5236_ ;
wire _1996_ ;
wire _1576_ ;
wire _1156_ ;
wire _487_ ;
wire _3722_ ;
wire _3302_ ;
wire _6194_ ;
wire _4927_ ;
wire _4507_ ;
wire _4680_ ;
wire _4260_ ;
wire _5885_ ;
wire _5465_ ;
wire _5045_ ;
wire _1385_ ;
wire _296_ ;
wire _3951_ ;
wire _3531_ ;
wire _3111_ ;
wire _4736_ ;
wire _4316_ ;
wire _15_ ;
wire _2802_ ;
wire _5694_ ;
wire _5274_ ;
wire _6059_ ;
wire _1194_ ;
wire _2399_ ;
wire _3760_ ;
wire _3340_ ;
wire _4965_ ;
wire _4545_ ;
wire _4125_ ;
wire _2611_ ;
wire _5083_ ;
wire _3816_ ;
wire _6288_ ;
wire _4774_ ;
wire _4354_ ;
wire _5979_ ;
wire _5559_ ;
wire _5139_ ;
wire _53_ ;
wire _1899_ ;
wire _1479_ ;
wire _1059_ ;
wire _2840_ ;
wire _2420_ ;
wire _2000_ ;
wire [1:0] \genblk1[4].u_ce.Yin1  ;
wire _3625_ ;
wire _3205_ ;
wire _6097_ ;
wire _4583_ ;
wire _4163_ ;
wire _602_ ;
wire \genblk1[3].u_ce.Vld  ;
wire _5788_ ;
wire _5368_ ;
wire _1288_ ;
wire _199_ ;
wire \u_ot.ISout_bF$buf1  ;
wire \genblk1[2].u_ce.Ain12b_11_bF$buf3  ;
wire _3854_ ;
wire _3434_ ;
wire _3014_ ;
wire _4639_ ;
wire _4219_ ;
wire _1920_ ;
wire _1500_ ;
wire _4392_ ;
wire _831_ ;
wire _411_ ;
wire _2705_ ;
wire _5597_ ;
wire _5177_ ;
wire _91_ ;
wire _1097_ ;
wire _3663_ ;
wire _3243_ ;
wire _4868_ ;
wire _4448_ ;
wire _4028_ ;
wire _640_ ;
wire _220_ ;
wire _2934_ ;
wire _2514_ ;
wire _3719_ ;
wire _2762__bF$buf0 ;
wire _2762__bF$buf1 ;
wire _2762__bF$buf2 ;
wire _2762__bF$buf3 ;
wire _2762__bF$buf4 ;
wire _3892_ ;
wire _3472_ ;
wire _3052_ ;
wire _4677_ ;
wire _4257_ ;
wire _2743_ ;
wire _2323_ ;
wire _3948_ ;
wire _3528_ ;
wire _3108_ ;
wire _9_ ;
wire _3281_ ;
wire _4486_ ;
wire _4066_ ;
wire _925_ ;
wire _505_ ;
wire _6212_ ;
wire _2972_ ;
wire _2552_ ;
wire _2132_ ;
wire _3757_ ;
wire _3337_ ;
wire _5903_ ;
wire _3090_ ;
wire _1823_ ;
wire _1403_ ;
wire _4295_ ;
wire _734_ ;
wire _314_ ;
wire _2608_ ;
wire _6021_ ;
wire _2781_ ;
wire _2361_ ;
wire _3986_ ;
wire _3566_ ;
wire _3146_ ;
wire _5712_ ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _2837_ ;
wire _2417_ ;
wire _6250_ ;
wire _2590_ ;
wire _2170_ ;
wire _3795_ ;
wire _3375_ ;
wire _5941_ ;
wire _5521_ ;
wire _5101_ ;
wire _6306_ ;
wire _1861_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _2646_ ;
wire _2226_ ;
wire _3184_ ;
wire _1917_ ;
wire _4389_ ;
wire _5750_ ;
wire _5330_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _6115_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _2875_ ;
wire _2455_ ;
wire _2035_ ;
wire _4601_ ;
wire _5806_ ;
wire _1726_ ;
wire _1306_ ;
wire _4198_ ;
wire _637_ ;
wire _217_ ;
wire _6344_ ;
wire _390_ ;
wire _2684_ ;
wire _2264_ ;
wire _3889_ ;
wire _3469_ ;
wire _3049_ ;
wire _4830_ ;
wire _4410_ ;
wire _5615_ ;
wire _1955_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire _6153_ ;
wire _2493_ ;
wire _2073_ ;
wire _3698_ ;
wire _3278_ ;
wire [11:0] \genblk1[5].u_ce.Ycalc  ;
wire _5844_ ;
wire _5424_ ;
wire _5004_ ;
wire _6209_ ;
wire _1764_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _2969_ ;
wire _2549_ ;
wire _2129_ ;
wire _3910_ ;
wire _3087_ ;
wire _5653_ ;
wire _5233_ ;
wire _6018_ ;
wire _1993_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _2778_ ;
wire _2358_ ;
wire _6191_ ;
wire \genblk1[6].u_ce.LoadCtl_0_bF$buf1  ;
wire _4924_ ;
wire _4504_ ;
wire \genblk1[5].u_ce.Vld_bF$buf1  ;
wire _5709_ ;
wire _1629_ ;
wire _1209_ ;
wire _5882_ ;
wire _5462_ ;
wire _5042_ ;
wire _6247_ ;
wire _1382_ ;
wire _293_ ;
wire _2587_ ;
wire _2167_ ;
wire _4733_ ;
wire _4313_ ;
wire _5938_ ;
wire _5518_ ;
wire _12_ ;
wire _1858_ ;
wire _1438_ ;
wire _1018_ ;
wire _5691_ ;
wire _5271_ ;
wire _769_ ;
wire _349_ ;
wire _6056_ ;
wire _1191_ ;
wire _2396_ ;
wire _4962_ ;
wire _4542_ ;
wire _4122_ ;
wire _5747_ ;
wire _5327_ ;
wire _1667_ ;
wire _1247_ ;
wire _5080_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _3813_ ;
wire _6285_ ;
wire _4771_ ;
wire _4351_ ;
wire _5976_ ;
wire _5556_ ;
wire _5136_ ;
wire _50_ ;
wire _1896_ ;
wire _1476_ ;
wire _1056_ ;
wire _387_ ;
wire _3622_ ;
wire _3202_ ;
wire _6094_ ;
wire _4827_ ;
wire _4407_ ;
wire [6:0] \genblk1[0].u_ce.LoadCtl  ;
wire _4580_ ;
wire _4160_ ;
wire _5785_ ;
wire _5365_ ;
wire _1285_ ;
wire _196_ ;
wire \genblk1[2].u_ce.Ain12b_11_bF$buf0  ;
wire _3851_ ;
wire _3431_ ;
wire _3011_ ;
wire _4636_ ;
wire _4216_ ;
wire _2702_ ;
wire _5594_ ;
wire _5174_ ;
wire _3907_ ;
wire _1094_ ;
wire [1:0] \a[4]  ;
wire _2299_ ;
wire _3660_ ;
wire _3240_ ;
wire _4865_ ;
wire _4445_ ;
wire _4025_ ;
wire _2931_ ;
wire _2511_ ;
wire _3716_ ;
wire _6188_ ;
wire [19:0] \u_pa.acc_reg  ;
wire _4674_ ;
wire _4254_ ;
wire _5879_ ;
wire _5459_ ;
wire _5039_ ;
wire _1799_ ;
wire _1379_ ;
wire _2740_ ;
wire _2320_ ;
wire _3945_ ;
wire _3525_ ;
wire _3105_ ;
wire _6_ ;
wire [1:0] \genblk1[2].u_ce.X_  ;
wire _4483_ ;
wire _4063_ ;
wire _922_ ;
wire _502_ ;
wire _5688_ ;
wire _5268_ ;
wire [1:0] \genblk1[0].u_ce.Ain0  ;
wire _1188_ ;
wire _3754_ ;
wire _3334_ ;
wire _4959_ ;
wire _4539_ ;
wire _4119_ ;
wire _5900_ ;
wire _1820_ ;
wire _1400_ ;
wire _4292_ ;
wire _731_ ;
wire _311_ ;
wire _2605_ ;
wire _5497_ ;
wire _5077_ ;
wire [6:0] \genblk1[5].u_ce.LoadCtl  ;
wire _3983_ ;
wire _3563_ ;
wire _3143_ ;
wire _4768_ ;
wire _4348_ ;
wire _47_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _2834_ ;
wire _2414_ ;
wire _3619_ ;
wire [11:0] \genblk1[0].u_ce.Xcalc  ;
wire _3792_ ;
wire _3372_ ;
wire _4997_ ;
wire _4577_ ;
wire _4157_ ;
wire \genblk1[4].u_ce.LoadCtl_0_bF$buf2  ;
wire _6303_ ;
wire _2643_ ;
wire _2223_ ;
wire [1:0] \u_ot.Xin1  ;
wire _3848_ ;
wire _3428_ ;
wire _3008_ ;
wire _3181_ ;
wire _1914_ ;
wire _4386_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _6112_ ;
wire _2872_ ;
wire _2452_ ;
wire _2032_ ;
wire _3657_ ;
wire _3237_ ;
wire _5803_ ;
wire _1723_ ;
wire _1303_ ;
wire _4195_ ;
wire _634_ ;
wire _214_ ;
wire _2928_ ;
wire _2508_ ;
wire _6341_ ;
wire _2681_ ;
wire _2261_ ;
wire _3886_ ;
wire _3466_ ;
wire _3046_ ;
wire _5612_ ;
wire _1952_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _2737_ ;
wire _2317_ ;
wire _6150_ ;
wire _2490_ ;
wire _2070_ ;
wire _3695_ ;
wire _3275_ ;
wire _5841_ ;
wire _5421_ ;
wire _5001_ ;
wire _919_ ;
wire _6206_ ;
wire _1761_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _2966_ ;
wire _2546_ ;
wire _2126_ ;
wire _3084_ ;
wire _1817_ ;
wire _4289_ ;
wire _5650_ ;
wire _5230_ ;
wire _728_ ;
wire _308_ ;
wire _6015_ ;
wire _1990_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _2775_ ;
wire _2355_ ;
wire _4921_ ;
wire _4501_ ;
wire _5706_ ;
wire \genblk1[3].u_ce.Vld_bF$buf4  ;
wire _1626_ ;
wire _1206_ ;
wire _4098_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _6244_ ;
wire _290_ ;
wire _2584_ ;
wire _2164_ ;
wire _3789_ ;
wire _3369_ ;
wire _4730_ ;
wire _4310_ ;
wire _5935_ ;
wire _5515_ ;
wire _1855_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _6053_ ;
wire _2393_ ;
wire _3598_ ;
wire _3178_ ;
wire \genblk1[0].u_ce.Ain12b_11_bF$buf3  ;
wire _5744_ ;
wire _5324_ ;
wire _6109_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire _2869_ ;
wire _2449_ ;
wire _2029_ ;
wire _3810_ ;
wire _6282_ ;
wire _5276__bF$buf0 ;
wire _5276__bF$buf1 ;
wire _5276__bF$buf2 ;
wire _5276__bF$buf3 ;
wire _5276__bF$buf4 ;
wire _5973_ ;
wire _5553_ ;
wire _5133_ ;
wire _6338_ ;
wire _1893_ ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _2678_ ;
wire _2258_ ;
wire [1:0] \genblk1[3].u_ce.Yin0  ;
wire clk_bF$buf70 ;
wire clk_bF$buf71 ;
wire clk_bF$buf72 ;
wire clk_bF$buf73 ;
wire clk_bF$buf74 ;
wire clk_bF$buf75 ;
wire _6091_ ;
wire _4824_ ;
wire _4404_ ;
wire _5609_ ;
wire _1949_ ;
wire _1529_ ;
wire _1109_ ;
wire _5782_ ;
wire _5362_ ;
wire [11:0] \genblk1[1].u_ce.Ain12b  ;
wire _6147_ ;
wire _1282_ ;
wire _193_ ;
wire _2487_ ;
wire _2067_ ;
wire _4633_ ;
wire _4213_ ;
wire _5838_ ;
wire _5418_ ;
wire _1758_ ;
wire _1338_ ;
wire _5591_ ;
wire _5171_ ;
wire _669_ ;
wire _249_ ;
wire _3904_ ;
wire _1091_ ;
wire _2296_ ;
wire _4862_ ;
wire _4442_ ;
wire _4022_ ;
wire _5647_ ;
wire _5227_ ;
wire _1987_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _3713_ ;
wire \genblk1[5].u_ce.Ain12b_11_bF$buf4  ;
wire _6185_ ;
wire _4918_ ;
wire _4474__bF$buf0 ;
wire _4474__bF$buf1 ;
wire _4474__bF$buf2 ;
wire _4474__bF$buf3 ;
wire _4474__bF$buf4 ;
wire _4671_ ;
wire _4251_ ;
wire _5876_ ;
wire _5456_ ;
wire _5036_ ;
wire \genblk1[4].u_ce.ISout  ;
wire _1796_ ;
wire _1376_ ;
wire _287_ ;
wire _2851__bF$buf0 ;
wire _2851__bF$buf1 ;
wire _2851__bF$buf2 ;
wire _2851__bF$buf3 ;
wire _2851__bF$buf4 ;
wire _2851__bF$buf5 ;
wire _3942_ ;
wire _3522_ ;
wire _3102_ ;
wire _3_ ;
wire _4727_ ;
wire _4307_ ;
wire _4480_ ;
wire _4060_ ;
wire _5685_ ;
wire _5265_ ;
wire [11:0] \genblk1[3].u_ce.Ain12b  ;
wire _1185_ ;
wire _3751_ ;
wire _3331_ ;
wire _4956_ ;
wire _4536_ ;
wire _4116_ ;
wire _2602_ ;
wire _5494_ ;
wire _5074_ ;
wire _3807_ ;
wire _6279_ ;
wire _2199_ ;
wire _3980_ ;
wire _3560_ ;
wire _3140_ ;
wire _4765_ ;
wire _4345_ ;
wire _44_ ;
wire _2831_ ;
wire _2411_ ;
wire _3616_ ;
wire _6088_ ;
wire _4994_ ;
wire _4574_ ;
wire _4154_ ;
wire _5779_ ;
wire _5359_ ;
wire _6300_ ;
wire _1699_ ;
wire _1279_ ;
wire _2640_ ;
wire _2220_ ;
wire _3845_ ;
wire _3425_ ;
wire _3005_ ;
wire _1911_ ;
wire _4383_ ;
wire _822_ ;
wire _402_ ;
wire _5588_ ;
wire _5168_ ;
wire _82_ ;
wire _1088_ ;
wire [1:0] \genblk1[0].u_ce.Xin1  ;
wire [11:0] \genblk1[5].u_ce.Ain12b  ;
wire _3654_ ;
wire _3234_ ;
wire _4859_ ;
wire _4439_ ;
wire _4019_ ;
wire _5800_ ;
wire _1720_ ;
wire _1300_ ;
wire _4192_ ;
wire \genblk1[0].u_ce.ISin  ;
wire _631_ ;
wire _211_ ;
wire _2925_ ;
wire _2505_ ;
wire _5397_ ;
wire _1024__bF$buf0 ;
wire _1024__bF$buf1 ;
wire _1024__bF$buf2 ;
wire _1024__bF$buf3 ;
wire _1024__bF$buf4 ;
wire _3883_ ;
wire _3463_ ;
wire _3043_ ;
wire _4668_ ;
wire _4248_ ;
wire _860_ ;
wire _440_ ;
wire _2734_ ;
wire _2314_ ;
wire _3939_ ;
wire _3519_ ;
wire _3692_ ;
wire _3272_ ;
wire _4897_ ;
wire _4477_ ;
wire _4057_ ;
wire _916_ ;
wire _6203_ ;
wire _2963_ ;
wire _2543_ ;
wire _2123_ ;
wire _3748_ ;
wire _3328_ ;
wire _3081_ ;
wire _1814_ ;
wire _4286_ ;
wire _725_ ;
wire _305_ ;
wire _6012_ ;
wire _2772_ ;
wire _2352_ ;
wire _3977_ ;
wire _3557_ ;
wire _3137_ ;
wire _5703_ ;
wire \genblk1[3].u_ce.Vld_bF$buf1  ;
wire _1623_ ;
wire _1203_ ;
wire _4095_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _2828_ ;
wire _2408_ ;
wire _6241_ ;
wire _2581_ ;
wire _2161_ ;
wire _3786_ ;
wire _3366_ ;
wire _5932_ ;
wire _5512_ ;
wire _1852_ ;
wire _1432_ ;
wire _1012_ ;
wire _763_ ;
wire _343_ ;
wire _2637_ ;
wire _2217_ ;
wire _6050_ ;
wire [19:0] FCW ;
wire _2390_ ;
wire _3595_ ;
wire _3175_ ;
wire \genblk1[0].u_ce.Ain12b_11_bF$buf0  ;
wire _1908_ ;
wire _5741_ ;
wire _5321_ ;
wire _819_ ;
wire _79_ ;
wire _6106_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _2866_ ;
wire _2446_ ;
wire _2026_ ;
wire _1717_ ;
wire _4189_ ;
wire _5970_ ;
wire _5550_ ;
wire _5130_ ;
wire _628_ ;
wire _208_ ;
wire _6335_ ;
wire _1890_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _2675_ ;
wire _2255_ ;
wire clk_bF$buf40 ;
wire clk_bF$buf41 ;
wire clk_bF$buf42 ;
wire clk_bF$buf43 ;
wire clk_bF$buf44 ;
wire clk_bF$buf45 ;
wire clk_bF$buf46 ;
wire clk_bF$buf47 ;
wire clk_bF$buf48 ;
wire clk_bF$buf49 ;
wire _4821_ ;
wire _4401_ ;
wire _5606_ ;
wire [1:0] \genblk1[5].u_ce.Ain1  ;
wire _1946_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _6144_ ;
wire _190_ ;
wire _2484_ ;
wire _2064_ ;
wire _3689_ ;
wire _3269_ ;
wire _4630_ ;
wire _4210_ ;
wire _5835_ ;
wire _5415_ ;
wire _1755_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _3901_ ;
wire _2293_ ;
wire _3498_ ;
wire _3078_ ;
wire _5644_ ;
wire _5224_ ;
wire _6009_ ;
wire _1984_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _2769_ ;
wire _2349_ ;
wire _3710_ ;
wire \genblk1[5].u_ce.Ain12b_11_bF$buf1  ;
wire _6182_ ;
wire _4915_ ;
wire _5873_ ;
wire _5453_ ;
wire _5033_ ;
wire _6238_ ;
wire _1793_ ;
wire _1373_ ;
wire _284_ ;
wire _2998_ ;
wire _2578_ ;
wire _2158_ ;
wire _0_ ;
wire _4724_ ;
wire _4304_ ;
wire _5929_ ;
wire _5509_ ;
wire [1:0] \genblk1[6].u_ce.Xin0  ;
wire _1849_ ;
wire _1429_ ;
wire _1009_ ;
wire _5682_ ;
wire _5262_ ;
wire \genblk1[2].u_ce.LoadCtl_0_bF$buf2  ;
wire _6047_ ;
wire _1182_ ;
wire _2387_ ;
wire _4953_ ;
wire _4533_ ;
wire _4113_ ;
wire _5738_ ;
wire _5318_ ;
wire _1658_ ;
wire _1238_ ;
wire _5491_ ;
wire _5071_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire _3804_ ;
wire _6276_ ;
wire _2196_ ;
wire _4762_ ;
wire _4342_ ;
wire [11:0] \genblk1[2].u_ce.Ycalc  ;
wire _5967_ ;
wire _5547_ ;
wire _5127_ ;
wire _41_ ;
wire _1887_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _3613_ ;
wire _6085_ ;
wire _4818_ ;
wire _4991_ ;
wire _4571_ ;
wire _4151_ ;
wire _5776_ ;
wire _5356_ ;
wire _1696_ ;
wire _1276_ ;
wire _187_ ;
wire _3842_ ;
wire _3422_ ;
wire _3002_ ;
wire _4627_ ;
wire _4207_ ;
wire _4380_ ;
wire _5585_ ;
wire _5165_ ;
wire _1085_ ;
wire _3651_ ;
wire _3231_ ;
wire _4856_ ;
wire _4436_ ;
wire _4016_ ;
wire _2922_ ;
wire _2502_ ;
wire _5394_ ;
wire _3707_ ;
wire _6179_ ;
wire _2099_ ;
wire _3880_ ;
wire _3460_ ;
wire _3040_ ;
wire [11:0] \genblk1[3].u_ce.Acalc  ;
wire _4665_ ;
wire _4245_ ;
wire _2731_ ;
wire _2311_ ;
wire \genblk1[1].u_ce.Vld_bF$buf2  ;
wire _3936_ ;
wire _3516_ ;
wire _4894_ ;
wire _4474_ ;
wire _4054_ ;
wire _913_ ;
wire _5679_ ;
wire _5259_ ;
wire _6200_ ;
wire _1599_ ;
wire _1179_ ;
wire _2960_ ;
wire _2540_ ;
wire _2120_ ;
wire [1:0] \genblk1[3].u_ce.X_  ;
wire _3745_ ;
wire _3325_ ;
wire _1811_ ;
wire _4283_ ;
wire _722_ ;
wire _302_ ;
wire _5488_ ;
wire _5068_ ;
wire _3974_ ;
wire _3554_ ;
wire _3134_ ;
wire _4759_ ;
wire _4339_ ;
wire _5700_ ;
wire _38_ ;
wire _1620_ ;
wire _1200_ ;
wire _4092_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _2825_ ;
wire _2405_ ;
wire _5297_ ;
wire _3783_ ;
wire _3363_ ;
wire _4988_ ;
wire _4568_ ;
wire _4148_ ;
wire \genblk1[1].u_ce.Vld  ;
wire _760_ ;
wire _340_ ;
wire _2634_ ;
wire _2214_ ;
wire _3839_ ;
wire _3419_ ;
wire _3592_ ;
wire _3172_ ;
wire _1905_ ;
wire _4797_ ;
wire _4377_ ;
wire _816_ ;
wire _76_ ;
wire _6103_ ;
wire _2863_ ;
wire _2443_ ;
wire _2023_ ;
wire _3648_ ;
wire _3228_ ;
wire _1714_ ;
wire _4186_ ;
wire _625_ ;
wire _205_ ;
wire _2919_ ;
wire _6332_ ;
wire _2672_ ;
wire _2252_ ;
wire _5365__bF$buf0 ;
wire _5365__bF$buf1 ;
wire _5365__bF$buf2 ;
wire clk_bF$buf10 ;
wire _5365__bF$buf3 ;
wire clk_bF$buf11 ;
wire _5365__bF$buf4 ;
wire clk_bF$buf12 ;
wire _5365__bF$buf5 ;
wire clk_bF$buf13 ;
wire clk_bF$buf14 ;
wire clk_bF$buf15 ;
wire clk_bF$buf16 ;
wire clk_bF$buf17 ;
wire clk_bF$buf18 ;
wire clk_bF$buf19 ;
wire _3877_ ;
wire _3457_ ;
wire _3037_ ;
wire \genblk1[3].u_ce.Ain12b_11_bF$buf4  ;
wire _5603_ ;
wire _1943_ ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _2728_ ;
wire _2308_ ;
wire _6141_ ;
wire _2481_ ;
wire _2061_ ;
wire _3686_ ;
wire _3266_ ;
wire _5832_ ;
wire _5412_ ;
wire _1752_ ;
wire _1332_ ;
wire _663_ ;
wire _243_ ;
wire _2957_ ;
wire _2537_ ;
wire _2117_ ;
wire _2290_ ;
wire _3495_ ;
wire _3075_ ;
wire _1808_ ;
wire _5641_ ;
wire _5221_ ;
wire _719_ ;
wire _6006_ ;
wire _1981_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _2766_ ;
wire _2346_ ;
wire _4912_ ;
wire _1617_ ;
wire _4089_ ;
wire [6:0] \u_ot.ISpipe  ;
wire _5870_ ;
wire _5450_ ;
wire _5030_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _6235_ ;
wire _1790_ ;
wire _1370_ ;
wire _281_ ;
wire _2995_ ;
wire _2575_ ;
wire _2155_ ;
wire _4721_ ;
wire _4301_ ;
wire _5926_ ;
wire _5506_ ;
wire _1846_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire _6044_ ;
wire _2384_ ;
wire _3589_ ;
wire _3169_ ;
wire _4950_ ;
wire _4530_ ;
wire _4110_ ;
wire _5735_ ;
wire _5315_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire _3801_ ;
wire _6273_ ;
wire _2193_ ;
wire \genblk1[0].u_ce.Rdy  ;
wire _3398_ ;
wire _5964_ ;
wire _5544_ ;
wire _5124_ ;
wire _6329_ ;
wire _1884_ ;
wire _1464_ ;
wire _1044_ ;
wire _795_ ;
wire _375_ ;
wire _2669_ ;
wire _2249_ ;
wire _3610_ ;
wire _6082_ ;
wire _4815_ ;
wire _5773_ ;
wire _5353_ ;
wire _6138_ ;
wire _1693_ ;
wire _1273_ ;
wire _184_ ;
wire _2898_ ;
wire _2478_ ;
wire _2058_ ;
wire _4624_ ;
wire _4204_ ;
wire _5829_ ;
wire _5409_ ;
wire _1749_ ;
wire _1329_ ;
wire _5582_ ;
wire _5162_ ;
wire _1082_ ;
wire _2287_ ;
wire _4853_ ;
wire _4433_ ;
wire _4013_ ;
wire _5638_ ;
wire _5218_ ;
wire _1978_ ;
wire _1558_ ;
wire _1138_ ;
wire _5391_ ;
wire _889_ ;
wire _469_ ;
wire _3704_ ;
wire _6176_ ;
wire _4909_ ;
wire _2096_ ;
wire _4662_ ;
wire _4242_ ;
wire _5867_ ;
wire _5447_ ;
wire _5027_ ;
wire _1787_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _3933_ ;
wire _3513_ ;
wire _4718_ ;
wire _4891_ ;
wire _4471_ ;
wire _4051_ ;
wire _910_ ;
wire _5676_ ;
wire _5256_ ;
wire _1596_ ;
wire _1176_ ;
wire _3742_ ;
wire _3322_ ;
wire _4947_ ;
wire _4527_ ;
wire _4107_ ;
wire _4280_ ;
wire _5485_ ;
wire _5065_ ;
wire _3971_ ;
wire _3551_ ;
wire _3131_ ;
wire _4756_ ;
wire _4336_ ;
wire _35_ ;
wire _2822_ ;
wire _2402_ ;
wire _5294_ ;
wire _3607_ ;
wire _6079_ ;
wire _3780_ ;
wire _3360_ ;
wire _4985_ ;
wire _4565_ ;
wire _4145_ ;
wire _2631_ ;
wire _2211_ ;
wire _3836_ ;
wire _3416_ ;
wire _1902_ ;
wire _4794_ ;
wire _4374_ ;
wire _813_ ;
wire \genblk1[1].u_ce.ISout  ;
wire _5999_ ;
wire _5579_ ;
wire _5159_ ;
wire _73_ ;
wire _6100_ ;
wire _1499_ ;
wire _1079_ ;
wire _2860_ ;
wire _2440_ ;
wire _2020_ ;
wire _3645_ ;
wire _3225_ ;
wire _1711_ ;
wire _4183_ ;
wire _622_ ;
wire _202_ ;
wire _2916_ ;
wire _5388_ ;
wire [1:0] \genblk1[1].u_ce.Yin1  ;
wire _3874_ ;
wire _3454_ ;
wire _3034_ ;
wire _4659_ ;
wire \genblk1[3].u_ce.Ain12b_11_bF$buf1  ;
wire _4239_ ;
wire _5600_ ;
wire [1:0] \genblk1[4].u_ce.Ain0  ;
wire _1940_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire [11:0] \genblk1[4].u_ce.Xcalc  ;
wire _2725_ ;
wire _2305_ ;
wire _5197_ ;
wire _3683_ ;
wire _3263_ ;
wire _4888_ ;
wire _4468_ ;
wire _4048_ ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _2954_ ;
wire _2534_ ;
wire _2114_ ;
wire _3739_ ;
wire _3319_ ;
wire \genblk1[0].u_ce.LoadCtl_0_bF$buf2  ;
wire _3492_ ;
wire _3072_ ;
wire _1805_ ;
wire _4697_ ;
wire _4277_ ;
wire _716_ ;
wire _6003_ ;
wire _2763_ ;
wire _2343_ ;
wire _3968_ ;
wire _3548_ ;
wire _3128_ ;
wire _1614_ ;
wire _4086_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _2819_ ;
wire _6232_ ;
wire _2992_ ;
wire _2572_ ;
wire _2152_ ;
wire _3777_ ;
wire _3357_ ;
wire _5923_ ;
wire _5503_ ;
wire _1843_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire _2628_ ;
wire _2208_ ;
wire _6041_ ;
wire _2381_ ;
wire _3586_ ;
wire _3166_ ;
wire _5732_ ;
wire _5312_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _2857_ ;
wire _2437_ ;
wire _2017_ ;
wire _6270_ ;
wire _2190_ ;
wire _3395_ ;
wire _1708_ ;
wire _5961_ ;
wire _5541_ ;
wire _5121_ ;
wire _619_ ;
wire _6326_ ;
wire _1881_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _2666_ ;
wire _2246_ ;
wire _4812_ ;
wire _1937_ ;
wire _1517_ ;
wire _5770_ ;
wire _5350_ ;
wire _848_ ;
wire _428_ ;
wire _6135_ ;
wire _1690_ ;
wire _1270_ ;
wire _181_ ;
wire _2895_ ;
wire _2475_ ;
wire _2055_ ;
wire _4621_ ;
wire _4201_ ;
wire [6:0] \genblk1[2].u_ce.LoadCtl  ;
wire _5826_ ;
wire _5406_ ;
wire _1746_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _2284_ ;
wire _3489_ ;
wire _3069_ ;
wire _4850_ ;
wire _4430_ ;
wire _4010_ ;
wire _5635_ ;
wire _5215_ ;
wire _1975_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire \genblk1[4].u_ce.Vld_bF$buf4  ;
wire _3701_ ;
wire _6173_ ;
wire _4906_ ;
wire _2093_ ;
wire _3298_ ;
wire _5864_ ;
wire _5444_ ;
wire _5024_ ;
wire _6229_ ;
wire _1784_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _2989_ ;
wire _2569_ ;
wire _2149_ ;
wire _3930_ ;
wire _3510_ ;
wire _4715_ ;
wire _5673_ ;
wire _5253_ ;
wire _6038_ ;
wire _1593_ ;
wire _1173_ ;
wire _2798_ ;
wire _2378_ ;
wire _4944_ ;
wire _4524_ ;
wire _4104_ ;
wire _5729_ ;
wire _5309_ ;
wire _1649_ ;
wire _1229_ ;
wire _5482_ ;
wire _5062_ ;
wire _6267_ ;
wire _2187_ ;
wire _4753_ ;
wire _4333_ ;
wire _5958_ ;
wire _5538_ ;
wire _5118_ ;
wire _32_ ;
wire _1878_ ;
wire _1458_ ;
wire _1038_ ;
wire _5291_ ;
wire _789_ ;
wire _369_ ;
wire _3604_ ;
wire _6076_ ;
wire _4809_ ;
wire _4982_ ;
wire _4562_ ;
wire _4142_ ;
wire _5767_ ;
wire _5347_ ;
wire \genblk1[1].u_ce.Ain12b_11_bF$buf4  ;
wire _1687_ ;
wire _1267_ ;
wire _598_ ;
wire _178_ ;
wire _3833_ ;
wire _3413_ ;
wire _4618_ ;
wire _4791_ ;
wire _4371_ ;
wire _810_ ;
wire _5996_ ;
wire _5576_ ;
wire _5156_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _3642_ ;
wire _3222_ ;
wire [1:0] \u_ot.Yin0  ;
wire _4847_ ;
wire _4427_ ;
wire _4007_ ;
wire _4180_ ;
wire _2913_ ;
wire _5385_ ;
wire _3871_ ;
wire _3451_ ;
wire _3031_ ;
wire _4656_ ;
wire _4236_ ;
wire _2722_ ;
wire _2302_ ;
wire _5194_ ;
wire _3927_ ;
wire _3507_ ;
wire [1:0] \a[6]  ;
wire _3680_ ;
wire _3260_ ;
wire _4885_ ;
wire _4465_ ;
wire _4045_ ;
wire _904_ ;
wire _2951_ ;
wire _2531_ ;
wire _2111_ ;
wire _3736_ ;
wire _3316_ ;
wire _1802_ ;
wire _4694_ ;
wire _4274_ ;
wire [1:0] \genblk1[4].u_ce.X_  ;
wire _713_ ;
wire _5899_ ;
wire _5479_ ;
wire _5059_ ;
wire _6000_ ;
wire _1399_ ;
wire _2760_ ;
wire _2340_ ;
wire _3965_ ;
wire _3545_ ;
wire _3125_ ;
wire _29_ ;
wire _1611_ ;
wire _4083_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _2816_ ;
wire _5288_ ;
wire _3774_ ;
wire _3354_ ;
wire _4979_ ;
wire _4559_ ;
wire _4139_ ;
wire _5920_ ;
wire _5500_ ;
wire _1840_ ;
wire _1420_ ;
wire _1000_ ;
wire [1:0] \genblk1[4].u_ce.Xin1  ;
wire _751_ ;
wire _331_ ;
wire _2625_ ;
wire _2205_ ;
wire _5097_ ;
wire [11:0] \genblk1[0].u_ce.Acalc  ;
wire _3583_ ;
wire _3163_ ;
wire _4788_ ;
wire _4368_ ;
wire _807_ ;
wire _67_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _2854_ ;
wire _2434_ ;
wire _2014_ ;
wire _3639_ ;
wire _3219_ ;
wire _3392_ ;
wire _1705_ ;
wire _4597_ ;
wire _4177_ ;
wire _616_ ;
wire _6323_ ;
wire _2663_ ;
wire _2243_ ;
wire _3868_ ;
wire _3448_ ;
wire _3028_ ;
wire _1934_ ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _2719_ ;
wire _6132_ ;
wire _2892_ ;
wire _2472_ ;
wire _2052_ ;
wire _3677_ ;
wire _3257_ ;
wire _5823_ ;
wire _5403_ ;
wire _1743_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire _2948_ ;
wire _2528_ ;
wire _2108_ ;
wire _2281_ ;
wire _3486_ ;
wire _3066_ ;
wire _5632_ ;
wire _5212_ ;
wire _1972_ ;
wire _1552_ ;
wire _1132_ ;
wire \genblk1[5].u_ce.LoadCtl_0_bF$buf2  ;
wire _883_ ;
wire _463_ ;
wire _2757_ ;
wire _2337_ ;
wire \genblk1[4].u_ce.Vld_bF$buf1  ;
wire _6170_ ;
wire _4903_ ;
wire _2090_ ;
wire _3295_ ;
wire _1608_ ;
wire _5861_ ;
wire _5441_ ;
wire _5021_ ;
wire _939_ ;
wire _519_ ;
wire _6226_ ;
wire _1781_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _4569__bF$buf0 ;
wire _4569__bF$buf1 ;
wire _4569__bF$buf2 ;
wire _4569__bF$buf3 ;
wire _2986_ ;
wire _4569__bF$buf4 ;
wire _2566_ ;
wire _4569__bF$buf5 ;
wire _2146_ ;
wire _4712_ ;
wire _5917_ ;
wire _1837_ ;
wire _1417_ ;
wire _5670_ ;
wire _5250_ ;
wire _748_ ;
wire _328_ ;
wire _6035_ ;
wire _1590_ ;
wire _1170_ ;
wire _2795_ ;
wire _2375_ ;
wire [11:0] \genblk1[0].u_ce.Ain12b  ;
wire _4941_ ;
wire _4521_ ;
wire _4101_ ;
wire _5726_ ;
wire _5306_ ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire _6264_ ;
wire _2184_ ;
wire _3389_ ;
wire _4750_ ;
wire _4330_ ;
wire _5955_ ;
wire _5535_ ;
wire _5115_ ;
wire _1875_ ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _3601_ ;
wire _6073_ ;
wire _4806_ ;
wire _3198_ ;
wire _5764_ ;
wire _5344_ ;
wire \genblk1[1].u_ce.Ain12b_11_bF$buf1  ;
wire _6129_ ;
wire _1684_ ;
wire _1264_ ;
wire _595_ ;
wire _175_ ;
wire _2889_ ;
wire _2469_ ;
wire _2049_ ;
wire _3830_ ;
wire _3410_ ;
wire _4615_ ;
wire _5993_ ;
wire _5573_ ;
wire _5153_ ;
wire _1493_ ;
wire _1073_ ;
wire _2698_ ;
wire _2278_ ;
wire _4844_ ;
wire _4424_ ;
wire _4004_ ;
wire [11:0] \genblk1[2].u_ce.Ain12b  ;
wire _5629_ ;
wire _5209_ ;
wire _1969_ ;
wire _1549_ ;
wire _1129_ ;
wire _2910_ ;
wire _5382_ ;
wire _6167_ ;
wire _2087_ ;
wire [11:0] \genblk1[6].u_ce.Ycalc  ;
wire [1:0] \genblk1[0].u_ce.Yin0  ;
wire _4653_ ;
wire _4233_ ;
wire _5858_ ;
wire _5438_ ;
wire _5018_ ;
wire _1778_ ;
wire _1358_ ;
wire _5191_ ;
wire _689_ ;
wire _269_ ;
wire _3924_ ;
wire _3504_ ;
wire _4709_ ;
wire _4882_ ;
wire _4462_ ;
wire _4042_ ;
wire _901_ ;
wire _5667_ ;
wire _5247_ ;
wire _1587_ ;
wire _1167_ ;
wire _498_ ;
wire _3733_ ;
wire _3313_ ;
wire _4938_ ;
wire _4518_ ;
wire \genblk1[6].u_ce.Ain12b_11_bF$buf2  ;
wire _4691_ ;
wire _4271_ ;
wire _710_ ;
wire _5896_ ;
wire _5476_ ;
wire _5056_ ;
wire _1396_ ;
wire _3962_ ;
wire _3542_ ;
wire _3122_ ;
wire _4747_ ;
wire _4327_ ;
wire [11:0] \genblk1[4].u_ce.Ain12b  ;
wire _26_ ;
wire _4080_ ;
wire _2813_ ;
wire _5285_ ;
wire \genblk1[3].u_ce.LoadCtl_0_bF$buf3  ;
wire _3771_ ;
wire _3351_ ;
wire _4976_ ;
wire _4556_ ;
wire _4136_ ;
wire _2622_ ;
wire _2202_ ;
wire _5094_ ;
wire _3827_ ;
wire _3407_ ;
wire _6299_ ;
wire _3580_ ;
wire _3160_ ;
wire _4785_ ;
wire _4365_ ;
wire _804_ ;
wire _64_ ;
wire _2851_ ;
wire _2431_ ;
wire _2011_ ;
wire _3636_ ;
wire _3216_ ;
wire _1702_ ;
wire _4594_ ;
wire _4174_ ;
wire _613_ ;
wire _2907_ ;
wire _5799_ ;
wire _5379_ ;
wire _6320_ ;
wire _1299_ ;
wire _2660_ ;
wire _2240_ ;
wire _3865_ ;
wire _3445_ ;
wire _3025_ ;
wire _1931_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _2716_ ;
wire _5188_ ;
wire _3674_ ;
wire _3254_ ;
wire _4879_ ;
wire _4459_ ;
wire _4039_ ;
wire _5820_ ;
wire _5400_ ;
wire _1740_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire _2945_ ;
wire _2525_ ;
wire _2105_ ;
wire _3483_ ;
wire _3063_ ;
wire _4688_ ;
wire _4268_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _2754_ ;
wire _2334_ ;
wire _3959_ ;
wire _3539_ ;
wire _3119_ ;
wire _4900_ ;
wire \genblk1[2].u_ce.Vld_bF$buf4  ;
wire [11:0] \genblk1[2].u_ce.Xin12b  ;
wire _3292_ ;
wire _1605_ ;
wire _4497_ ;
wire _4077_ ;
wire _936_ ;
wire _516_ ;
wire _6223_ ;
wire _2983_ ;
wire _2563_ ;
wire _2143_ ;
wire _3768_ ;
wire _3348_ ;
wire _5914_ ;
wire _1834_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _2619_ ;
wire _6032_ ;
wire _2792_ ;
wire _2372_ ;
wire _3997_ ;
wire _3577_ ;
wire _3157_ ;
wire _5723_ ;
wire _5303_ ;
wire _1643_ ;
wire _1223_ ;
wire [11:0] \genblk1[1].u_ce.Xcalc  ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire _2848_ ;
wire _2428_ ;
wire _2008_ ;
wire _6261_ ;
wire _2181_ ;
wire _3386_ ;
wire _5952_ ;
wire _5532_ ;
wire _5112_ ;
wire _6317_ ;
wire _1872_ ;
wire _1452_ ;
wire _1032_ ;
wire _783_ ;
wire _363_ ;
wire _2657_ ;
wire _2237_ ;
wire _6070_ ;
wire _4803_ ;
wire _3195_ ;
wire [11:0] \genblk1[4].u_ce.Xin12b  ;
wire _1928_ ;
wire _1508_ ;
wire _5761_ ;
wire _5341_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _6126_ ;
wire _1681_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _2886_ ;
wire _2466_ ;
wire _2046_ ;
wire _4612_ ;
wire _5817_ ;
wire _1737_ ;
wire _1317_ ;
wire Vld ;
wire _5990_ ;
wire _5570_ ;
wire _5150_ ;
wire _648_ ;
wire _228_ ;
wire _1490_ ;
wire _1070_ ;
wire _2695_ ;
wire _2275_ ;
wire _4841_ ;
wire _4421_ ;
wire _4001_ ;
wire _5626_ ;
wire _5206_ ;
wire _1966_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _6164_ ;
wire _2084_ ;
wire _3289_ ;
wire _4650_ ;
wire _4230_ ;
wire _5855_ ;
wire _5435_ ;
wire _5015_ ;
wire [1:0] \genblk1[2].u_ce.Ain1  ;
wire _1775_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire _3921_ ;
wire _3501_ ;
wire _4706_ ;
wire _3098_ ;
wire [11:0] \genblk1[6].u_ce.Xin12b  ;
wire _5664_ ;
wire _5244_ ;
wire _6029_ ;
wire _1584_ ;
wire _1164_ ;
wire _495_ ;
wire _2789_ ;
wire _2369_ ;
wire _3730_ ;
wire _3310_ ;
wire _4935_ ;
wire _4515_ ;
wire _5893_ ;
wire _5473_ ;
wire _5053_ ;
wire _6258_ ;
wire _1393_ ;
wire _2598_ ;
wire _2178_ ;
wire _4744_ ;
wire _4324_ ;
wire _5949_ ;
wire _5529_ ;
wire _5109_ ;
wire _23_ ;
wire _1869_ ;
wire _1449_ ;
wire _1029_ ;
wire _2810_ ;
wire _5282_ ;
wire _6067_ ;
wire \genblk1[3].u_ce.LoadCtl_0_bF$buf0  ;
wire _4973_ ;
wire _4553_ ;
wire _4133_ ;
wire _5758_ ;
wire _5338_ ;
wire _1678_ ;
wire _1258_ ;
wire [1:0] \genblk1[3].u_ce.Xin0  ;
wire _5091_ ;
wire _589_ ;
wire _169_ ;
wire _3824_ ;
wire _3404_ ;
wire _6296_ ;
wire _4609_ ;
wire _4782_ ;
wire _4362_ ;
wire _801_ ;
wire _5987_ ;
wire _5567_ ;
wire _5147_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _398_ ;
wire _3633_ ;
wire _3213_ ;
wire _4838_ ;
wire _4418_ ;
wire _4591_ ;
wire _4171_ ;
wire _610_ ;
wire _2904_ ;
wire _5796_ ;
wire _5376_ ;
wire _1296_ ;
wire _3862_ ;
wire _3442_ ;
wire _3022_ ;
wire _4647_ ;
wire _4227_ ;
wire _2713_ ;
wire _5185_ ;
wire _3918_ ;
wire _3671_ ;
wire _3251_ ;
wire _4876_ ;
wire _4456_ ;
wire _4036_ ;
wire _2942_ ;
wire _2522_ ;
wire _2102_ ;
wire _3727_ ;
wire _3307_ ;
wire _6199_ ;
wire _3480_ ;
wire _3060_ ;
wire _4685_ ;
wire _4265_ ;
wire _704_ ;
wire _2751_ ;
wire _2331_ ;
wire _3956_ ;
wire _3536_ ;
wire _3116_ ;
wire \genblk1[2].u_ce.Vld_bF$buf1  ;
wire [1:0] \genblk1[5].u_ce.X_  ;
wire _1602_ ;
wire _4494_ ;
wire _4074_ ;
wire _933_ ;
wire _513_ ;
wire _2807_ ;
wire _5699_ ;
wire _5279_ ;
wire _6220_ ;
wire _1199_ ;
wire _2980_ ;
wire _2560_ ;
wire _2140_ ;
wire _3765_ ;
wire _3345_ ;
wire _5911_ ;
wire _1831_ ;
wire _1411_ ;
wire _742_ ;
wire _322_ ;
wire _2616_ ;
wire _5088_ ;
wire _3994_ ;
wire _3574_ ;
wire _3154_ ;
wire _4779_ ;
wire _4359_ ;
wire _5720_ ;
wire _5300_ ;
wire _58_ ;
wire _1640_ ;
wire _1220_ ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _2845_ ;
wire [1:0] \genblk1[5].u_ce.Yin1  ;
wire _2425_ ;
wire _2005_ ;
wire _3383_ ;
wire _4588_ ;
wire _4168_ ;
wire _607_ ;
wire _6314_ ;
wire _780_ ;
wire _360_ ;
wire _2654_ ;
wire _2234_ ;
wire _3859_ ;
wire _3439_ ;
wire _3019_ ;
wire _4800_ ;
wire _3192_ ;
wire _1925_ ;
wire _1505_ ;
wire _4397_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _6123_ ;
wire _2883_ ;
wire _2463_ ;
wire _2043_ ;
wire _3668_ ;
wire _3248_ ;
wire _5814_ ;
wire _1734_ ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire _2939_ ;
wire _2519_ ;
wire _2692_ ;
wire _2272_ ;
wire _3897_ ;
wire _3477_ ;
wire _3057_ ;
wire _5623_ ;
wire _5203_ ;
wire _1963_ ;
wire _1543_ ;
wire \genblk1[4].u_ce.Ain12b_11_bF$buf2  ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _2748_ ;
wire _2328_ ;
wire _6161_ ;
wire _2081_ ;
wire _3286_ ;
wire _5852_ ;
wire _5432_ ;
wire _5012_ ;
wire _6217_ ;
wire _1772_ ;
wire _1352_ ;
wire _683_ ;
wire _263_ ;
wire _2977_ ;
wire _2557_ ;
wire _2137_ ;
wire _4703_ ;
wire _5908_ ;
wire _3095_ ;
wire \genblk1[1].u_ce.LoadCtl_0_bF$buf3  ;
wire _1828_ ;
wire _1408_ ;
wire _5661_ ;
wire _5241_ ;
wire _739_ ;
wire _319_ ;
wire _6026_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _2786_ ;
wire _2366_ ;
wire _4932_ ;
wire _4512_ ;
wire _5717_ ;
wire _1637_ ;
wire _1217_ ;
wire _5890_ ;
wire _5470_ ;
wire _5050_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _6255_ ;
wire _1390_ ;
wire _2595_ ;
wire _2175_ ;
wire _4741_ ;
wire _4321_ ;
wire _5946_ ;
wire _5526_ ;
wire _5106_ ;
wire _20_ ;
wire _1866_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire _6064_ ;
wire _3189_ ;
wire _4970_ ;
wire _4550_ ;
wire _4130_ ;
wire _5755_ ;
wire _5335_ ;
wire _1675_ ;
wire _1255_ ;
wire _586_ ;
wire _166_ ;
wire _3821_ ;
wire _3401_ ;
wire _6293_ ;
wire _4606_ ;
wire _5984_ ;
wire _5564_ ;
wire _5144_ ;
wire _1484_ ;
wire _1064_ ;
wire _395_ ;
wire [1:0] \a[1]  ;
wire _2689_ ;
wire _2269_ ;
wire _164__bF$buf0 ;
wire _164__bF$buf1 ;
wire _164__bF$buf2 ;
wire _164__bF$buf3 ;
wire _164__bF$buf4 ;
wire _3630_ ;
wire _3210_ ;
wire _4835_ ;
wire _4415_ ;
wire _2901_ ;
wire _5793_ ;
wire _5373_ ;
wire _6158_ ;
wire _1293_ ;
wire _2498_ ;
wire _2078_ ;
wire _4644_ ;
wire _4224_ ;
wire _5849_ ;
wire _5429_ ;
wire _5009_ ;
wire \genblk1[0].u_ce.Vld_bF$buf2  ;
wire _1769_ ;
wire _1349_ ;
wire _2710_ ;
wire _5182_ ;
wire _3915_ ;
wire _4873_ ;
wire _4453_ ;
wire _4033_ ;
wire _5658_ ;
wire _5238_ ;
wire _1998_ ;
wire _1578_ ;
wire _1158_ ;
wire _489_ ;
wire _3724_ ;
wire _3304_ ;
wire _6196_ ;
wire _4929_ ;
wire _4509_ ;
wire _4682_ ;
wire _4262_ ;
wire _701_ ;
wire _5887_ ;
wire _5467_ ;
wire _5047_ ;
wire _1387_ ;
wire _298_ ;
wire _3953_ ;
wire _3533_ ;
wire _3113_ ;
wire _4738_ ;
wire _4318_ ;
wire _17_ ;
wire _4491_ ;
wire _4071_ ;
wire _930_ ;
wire _510_ ;
wire _2804_ ;
wire _5696_ ;
wire _5276_ ;
wire _1196_ ;
wire _3762_ ;
wire _3342_ ;
wire _4967_ ;
wire _4547_ ;
wire _4127_ ;
wire _2613_ ;
wire _5085_ ;
wire _3818_ ;
wire [11:0] \genblk1[3].u_ce.Ycalc  ;
wire _3991_ ;
wire _3571_ ;
wire _3151_ ;
wire _4776_ ;
wire _4356_ ;
wire _55_ ;
wire _2842_ ;
wire _2422_ ;
wire _2002_ ;
wire _3627_ ;
wire _3207_ ;
wire _6099_ ;
wire _3380_ ;
wire _4585_ ;
wire _4165_ ;
wire _604_ ;
wire _6311_ ;
wire _2651_ ;
wire _2231_ ;
wire \u_ot.ISout_bF$buf3  ;
wire _3856_ ;
wire _3436_ ;
wire _3016_ ;
wire _1922_ ;
wire _1502_ ;
wire _4394_ ;
wire _833_ ;
wire _413_ ;
wire _2707_ ;
wire _5599_ ;
wire _5179_ ;
wire _93_ ;
wire _6120_ ;
wire _1099_ ;
wire _2880_ ;
wire _2460_ ;
wire _2040_ ;
wire _3665_ ;
wire _3245_ ;
wire _5811_ ;
wire _1731_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _2936_ ;
wire _2516_ ;
wire [11:0] \genblk1[4].u_ce.Acalc  ;
wire _3894_ ;
wire _3474_ ;
wire _3054_ ;
wire [6:0] \genblk1[4].u_ce.LoadCtl  ;
wire _4679_ ;
wire _4259_ ;
wire _5620_ ;
wire _5200_ ;
wire _1960_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _2745_ ;
wire _2325_ ;
wire _3283_ ;
wire _4488_ ;
wire _4068_ ;
wire _927_ ;
wire _507_ ;
wire _6214_ ;
wire [1:0] \genblk1[1].u_ce.Ain0  ;
wire _680_ ;
wire _260_ ;
wire _2974_ ;
wire _2554_ ;
wire _2134_ ;
wire _3759_ ;
wire _3339_ ;
wire _4700_ ;
wire _5905_ ;
wire _3092_ ;
wire \genblk1[1].u_ce.LoadCtl_0_bF$buf0  ;
wire _1825_ ;
wire _1405_ ;
wire _4297_ ;
wire _736_ ;
wire _316_ ;
wire _6023_ ;
wire _2783_ ;
wire _2363_ ;
wire _3988_ ;
wire _3568_ ;
wire _3148_ ;
wire _5714_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _2839_ ;
wire _2419_ ;
wire _6252_ ;
wire _2592_ ;
wire _2172_ ;
wire _3797_ ;
wire _3377_ ;
wire _5943_ ;
wire _5523_ ;
wire _5103_ ;
wire _6308_ ;
wire _1863_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _2648_ ;
wire _2228_ ;
wire _6061_ ;
wire _3186_ ;
wire _1919_ ;
wire _5752_ ;
wire _5332_ ;
wire _6117_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _2877_ ;
wire _2457_ ;
wire _2037_ ;
wire _6290_ ;
wire _4603_ ;
wire _5808_ ;
wire _1728_ ;
wire _1308_ ;
wire _5981_ ;
wire _5561_ ;
wire _5141_ ;
wire _639_ ;
wire _219_ ;
wire _6346_ ;
wire _1481_ ;
wire _1061_ ;
wire _392_ ;
wire _2686_ ;
wire _2266_ ;
wire _4832_ ;
wire _4412_ ;
wire _5617_ ;
wire _1957_ ;
wire _1537_ ;
wire _1117_ ;
wire _5790_ ;
wire _5370_ ;
wire _868_ ;
wire _448_ ;
wire _6155_ ;
wire _1290_ ;
wire _2495_ ;
wire _2075_ ;
wire _4641_ ;
wire _4221_ ;
wire [11:0] _5846_ ;
wire _5426_ ;
wire _5006_ ;
wire _1766_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _3912_ ;
wire _3089_ ;
wire _4870_ ;
wire _4450_ ;
wire _4030_ ;
wire _5655_ ;
wire _5235_ ;
wire _1995_ ;
wire _1575_ ;
wire _1155_ ;
wire _486_ ;
wire _3721_ ;
wire _3301_ ;
wire _6193_ ;
wire \genblk1[6].u_ce.LoadCtl_0_bF$buf3  ;
wire _4926_ ;
wire _4506_ ;
wire \genblk1[5].u_ce.Vld_bF$buf3  ;
wire _5884_ ;
wire _5464_ ;
wire _5044_ ;
wire _6249_ ;
wire _1384_ ;
wire _295_ ;
wire _2589_ ;
wire _2169_ ;
wire _3950_ ;
wire _3530_ ;
wire _3110_ ;
wire _4735_ ;
wire _4315_ ;
wire _14_ ;
wire _2801_ ;
wire _5693_ ;
wire _5273_ ;
wire _6058_ ;
wire _1193_ ;
wire _2398_ ;
wire _4964_ ;
wire _4544_ ;
wire _4124_ ;
wire _5749_ ;
wire _5329_ ;
wire _1669_ ;
wire _1249_ ;
wire _2610_ ;
wire _5082_ ;
wire _3815_ ;
wire _6287_ ;
wire _4773_ ;
wire _4353_ ;
wire _5978_ ;
wire _5558_ ;
wire _5138_ ;
wire _52_ ;
wire _1898_ ;
wire _1478_ ;
wire _1058_ ;
wire [1:0] \genblk1[4].u_ce.Yin0  ;
wire _389_ ;
wire _3624_ ;
wire _3204_ ;
wire _6096_ ;
wire _4829_ ;
wire _4409_ ;
wire _4582_ ;
wire _4162_ ;
wire _601_ ;
wire _5787_ ;
wire _5367_ ;
wire _1287_ ;
wire _198_ ;
wire \u_ot.ISout_bF$buf0  ;
wire \genblk1[2].u_ce.Ain12b_11_bF$buf2  ;
wire _3853_ ;
wire _3433_ ;
wire _3013_ ;
wire _4638_ ;
wire _4218_ ;
wire _4391_ ;
wire _830_ ;
wire _410_ ;
wire _2704_ ;
wire _5596_ ;
wire _5176_ ;
wire _90_ ;
wire _3909_ ;
wire _1096_ ;
wire _3662_ ;
wire _3242_ ;
wire _4867_ ;
wire _4447_ ;
wire _4027_ ;
wire _2933_ ;
wire _2513_ ;
wire _3718_ ;
wire _3891_ ;
wire _3471_ ;
wire _3051_ ;
wire _4676_ ;
wire _4256_ ;
wire _2742_ ;
wire _2322_ ;
wire _3947_ ;
wire _3527_ ;
wire _3107_ ;
wire _8_ ;
wire _3280_ ;
wire _4485_ ;
wire _4065_ ;
wire _924_ ;
wire _504_ ;
wire _6211_ ;
wire [1:0] \genblk1[6].u_ce.X_  ;
wire _2971_ ;
wire _2551_ ;
wire _2131_ ;
wire _3756_ ;
wire _3336_ ;
wire [11:0] \u_ot.Ycalc  ;
wire _5902_ ;
wire _1822_ ;
wire _1402_ ;
wire _4294_ ;
wire _733_ ;
wire _313_ ;
wire _2607_ ;
wire _5499_ ;
wire _5079_ ;
wire _6020_ ;
wire _2780_ ;
wire _2360_ ;
wire _3985_ ;
wire _3565_ ;
wire _3145_ ;
wire _1057__bF$buf0 ;
wire _5711_ ;
wire _1057__bF$buf1 ;
wire _1057__bF$buf2 ;
wire _1057__bF$buf3 ;
wire _49_ ;
wire _1631_ ;
wire _1211_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _2836_ ;
wire _2416_ ;
wire _3794_ ;
wire _3374_ ;
wire _4999_ ;
wire _4579_ ;
wire _4159_ ;
wire _5940_ ;
wire \genblk1[4].u_ce.LoadCtl_0_bF$buf4  ;
wire _5520_ ;
wire _5100_ ;
wire _6305_ ;
wire _1860_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _2645_ ;
wire _2225_ ;
wire _3183_ ;
wire _1916_ ;
wire _4388_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _6114_ ;
wire [1:0] \genblk1[1].u_ce.Xin1  ;
wire _580_ ;
wire _160_ ;
wire _2874_ ;
wire _2454_ ;
wire _2034_ ;
wire _3659_ ;
wire _3239_ ;
wire _4600_ ;
wire _5805_ ;
wire _1725_ ;
wire _1305_ ;
wire _4197_ ;
wire _636_ ;
wire _216_ ;
wire _6343_ ;
wire _2683_ ;
wire _2263_ ;
wire _3888_ ;
wire _3468_ ;
wire _3048_ ;
wire _5614_ ;
wire _1954_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _2739_ ;
wire _2319_ ;
wire _6152_ ;
wire _253__bF$buf0 ;
wire _253__bF$buf1 ;
wire _253__bF$buf2 ;
wire _253__bF$buf3 ;
wire _253__bF$buf4 ;
wire _253__bF$buf5 ;
wire _2492_ ;
wire _2072_ ;
wire _3697_ ;
wire _3277_ ;
wire _5843_ ;
wire _5423_ ;
wire _5003_ ;
wire _6208_ ;
wire _1763_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _2968_ ;
wire _2548_ ;
wire _2128_ ;
wire _3086_ ;
wire _1819_ ;
wire _5652_ ;
wire _5232_ ;
wire _6017_ ;
wire _1992_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire _2777_ ;
wire _2357_ ;
wire _6190_ ;
wire \genblk1[6].u_ce.LoadCtl_0_bF$buf0  ;
wire _4923_ ;
wire _4503_ ;
wire \genblk1[5].u_ce.Vld_bF$buf0  ;
wire _5708_ ;
wire _1628_ ;
wire _1208_ ;
wire _5881_ ;
wire _5461_ ;
wire _5041_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _6246_ ;
wire _1381_ ;
wire _292_ ;
wire _2586_ ;
wire _2166_ ;
wire _4732_ ;
wire _4312_ ;
wire _6047__bF$buf0 ;
wire _6047__bF$buf1 ;
wire _6047__bF$buf2 ;
wire _6047__bF$buf3 ;
wire _5937_ ;
wire _5517_ ;
wire _11_ ;
wire _1857_ ;
wire _1437_ ;
wire _1017_ ;
wire _5690_ ;
wire _5270_ ;
wire _768_ ;
wire _348_ ;
wire _6055_ ;
wire _1190_ ;
wire _2395_ ;
wire _4961_ ;
wire _4541_ ;
wire _4121_ ;
wire _5746_ ;
wire _5326_ ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _3812_ ;
wire _6284_ ;
wire _4770_ ;
wire _4350_ ;
wire _5975_ ;
wire _5555_ ;
wire _5135_ ;
wire _1895_ ;
wire _1475_ ;
wire _1055_ ;
wire _386_ ;
wire _3621_ ;
wire _3201_ ;
wire _6093_ ;
wire _4826_ ;
wire _4406_ ;
wire _5784_ ;
wire _5364_ ;
wire _6149_ ;
wire _1284_ ;
wire _195_ ;
wire _2489_ ;
wire _2069_ ;
wire _3850_ ;
wire _3430_ ;
wire _3010_ ;
wire _4635_ ;
wire _4215_ ;
wire _2701_ ;
wire _5593_ ;
wire _5173_ ;
wire _3906_ ;
wire _1093_ ;
wire _2298_ ;
wire _3622__bF$buf0 ;
wire _3622__bF$buf1 ;
wire _3622__bF$buf2 ;
wire _3622__bF$buf3 ;
wire _3622__bF$buf4 ;
wire _4864_ ;
wire _4444_ ;
wire _4024_ ;
wire _5649_ ;
wire _5229_ ;
wire _1989_ ;
wire _1569_ ;
wire _1149_ ;
wire _2930_ ;
wire _2510_ ;
wire _3715_ ;
wire _6187_ ;
wire _4673_ ;
wire _4253_ ;
wire _5878_ ;
wire _5458_ ;
wire _5038_ ;
wire _1798_ ;
wire _1378_ ;
wire _289_ ;
wire _3944_ ;
wire _3524_ ;
wire _3104_ ;
wire _5_ ;
wire _4729_ ;
wire _4309_ ;
wire _4482_ ;
wire _4062_ ;
wire _921_ ;
wire _501_ ;
wire _5687_ ;
wire _5267_ ;
wire _1187_ ;
wire _3753_ ;
wire _3333_ ;
wire _4958_ ;
wire _4538_ ;
wire _4118_ ;
wire _4291_ ;
wire _730_ ;
wire _310_ ;
wire _2604_ ;
wire _5496_ ;
wire _5076_ ;
wire _3809_ ;
wire _3982_ ;
wire _3562_ ;
wire _3142_ ;
wire _4767_ ;
wire _4347_ ;
wire _46_ ;
wire _2833_ ;
wire _2413_ ;
wire _3618_ ;
wire _3791_ ;
wire _3371_ ;
wire _4996_ ;
wire _4576_ ;
wire _4156_ ;
wire \genblk1[4].u_ce.LoadCtl_0_bF$buf1  ;
wire _6302_ ;
wire _2642_ ;
wire _2222_ ;
wire [1:0] \u_ot.Xin0  ;
wire _3847_ ;
wire _3427_ ;
wire _3007_ ;
wire _3180_ ;
wire _1913_ ;
wire _4385_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _6111_ ;
wire [11:0] \genblk1[1].u_ce.Xin12b  ;
wire _2871_ ;
wire _2451_ ;
wire _2031_ ;
wire _3656_ ;
wire _3236_ ;
wire _5802_ ;
wire _1722_ ;
wire _1302_ ;
wire _4194_ ;
wire _633_ ;
wire _213_ ;
wire _2927_ ;
wire _2507_ ;
wire _5399_ ;
wire _6340_ ;
wire _2680_ ;
wire _2260_ ;
wire _3885_ ;
wire _3465_ ;
wire _3045_ ;
wire _5611_ ;
wire _1951_ ;
wire _1531_ ;
wire _1111_ ;
wire _862_ ;
wire _442_ ;
wire _2736_ ;
wire _2316_ ;
wire [11:0] \genblk1[0].u_ce.Ycalc  ;
wire _3694_ ;
wire _3274_ ;
wire _4899_ ;
wire _4479_ ;
wire _4059_ ;
wire _5840_ ;
wire _5420_ ;
wire _5000_ ;
wire _918_ ;
wire _6205_ ;
wire _1760_ ;
wire _1340_ ;
wire _671_ ;
wire _251_ ;
wire _2965_ ;
wire _2545_ ;
wire _2125_ ;
wire _6133__bF$buf0 ;
wire _6133__bF$buf1 ;
wire _6133__bF$buf2 ;
wire _6133__bF$buf3 ;
wire _3083_ ;
wire _1816_ ;
wire _4288_ ;
wire _727_ ;
wire _307_ ;
wire _6014_ ;
wire [11:0] \genblk1[3].u_ce.Xin12b  ;
wire _480_ ;
wire _2774_ ;
wire _2354_ ;
wire _3979_ ;
wire _3559_ ;
wire _3139_ ;
wire _4920_ ;
wire _4500_ ;
wire _5705_ ;
wire \genblk1[3].u_ce.Vld_bF$buf3  ;
wire _1625_ ;
wire _1205_ ;
wire _4097_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _6243_ ;
wire _2583_ ;
wire _2163_ ;
wire _3788_ ;
wire _3368_ ;
wire _5934_ ;
wire _5514_ ;
wire _1854_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _2639_ ;
wire _2219_ ;
wire [11:0] \genblk1[1].u_ce.Acalc  ;
wire _6052_ ;
wire _2392_ ;
wire _3597_ ;
wire _3177_ ;
wire \genblk1[0].u_ce.Ain12b_11_bF$buf2  ;
wire _5743_ ;
wire _5323_ ;
wire _6108_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _2868_ ;
wire _2448_ ;
wire _2028_ ;
wire _6281_ ;
wire _1719_ ;
wire _5972_ ;
wire _5552_ ;
wire _5132_ ;
wire _6337_ ;
wire _1892_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _2677_ ;
wire _2257_ ;
wire clk_bF$buf60 ;
wire clk_bF$buf61 ;
wire clk_bF$buf62 ;
wire clk_bF$buf63 ;
wire clk_bF$buf64 ;
wire clk_bF$buf65 ;
wire clk_bF$buf66 ;
wire clk_bF$buf67 ;
wire clk_bF$buf68 ;
wire clk_bF$buf69 ;
wire [11:0] \genblk1[5].u_ce.Xin12b  ;
wire _6090_ ;
wire _4823_ ;
wire _4403_ ;
wire _5608_ ;
wire _1948_ ;
wire _1528_ ;
wire _1108_ ;
wire _5781_ ;
wire _5361_ ;
wire _859_ ;
wire _439_ ;
wire _6146_ ;
wire _1281_ ;
wire _192_ ;
wire _2486_ ;
wire _2066_ ;
wire _4632_ ;
wire _4212_ ;
wire _5837_ ;
wire _5417_ ;
wire _1757_ ;
wire _1337_ ;
wire _5590_ ;
wire _5170_ ;
wire _668_ ;
wire _248_ ;
wire _3903_ ;
wire _1090_ ;
wire _2295_ ;
wire _4861_ ;
wire _4441_ ;
wire _4021_ ;
wire _5646_ ;
wire _5226_ ;
wire _1986_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _3712_ ;
wire \genblk1[5].u_ce.Ain12b_11_bF$buf3  ;
wire _6184_ ;
wire _4917_ ;
wire _2756__bF$buf0 ;
wire _2756__bF$buf1 ;
wire _2756__bF$buf2 ;
wire _2756__bF$buf3 ;
wire _2756__bF$buf4 ;
wire _4670_ ;
wire _4250_ ;
wire _5875_ ;
wire _5455_ ;
wire _5035_ ;
wire _1795_ ;
wire _1375_ ;
wire _286_ ;
wire _3941_ ;
wire _3521_ ;
wire _3101_ ;
wire _2_ ;
wire _4726_ ;
wire _4306_ ;
wire _5684_ ;
wire _5264_ ;
wire \genblk1[2].u_ce.LoadCtl_0_bF$buf4  ;
wire _6049_ ;
wire _1184_ ;
wire _2389_ ;
wire _3750_ ;
wire _3330_ ;
wire _4955_ ;
wire _4535_ ;
wire _4115_ ;
wire _2601_ ;
wire _5493_ ;
wire _5073_ ;
wire _3806_ ;
wire _6278_ ;
wire _2198_ ;
wire _4764_ ;
wire _4344_ ;
wire _5969_ ;
wire _5549_ ;
wire _5129_ ;
wire _43_ ;
wire _1889_ ;
wire _1469_ ;
wire _1049_ ;
wire _2830_ ;
wire _2410_ ;
wire _3615_ ;
wire _6087_ ;
wire _4993_ ;
wire _4573_ ;
wire _4153_ ;
wire _5778_ ;
wire _5358_ ;
wire _1698_ ;
wire _1278_ ;
wire _189_ ;
wire _3844_ ;
wire _3424_ ;
wire _3004_ ;
wire _4629_ ;
wire _4209_ ;
wire _1910_ ;
wire _4382_ ;
wire _821_ ;
wire _401_ ;
wire _5587_ ;
wire _5167_ ;
wire _81_ ;
wire _1087_ ;
wire [1:0] \genblk1[0].u_ce.Xin0  ;
wire _3653_ ;
wire _3233_ ;
wire _4858_ ;
wire _4438_ ;
wire _4018_ ;
wire _4191_ ;
wire _630_ ;
wire _210_ ;
wire _2924_ ;
wire _2504_ ;
wire _5396_ ;
wire _3709_ ;
wire _3882_ ;
wire _3462_ ;
wire _3042_ ;
wire _4667_ ;
wire _4247_ ;
wire _2733_ ;
wire _2313_ ;
wire \genblk1[1].u_ce.Vld_bF$buf4  ;
wire _3938_ ;
wire _3518_ ;
wire _3691_ ;
wire _3271_ ;
wire _4896_ ;
wire _4476_ ;
wire _4056_ ;
wire _915_ ;
wire _6202_ ;
wire _2962_ ;
wire _2542_ ;
wire _2122_ ;
wire _3747_ ;
wire _3327_ ;
wire _3080_ ;
wire _1813_ ;
wire _4285_ ;
wire _724_ ;
wire _304_ ;
wire _6011_ ;
wire _2771_ ;
wire _2351_ ;
wire _3976_ ;
wire _3556_ ;
wire _3136_ ;
wire _5702_ ;
wire \genblk1[3].u_ce.Vld_bF$buf0  ;
wire _1622_ ;
wire _1202_ ;
wire _4094_ ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _2827_ ;
wire _2407_ ;
wire _5299_ ;
wire _6240_ ;
wire _2580_ ;
wire _2160_ ;
wire _3785_ ;
wire _3365_ ;
wire _5931_ ;
wire _5511_ ;
wire _1851_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire _2636_ ;
wire _2216_ ;
wire _3594_ ;
wire _3174_ ;
wire _1907_ ;
wire _4799_ ;
wire _4379_ ;
wire _5740_ ;
wire _5320_ ;
wire _818_ ;
wire _78_ ;
wire _6105_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _2865_ ;
wire _2445_ ;
wire _2025_ ;
wire _1716_ ;
wire _4188_ ;
wire _627_ ;
wire _207_ ;
wire _6334_ ;
wire _380_ ;
wire _2674_ ;
wire _2254_ ;
wire clk_bF$buf30 ;
wire clk_bF$buf31 ;
wire clk_bF$buf32 ;
wire clk_bF$buf33 ;
wire clk_bF$buf34 ;
wire clk_bF$buf35 ;
wire clk_bF$buf36 ;
wire clk_bF$buf37 ;
wire [1:0] \genblk1[2].u_ce.Yin1  ;
wire clk_bF$buf38 ;
wire clk_bF$buf39 ;
wire _3879_ ;
wire _3459_ ;
wire _3039_ ;
wire _4820_ ;
wire _4400_ ;
wire _5605_ ;
wire [1:0] \genblk1[5].u_ce.Ain0  ;
wire _1945_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _6143_ ;
wire _2483_ ;
wire _2063_ ;
wire _3688_ ;
wire _3268_ ;
wire _5834_ ;
wire _5414_ ;
wire _1754_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _2959_ ;
wire _2539_ ;
wire _2119_ ;
wire _3900_ ;
wire _2292_ ;
wire _3497_ ;
wire _3077_ ;
wire _5643_ ;
wire _5223_ ;
wire _6008_ ;
wire _1983_ ;
wire _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _2768_ ;
wire _2348_ ;
wire \genblk1[5].u_ce.Ain12b_11_bF$buf0  ;
wire _6181_ ;
wire _4914_ ;
wire _1619_ ;
wire _5872_ ;
wire _5452_ ;
wire _5032_ ;
wire _6237_ ;
wire _1792_ ;
wire _1372_ ;
wire _283_ ;
wire _2997_ ;
wire _2577_ ;
wire _2157_ ;
wire _4723_ ;
wire _4303_ ;
wire _5928_ ;
wire _5508_ ;
wire _1848_ ;
wire _1428_ ;
wire _1008_ ;
wire _5681_ ;
wire _5261_ ;
wire _759_ ;
wire _339_ ;
wire \genblk1[2].u_ce.LoadCtl_0_bF$buf1  ;
wire _6046_ ;
wire _1181_ ;
wire _2386_ ;
wire _4952_ ;
wire _4532_ ;
wire _4112_ ;
wire _5737_ ;
wire _5317_ ;
wire _1657_ ;
wire _1237_ ;
wire _5490_ ;
wire _5070_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _3803_ ;
wire _6275_ ;
wire _2195_ ;
wire _4761_ ;
wire _4341_ ;
wire _5966_ ;
wire _5546_ ;
wire _5126_ ;
wire _40_ ;
wire _1886_ ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire _3612_ ;
wire _6084_ ;
wire _4817_ ;
wire _4990_ ;
wire _4570_ ;
wire _4150_ ;
wire _5775_ ;
wire _5355_ ;
wire _1695_ ;
wire _1275_ ;
wire _186_ ;
wire _3841_ ;
wire _3421_ ;
wire _3001_ ;
wire _4626_ ;
wire _4206_ ;
wire _5584_ ;
wire _5164_ ;
wire _1084_ ;
wire _3628__bF$buf0 ;
wire _3628__bF$buf1 ;
wire _3628__bF$buf2 ;
wire _3628__bF$buf3 ;
wire _3628__bF$buf4 ;
wire [1:0] \a[3]  ;
wire _2289_ ;
wire _3650_ ;
wire _3230_ ;
wire _4855_ ;
wire _4435_ ;
wire _4015_ ;
wire _2921_ ;
wire _2501_ ;
wire _5393_ ;
wire _3706_ ;
wire _6178_ ;
wire _2098_ ;
wire _4664_ ;
wire _4244_ ;
wire _5869_ ;
wire _5449_ ;
wire _5029_ ;
wire _1789_ ;
wire _1369_ ;
wire _2730_ ;
wire _2310_ ;
wire \genblk1[1].u_ce.Vld_bF$buf1  ;
wire _3935_ ;
wire _3515_ ;
wire [6:0] \genblk1[6].u_ce.LoadCtl  ;
wire _4893_ ;
wire _4473_ ;
wire _4053_ ;
wire _912_ ;
wire _5678_ ;
wire _5258_ ;
wire _1598_ ;
wire _1178_ ;
wire [1:0] \genblk1[0].u_ce.Y_  ;
wire _3744_ ;
wire _3324_ ;
wire _4949_ ;
wire _4529_ ;
wire _4109_ ;
wire _1810_ ;
wire _4282_ ;
wire _721_ ;
wire _301_ ;
wire _5487_ ;
wire _5067_ ;
wire _3973_ ;
wire _3553_ ;
wire _3133_ ;
wire _4758_ ;
wire _4338_ ;
wire _37_ ;
wire _4091_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _2824_ ;
wire _2404_ ;
wire _5296_ ;
wire _3609_ ;
wire _3782_ ;
wire _3362_ ;
wire _4987_ ;
wire _4567_ ;
wire _4147_ ;
wire _2633_ ;
wire _2213_ ;
wire _3838_ ;
wire _3418_ ;
wire _3591_ ;
wire _3171_ ;
wire _1904_ ;
wire _4796_ ;
wire _4376_ ;
wire _815_ ;
wire _75_ ;
wire _6102_ ;
wire _2862_ ;
wire _2442_ ;
wire _2022_ ;
wire _3647_ ;
wire _3227_ ;
wire _1713_ ;
wire _4185_ ;
wire _624_ ;
wire _204_ ;
wire _2918_ ;
wire \genblk1[6].u_ce.Vld  ;
wire _6331_ ;
wire _2671_ ;
wire _2251_ ;
wire _3876_ ;
wire _3456_ ;
wire _3036_ ;
wire \genblk1[3].u_ce.Ain12b_11_bF$buf3  ;
wire _5602_ ;
wire _1942_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _2727_ ;
wire _2307_ ;
wire _5199_ ;
wire _6140_ ;
wire _2480_ ;
wire _2060_ ;
wire _3685_ ;
wire _3265_ ;
wire _5831_ ;
wire _5411_ ;
wire _909_ ;
wire _1751_ ;
wire _1331_ ;
wire _662_ ;
wire _242_ ;
wire _2956_ ;
wire _2536_ ;
wire _2116_ ;
wire \genblk1[0].u_ce.LoadCtl_0_bF$buf4  ;
wire _3494_ ;
wire _3074_ ;
wire _1807_ ;
wire _4699_ ;
wire _4279_ ;
wire _5640_ ;
wire _5220_ ;
wire _718_ ;
wire _6005_ ;
wire _1980_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _2765_ ;
wire _2345_ ;
wire _4911_ ;
wire _1616_ ;
wire _4088_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _6234_ ;
wire _280_ ;
wire _2994_ ;
wire _2574_ ;
wire _2154_ ;
wire _3779_ ;
wire _3359_ ;
wire _4720_ ;
wire _4300_ ;
wire _5925_ ;
wire _5505_ ;
wire _1845_ ;
wire [1:0] \genblk1[5].u_ce.Xin1  ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire _6043_ ;
wire _2383_ ;
wire _3588_ ;
wire _3168_ ;
wire _5734_ ;
wire _5314_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _2859_ ;
wire _2439_ ;
wire _2019_ ;
wire _3800_ ;
wire _6272_ ;
wire _2192_ ;
wire _3397_ ;
wire _5963_ ;
wire _5543_ ;
wire _5123_ ;
wire _6328_ ;
wire _1883_ ;
wire _1463_ ;
wire _1043_ ;
wire _794_ ;
wire _374_ ;
wire _2668_ ;
wire _2248_ ;
wire _6081_ ;
wire _4814_ ;
wire _1939_ ;
wire _1519_ ;
wire _5772_ ;
wire _5352_ ;
wire _6137_ ;
wire _1692_ ;
wire _1272_ ;
wire _183_ ;
wire _2897_ ;
wire _2477_ ;
wire _2057_ ;
wire _4623_ ;
wire _4203_ ;
wire _5828_ ;
wire _5408_ ;
wire _1748_ ;
wire _1328_ ;
wire _5581_ ;
wire _5161_ ;
wire _659_ ;
wire _239_ ;
wire _1081_ ;
wire _2286_ ;
wire _4852_ ;
wire _4432_ ;
wire _4012_ ;
wire _5637_ ;
wire _5217_ ;
wire _1977_ ;
wire _1557_ ;
wire _1137_ ;
wire _5390_ ;
wire _888_ ;
wire _468_ ;
wire _3703_ ;
wire _6175_ ;
wire _4908_ ;
wire _2095_ ;
wire _4661_ ;
wire _4241_ ;
wire _5866_ ;
wire _5446_ ;
wire _5026_ ;
wire _1786_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _3932_ ;
wire _3512_ ;
wire _4717_ ;
wire _4890_ ;
wire _4470_ ;
wire _4050_ ;
wire _5675_ ;
wire _5255_ ;
wire _1595_ ;
wire _1175_ ;
wire _3741_ ;
wire _3321_ ;
wire _4946_ ;
wire _4526_ ;
wire _4106_ ;
wire _191__bF$buf0 ;
wire _191__bF$buf1 ;
wire _191__bF$buf2 ;
wire _191__bF$buf3 ;
wire _5484_ ;
wire _5064_ ;
wire _6269_ ;
wire _2189_ ;
wire _3970_ ;
wire _3550_ ;
wire _3130_ ;
wire _4755_ ;
wire _4335_ ;
wire _34_ ;
wire _2821_ ;
wire _2401_ ;
wire _5293_ ;
wire _3606_ ;
wire _6078_ ;
wire _4984_ ;
wire _4564_ ;
wire _4144_ ;
wire _5769_ ;
wire _5349_ ;
wire _1689_ ;
wire _1269_ ;
wire _2630_ ;
wire _2210_ ;
wire _3835_ ;
wire _3415_ ;
wire _1901_ ;
wire _4793_ ;
wire _4373_ ;
wire _812_ ;
wire _5998_ ;
wire _5578_ ;
wire _5158_ ;
wire _72_ ;
wire _1498_ ;
wire _1078_ ;
wire _3644_ ;
wire _3224_ ;
wire _4849_ ;
wire _4429_ ;
wire _4009_ ;
wire _1710_ ;
wire _4182_ ;
wire _621_ ;
wire _201_ ;
wire _2915_ ;
wire _5387_ ;
wire [1:0] \genblk1[1].u_ce.Yin0  ;
wire _3873_ ;
wire _3453_ ;
wire _3033_ ;
wire _4658_ ;
wire \genblk1[3].u_ce.Ain12b_11_bF$buf0  ;
wire _4238_ ;
wire _850_ ;
wire _430_ ;
wire _2724_ ;
wire _2304_ ;
wire _5196_ ;
wire _3929_ ;
wire _3509_ ;
wire _3682_ ;
wire _3262_ ;
wire _4887_ ;
wire _4467_ ;
wire _4047_ ;
wire _906_ ;
wire _2953_ ;
wire _2533_ ;
wire _2113_ ;
wire _3738_ ;
wire _3318_ ;
wire \genblk1[0].u_ce.LoadCtl_0_bF$buf1  ;
wire _3491_ ;
wire _3071_ ;
wire _1804_ ;
wire _4696_ ;
wire _4276_ ;
wire _715_ ;
wire _6002_ ;
wire _2762_ ;
wire _2342_ ;
wire _3967_ ;
wire _3547_ ;
wire _3127_ ;
wire _1613_ ;
wire _4085_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _2818_ ;
wire _6231_ ;
wire _2991_ ;
wire _2571_ ;
wire _2151_ ;
wire _3776_ ;
wire _3356_ ;
wire _5922_ ;
wire _5502_ ;
wire _1842_ ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire _333_ ;
wire _2627_ ;
wire _2207_ ;
wire _5099_ ;
wire _6040_ ;
wire _2380_ ;
wire _3585_ ;
wire _3165_ ;
wire _5731_ ;
wire _5311_ ;
wire _809_ ;
wire _69_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _2856_ ;
wire _2436_ ;
wire _2016_ ;
wire _3394_ ;
wire _1707_ ;
wire _4599_ ;
wire _4179_ ;
wire _5960_ ;
wire _5540_ ;
wire _5120_ ;
wire _618_ ;
wire _6325_ ;
wire _1880_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _2665_ ;
wire _2245_ ;
wire _4811_ ;
wire _1936_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire _6134_ ;
wire _180_ ;
wire _2894_ ;
wire _2474_ ;
wire _2054_ ;
wire _3679_ ;
wire _3259_ ;
wire _4620_ ;
wire _4200_ ;
wire _5825_ ;
wire _5405_ ;
wire _1745_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _2283_ ;
wire [6:0] \u_ot.LoadCtl  ;
wire _3488_ ;
wire _3068_ ;
wire _5634_ ;
wire _5214_ ;
wire _1974_ ;
wire _1554_ ;
wire _1134_ ;
wire \genblk1[5].u_ce.LoadCtl_0_bF$buf4  ;
wire _885_ ;
wire _465_ ;
wire _3717__bF$buf0 ;
wire _3717__bF$buf1 ;
wire _3717__bF$buf2 ;
wire _2759_ ;
wire _3717__bF$buf3 ;
wire _2339_ ;
wire _3717__bF$buf4 ;
wire _3717__bF$buf5 ;
wire \genblk1[4].u_ce.Vld_bF$buf3  ;
wire _3700_ ;
wire _6172_ ;
wire _4905_ ;
wire _2092_ ;
wire _3297_ ;
wire _5863_ ;
wire _5443_ ;
wire _5023_ ;
wire _6228_ ;
wire _1783_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _2988_ ;
wire _2568_ ;
wire _2148_ ;
wire _4714_ ;
wire _5919_ ;
wire _1839_ ;
wire _1419_ ;
wire _5672_ ;
wire _5252_ ;
wire _6037_ ;
wire _1592_ ;
wire _1172_ ;
wire _2797_ ;
wire _2377_ ;
wire _4943_ ;
wire _4523_ ;
wire _4103_ ;
wire _5728_ ;
wire _5308_ ;
wire _1648_ ;
wire _1228_ ;
wire _5481_ ;
wire _5061_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _6266_ ;
wire _2186_ ;
wire _4752_ ;
wire _4332_ ;
wire _5957_ ;
wire _5537_ ;
wire _5117_ ;
wire _31_ ;
wire _1877_ ;
wire _1457_ ;
wire _1037_ ;
wire _5290_ ;
wire _788_ ;
wire _368_ ;
wire _3603_ ;
wire _6075_ ;
wire _4808_ ;
wire _4981_ ;
wire _4561_ ;
wire _4141_ ;
wire _5766_ ;
wire _5346_ ;
wire \genblk1[1].u_ce.Ain12b_11_bF$buf3  ;
wire _1686_ ;
wire _1266_ ;
wire _597_ ;
wire _177_ ;
wire _3832_ ;
wire _3412_ ;
wire _4617_ ;
wire _4790_ ;
wire _4370_ ;
wire _5995_ ;
wire _5575_ ;
wire _5155_ ;
wire _1495_ ;
wire _1075_ ;
wire _3641_ ;
wire _3221_ ;
wire _4846_ ;
wire _4426_ ;
wire _4006_ ;
wire _2912_ ;
wire _5384_ ;
wire _6169_ ;
wire _2089_ ;
wire _3870_ ;
wire _3450_ ;
wire _3030_ ;
wire _4655_ ;
wire _4235_ ;
wire [1:0] \genblk1[3].u_ce.Ain1  ;
wire _2721_ ;
wire _2301_ ;
wire _5193_ ;
wire _3926_ ;
wire _3506_ ;
wire _4884_ ;
wire _4464_ ;
wire _4044_ ;
wire _903_ ;
wire _5669_ ;
wire _5249_ ;
wire _1589_ ;
wire _1169_ ;
wire _2950_ ;
wire _2530_ ;
wire _2110_ ;
wire _3735_ ;
wire _3315_ ;
wire _1801_ ;
wire _4693_ ;
wire _4273_ ;
wire _712_ ;
wire [1:0] \genblk1[1].u_ce.Y_  ;
wire _5898_ ;
wire _5478_ ;
wire _5058_ ;
wire _1398_ ;
wire _3964_ ;
wire _3544_ ;
wire _3124_ ;
wire [11:0] \genblk1[0].u_ce.Xin12b  ;
wire _4749_ ;
wire _4329_ ;
wire _28_ ;
wire _1610_ ;
wire _4082_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _2815_ ;
wire _5287_ ;
wire _3773_ ;
wire _3353_ ;
wire _4978_ ;
wire _4558_ ;
wire _4138_ ;
wire [1:0] \genblk1[4].u_ce.Xin0  ;
wire _750_ ;
wire _330_ ;
wire _2624_ ;
wire _2204_ ;
wire _5096_ ;
wire _3829_ ;
wire _3409_ ;
wire _3582_ ;
wire _3162_ ;
wire _4787_ ;
wire _4367_ ;
wire _806_ ;
wire _66_ ;
wire _2853_ ;
wire _2433_ ;
wire _2013_ ;
wire _3638_ ;
wire _3218_ ;
wire _3391_ ;
wire _1704_ ;
wire _4596_ ;
wire _4176_ ;
wire _615_ ;
wire _2909_ ;
wire _6322_ ;
wire _2662_ ;
wire _2242_ ;
wire _3867_ ;
wire _3447_ ;
wire _3027_ ;
wire _1933_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _2718_ ;
wire _6131_ ;
wire _2891_ ;
wire _2471_ ;
wire _2051_ ;
wire _3676_ ;
wire _3256_ ;
wire _5822_ ;
wire _5402_ ;
wire _1742_ ;
wire _1322_ ;
wire _653_ ;
wire _233_ ;
wire _2947_ ;
wire _2527_ ;
wire _2107_ ;
wire _2280_ ;
wire _3485_ ;
wire _3065_ ;
wire _5631_ ;
wire _5211_ ;
wire _709_ ;
wire _1971_ ;
wire _1551_ ;
wire _1131_ ;
wire \genblk1[5].u_ce.LoadCtl_0_bF$buf1  ;
wire _882_ ;
wire _462_ ;
wire _2756_ ;
wire _2336_ ;
wire \genblk1[4].u_ce.Vld_bF$buf0  ;
wire _4902_ ;
wire _3294_ ;
wire _1607_ ;
wire _4499_ ;
wire _4079_ ;
wire _5860_ ;
wire _5440_ ;
wire _5020_ ;
wire _938_ ;
wire _518_ ;
wire _6225_ ;
wire _1780_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _2985_ ;
wire _2565_ ;
wire _2145_ ;
wire _4711_ ;
wire _5916_ ;
wire _1836_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _6034_ ;
wire _2794_ ;
wire _2374_ ;
wire _3999_ ;
wire _3579_ ;
wire _3159_ ;
wire _4940_ ;
wire _4520_ ;
wire _4100_ ;
wire _5725_ ;
wire _5305_ ;
wire _1645_ ;
wire _1225_ ;
wire [1:0] \genblk1[6].u_ce.Yin1  ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire _6263_ ;
wire _2183_ ;
wire _3388_ ;
wire _5954_ ;
wire _5534_ ;
wire _5114_ ;
wire _6319_ ;
wire _1874_ ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _2659_ ;
wire _2239_ ;
wire _3600_ ;
wire _6072_ ;
wire _4805_ ;
wire [11:0] \genblk1[3].u_ce.Yin12b  ;
wire _3197_ ;
wire _5763_ ;
wire _5343_ ;
wire \genblk1[1].u_ce.Ain12b_11_bF$buf0  ;
wire _6128_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _2888_ ;
wire _2468_ ;
wire _2048_ ;
wire _4614_ ;
wire [11:0] \u_ot.Xin12b  ;
wire _5819_ ;
wire _1739_ ;
wire _1319_ ;
wire _5992_ ;
wire _5572_ ;
wire _5152_ ;
wire _1492_ ;
wire _1072_ ;
wire _2697_ ;
wire _2277_ ;
wire _4843_ ;
wire _4423_ ;
wire _4003_ ;
wire _5628_ ;
wire _5208_ ;
wire _1968_ ;
wire _1548_ ;
wire _1128_ ;
wire _5381_ ;
wire _879_ ;
wire _459_ ;
wire _6166_ ;
wire _2086_ ;
wire _4652_ ;
wire _4232_ ;
wire _5857_ ;
wire _5437_ ;
wire _5017_ ;
wire _1777_ ;
wire _1357_ ;
wire _5190_ ;
wire _688_ ;
wire _268_ ;
wire _3923_ ;
wire _3503_ ;
wire _4708_ ;
wire [11:0] \genblk1[5].u_ce.Yin12b  ;
wire _4881_ ;
wire _4461_ ;
wire _4041_ ;
wire _900_ ;
wire _5666_ ;
wire _5246_ ;
wire _1586_ ;
wire _1166_ ;
wire _497_ ;
wire _3732_ ;
wire _3312_ ;
wire _4937_ ;
wire _4517_ ;
wire \genblk1[6].u_ce.Ain12b_11_bF$buf1  ;
wire _4690_ ;
wire _4270_ ;
wire _5895_ ;
wire _5475_ ;
wire _5055_ ;
wire _1395_ ;
wire _3961_ ;
wire _3541_ ;
wire _3121_ ;
wire _4746_ ;
wire _4326_ ;
wire _25_ ;
wire _2812_ ;
wire _5284_ ;
wire _6069_ ;
wire \genblk1[3].u_ce.LoadCtl_0_bF$buf2  ;
wire _3770_ ;
wire _3350_ ;
wire _4975_ ;
wire _4555_ ;
wire _4135_ ;
wire _2621_ ;
wire _2201_ ;
wire _5093_ ;
wire _3826_ ;
wire _3406_ ;
wire _6298_ ;
wire _4784_ ;
wire _4364_ ;
wire _803_ ;
wire _5989_ ;
wire _5569_ ;
wire _5149_ ;
wire _63_ ;
wire _1489_ ;
wire _1069_ ;
wire _2850_ ;
wire _2430_ ;
wire _2010_ ;
wire _3635_ ;
wire _3215_ ;
wire \genblk1[5].u_ce.ISout  ;
wire _1701_ ;
wire _4593_ ;
wire _4173_ ;
wire _612_ ;
wire _2906_ ;
wire _5798_ ;
wire _5378_ ;
wire _1298_ ;
wire _3864_ ;
wire _3444_ ;
wire _3024_ ;
wire _4649_ ;
wire _4229_ ;
wire _1930_ ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _2715_ ;
wire _5187_ ;
wire _3673_ ;
wire _3253_ ;
wire _4878_ ;
wire _4458_ ;
wire _4038_ ;
wire _650_ ;
wire _230_ ;
wire _2944_ ;
wire _2524_ ;
wire _2104_ ;
wire _3729_ ;
wire _3309_ ;
wire _3482_ ;
wire _3062_ ;
wire _4687_ ;
wire _4267_ ;
wire _706_ ;
wire _2753_ ;
wire _2333_ ;
wire _3958_ ;
wire _3538_ ;
wire _3118_ ;
wire \genblk1[2].u_ce.Vld_bF$buf3  ;
wire _3291_ ;
wire _1604_ ;
wire _4496_ ;
wire _4076_ ;
wire _935_ ;
wire _515_ ;
wire _2809_ ;
wire _6222_ ;
wire _2982_ ;
wire _2562_ ;
wire _2142_ ;
wire _3767_ ;
wire _3347_ ;
wire _5913_ ;
wire _1833_ ;
wire _1413_ ;
wire _744_ ;
wire _324_ ;
wire _2618_ ;
wire _6031_ ;
wire _2791_ ;
wire _2371_ ;
wire _3996_ ;
wire _3576_ ;
wire _3156_ ;
wire _5722_ ;
wire _5302_ ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _2847_ ;
wire _2427_ ;
wire _2007_ ;
wire _6260_ ;
wire _2180_ ;
wire _3385_ ;
wire _5951_ ;
wire _5531_ ;
wire _5111_ ;
wire _609_ ;
wire \genblk1[4].u_ce.Vld  ;
wire _6316_ ;
wire _1871_ ;
wire _1451_ ;
wire _1031_ ;
wire _782_ ;
wire _362_ ;
wire _2656_ ;
wire _2236_ ;
wire _4802_ ;
wire _3194_ ;
wire _1927_ ;
wire _1507_ ;
wire _4399_ ;
wire _5760_ ;
wire _5340_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _6125_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _2885_ ;
wire _2465_ ;
wire _2045_ ;
wire _4611_ ;
wire _5816_ ;
wire _1736_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire _2694_ ;
wire _2274_ ;
wire _3899_ ;
wire _3479_ ;
wire _3059_ ;
wire _4840_ ;
wire _4420_ ;
wire _4000_ ;
wire _5625_ ;
wire _5205_ ;
wire _1965_ ;
wire _1545_ ;
wire \genblk1[4].u_ce.Ain12b_11_bF$buf4  ;
wire _1125_ ;
wire _876_ ;
wire _456_ ;
wire _6163_ ;
wire _2083_ ;
wire _3288_ ;
wire _5854_ ;
wire _5434_ ;
wire _5014_ ;
wire [1:0] \genblk1[2].u_ce.Ain0  ;
wire _6219_ ;
wire _1774_ ;
wire _1354_ ;
wire _685_ ;
wire _265_ ;
wire _2979_ ;
wire _2559_ ;
wire _2139_ ;
wire _3920_ ;
wire _3500_ ;
wire _4705_ ;
wire _3097_ ;
wire _5663_ ;
wire _5243_ ;
wire _6028_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _2788_ ;
wire _2368_ ;
wire _4934_ ;
wire _4514_ ;
wire _5719_ ;
wire _1639_ ;
wire _1219_ ;
wire _5892_ ;
wire _5472_ ;
wire _5052_ ;
wire _6257_ ;
wire _1392_ ;
wire _2597_ ;
wire _2177_ ;
wire \u_ot.ISout  ;
wire _4743_ ;
wire _4323_ ;
wire _5948_ ;
wire _5528_ ;
wire _5108_ ;
wire _22_ ;
wire [11:0] \genblk1[2].u_ce.Acalc  ;
wire _1868_ ;
wire _1448_ ;
wire _1028_ ;
wire _5281_ ;
wire _779_ ;
wire _359_ ;
wire _6066_ ;

CLKBUF1 CLKBUF1_insert336 (
    .A(clk),
    .Y(clk_hier0_bF$buf0)
);

CLKBUF1 CLKBUF1_insert335 (
    .A(clk),
    .Y(clk_hier0_bF$buf1)
);

CLKBUF1 CLKBUF1_insert334 (
    .A(clk),
    .Y(clk_hier0_bF$buf2)
);

CLKBUF1 CLKBUF1_insert333 (
    .A(clk),
    .Y(clk_hier0_bF$buf3)
);

CLKBUF1 CLKBUF1_insert332 (
    .A(clk),
    .Y(clk_hier0_bF$buf4)
);

CLKBUF1 CLKBUF1_insert331 (
    .A(clk),
    .Y(clk_hier0_bF$buf5)
);

CLKBUF1 CLKBUF1_insert330 (
    .A(clk),
    .Y(clk_hier0_bF$buf6)
);

CLKBUF1 CLKBUF1_insert329 (
    .A(clk),
    .Y(clk_hier0_bF$buf7)
);

BUFX2 BUFX2_insert328 (
    .A(\u_ot.ISout ),
    .Y(\u_ot.ISout_bF$buf0 )
);

BUFX2 BUFX2_insert327 (
    .A(\u_ot.ISout ),
    .Y(\u_ot.ISout_bF$buf1 )
);

BUFX2 BUFX2_insert326 (
    .A(\u_ot.ISout ),
    .Y(\u_ot.ISout_bF$buf2 )
);

BUFX2 BUFX2_insert325 (
    .A(\u_ot.ISout ),
    .Y(\u_ot.ISout_bF$buf3 )
);

BUFX2 BUFX2_insert324 (
    .A(\u_ot.ISout ),
    .Y(\u_ot.ISout_bF$buf4 )
);

BUFX2 BUFX2_insert323 (
    .A(\genblk1[4].u_ce.Vld ),
    .Y(\genblk1[4].u_ce.Vld_bF$buf0 )
);

BUFX2 BUFX2_insert322 (
    .A(\genblk1[4].u_ce.Vld ),
    .Y(\genblk1[4].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert321 (
    .A(\genblk1[4].u_ce.Vld ),
    .Y(\genblk1[4].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert320 (
    .A(\genblk1[4].u_ce.Vld ),
    .Y(\genblk1[4].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert319 (
    .A(\genblk1[4].u_ce.Vld ),
    .Y(\genblk1[4].u_ce.Vld_bF$buf4 )
);

BUFX2 BUFX2_insert318 (
    .A(\genblk1[4].u_ce.LoadCtl [0]),
    .Y(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert317 (
    .A(\genblk1[4].u_ce.LoadCtl [0]),
    .Y(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert316 (
    .A(\genblk1[4].u_ce.LoadCtl [0]),
    .Y(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert315 (
    .A(\genblk1[4].u_ce.LoadCtl [0]),
    .Y(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert314 (
    .A(\genblk1[4].u_ce.LoadCtl [0]),
    .Y(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 )
);

BUFX2 BUFX2_insert313 (
    .A(_2756_),
    .Y(_2756__bF$buf0)
);

BUFX2 BUFX2_insert312 (
    .A(_2756_),
    .Y(_2756__bF$buf1)
);

BUFX2 BUFX2_insert311 (
    .A(_2756_),
    .Y(_2756__bF$buf2)
);

BUFX2 BUFX2_insert310 (
    .A(_2756_),
    .Y(_2756__bF$buf3)
);

BUFX2 BUFX2_insert309 (
    .A(_2756_),
    .Y(_2756__bF$buf4)
);

BUFX2 BUFX2_insert308 (
    .A(\genblk1[0].u_ce.LoadCtl [0]),
    .Y(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert307 (
    .A(\genblk1[0].u_ce.LoadCtl [0]),
    .Y(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert306 (
    .A(\genblk1[0].u_ce.LoadCtl [0]),
    .Y(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert305 (
    .A(\genblk1[0].u_ce.LoadCtl [0]),
    .Y(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert304 (
    .A(\genblk1[0].u_ce.LoadCtl [0]),
    .Y(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 )
);

BUFX2 BUFX2_insert303 (
    .A(_2762_),
    .Y(_2762__bF$buf0)
);

BUFX2 BUFX2_insert302 (
    .A(_2762_),
    .Y(_2762__bF$buf1)
);

BUFX2 BUFX2_insert301 (
    .A(_2762_),
    .Y(_2762__bF$buf2)
);

BUFX2 BUFX2_insert300 (
    .A(_2762_),
    .Y(_2762__bF$buf3)
);

BUFX2 BUFX2_insert299 (
    .A(_2762_),
    .Y(_2762__bF$buf4)
);

BUFX2 BUFX2_insert298 (
    .A(\genblk1[4].u_ce.Ain12b [11]),
    .Y(\genblk1[4].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert297 (
    .A(\genblk1[4].u_ce.Ain12b [11]),
    .Y(\genblk1[4].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert296 (
    .A(\genblk1[4].u_ce.Ain12b [11]),
    .Y(\genblk1[4].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert295 (
    .A(\genblk1[4].u_ce.Ain12b [11]),
    .Y(\genblk1[4].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert294 (
    .A(\genblk1[4].u_ce.Ain12b [11]),
    .Y(\genblk1[4].u_ce.Ain12b_11_bF$buf4 )
);

BUFX2 BUFX2_insert293 (
    .A(_5270_),
    .Y(_5270__bF$buf0)
);

BUFX2 BUFX2_insert292 (
    .A(_5270_),
    .Y(_5270__bF$buf1)
);

BUFX2 BUFX2_insert291 (
    .A(_5270_),
    .Y(_5270__bF$buf2)
);

BUFX2 BUFX2_insert290 (
    .A(_5270_),
    .Y(_5270__bF$buf3)
);

BUFX2 BUFX2_insert289 (
    .A(\genblk1[0].u_ce.Ain12b [11]),
    .Y(\genblk1[0].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert288 (
    .A(\genblk1[0].u_ce.Ain12b [11]),
    .Y(\genblk1[0].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert287 (
    .A(\genblk1[0].u_ce.Ain12b [11]),
    .Y(\genblk1[0].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert286 (
    .A(\genblk1[0].u_ce.Ain12b [11]),
    .Y(\genblk1[0].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert285 (
    .A(\genblk1[0].u_ce.Ain12b [11]),
    .Y(\genblk1[0].u_ce.Ain12b_11_bF$buf4 )
);

BUFX2 BUFX2_insert284 (
    .A(_5276_),
    .Y(_5276__bF$buf0)
);

BUFX2 BUFX2_insert283 (
    .A(_5276_),
    .Y(_5276__bF$buf1)
);

BUFX2 BUFX2_insert282 (
    .A(_5276_),
    .Y(_5276__bF$buf2)
);

BUFX2 BUFX2_insert281 (
    .A(_5276_),
    .Y(_5276__bF$buf3)
);

BUFX2 BUFX2_insert280 (
    .A(_5276_),
    .Y(_5276__bF$buf4)
);

BUFX2 BUFX2_insert279 (
    .A(_2789_),
    .Y(_2789__bF$buf0)
);

BUFX2 BUFX2_insert278 (
    .A(_2789_),
    .Y(_2789__bF$buf1)
);

BUFX2 BUFX2_insert277 (
    .A(_2789_),
    .Y(_2789__bF$buf2)
);

BUFX2 BUFX2_insert276 (
    .A(_2789_),
    .Y(_2789__bF$buf3)
);

BUFX2 BUFX2_insert275 (
    .A(_5303_),
    .Y(_5303__bF$buf0)
);

BUFX2 BUFX2_insert274 (
    .A(_5303_),
    .Y(_5303__bF$buf1)
);

BUFX2 BUFX2_insert273 (
    .A(_5303_),
    .Y(_5303__bF$buf2)
);

BUFX2 BUFX2_insert272 (
    .A(_5303_),
    .Y(_5303__bF$buf3)
);

BUFX2 BUFX2_insert271 (
    .A(_2851_),
    .Y(_2851__bF$buf0)
);

BUFX2 BUFX2_insert270 (
    .A(_2851_),
    .Y(_2851__bF$buf1)
);

BUFX2 BUFX2_insert269 (
    .A(_2851_),
    .Y(_2851__bF$buf2)
);

BUFX2 BUFX2_insert268 (
    .A(_2851_),
    .Y(_2851__bF$buf3)
);

BUFX2 BUFX2_insert267 (
    .A(_2851_),
    .Y(_2851__bF$buf4)
);

BUFX2 BUFX2_insert266 (
    .A(_2851_),
    .Y(_2851__bF$buf5)
);

BUFX2 BUFX2_insert265 (
    .A(\genblk1[3].u_ce.LoadCtl [0]),
    .Y(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert264 (
    .A(\genblk1[3].u_ce.LoadCtl [0]),
    .Y(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert263 (
    .A(\genblk1[3].u_ce.LoadCtl [0]),
    .Y(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert262 (
    .A(\genblk1[3].u_ce.LoadCtl [0]),
    .Y(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert261 (
    .A(\genblk1[3].u_ce.LoadCtl [0]),
    .Y(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 )
);

BUFX2 BUFX2_insert260 (
    .A(\genblk1[2].u_ce.LoadCtl [0]),
    .Y(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert259 (
    .A(\genblk1[2].u_ce.LoadCtl [0]),
    .Y(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert258 (
    .A(\genblk1[2].u_ce.LoadCtl [0]),
    .Y(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert257 (
    .A(\genblk1[2].u_ce.LoadCtl [0]),
    .Y(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert256 (
    .A(\genblk1[2].u_ce.LoadCtl [0]),
    .Y(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 )
);

BUFX2 BUFX2_insert255 (
    .A(\genblk1[1].u_ce.Vld ),
    .Y(\genblk1[1].u_ce.Vld_bF$buf0 )
);

BUFX2 BUFX2_insert254 (
    .A(\genblk1[1].u_ce.Vld ),
    .Y(\genblk1[1].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert253 (
    .A(\genblk1[1].u_ce.Vld ),
    .Y(\genblk1[1].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert252 (
    .A(\genblk1[1].u_ce.Vld ),
    .Y(\genblk1[1].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert251 (
    .A(\genblk1[1].u_ce.Vld ),
    .Y(\genblk1[1].u_ce.Vld_bF$buf4 )
);

BUFX2 BUFX2_insert250 (
    .A(_4474_),
    .Y(_4474__bF$buf0)
);

BUFX2 BUFX2_insert249 (
    .A(_4474_),
    .Y(_4474__bF$buf1)
);

BUFX2 BUFX2_insert248 (
    .A(_4474_),
    .Y(_4474__bF$buf2)
);

BUFX2 BUFX2_insert247 (
    .A(_4474_),
    .Y(_4474__bF$buf3)
);

BUFX2 BUFX2_insert246 (
    .A(_4474_),
    .Y(_4474__bF$buf4)
);

BUFX2 BUFX2_insert245 (
    .A(_6047_),
    .Y(_6047__bF$buf0)
);

BUFX2 BUFX2_insert244 (
    .A(_6047_),
    .Y(_6047__bF$buf1)
);

BUFX2 BUFX2_insert243 (
    .A(_6047_),
    .Y(_6047__bF$buf2)
);

BUFX2 BUFX2_insert242 (
    .A(_6047_),
    .Y(_6047__bF$buf3)
);

BUFX2 BUFX2_insert241 (
    .A(_1890_),
    .Y(_1890__bF$buf0)
);

BUFX2 BUFX2_insert240 (
    .A(_1890_),
    .Y(_1890__bF$buf1)
);

BUFX2 BUFX2_insert239 (
    .A(_1890_),
    .Y(_1890__bF$buf2)
);

BUFX2 BUFX2_insert238 (
    .A(_1890_),
    .Y(_1890__bF$buf3)
);

BUFX2 BUFX2_insert237 (
    .A(_1890_),
    .Y(_1890__bF$buf4)
);

BUFX2 BUFX2_insert236 (
    .A(\genblk1[3].u_ce.Ain12b [11]),
    .Y(\genblk1[3].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert235 (
    .A(\genblk1[3].u_ce.Ain12b [11]),
    .Y(\genblk1[3].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert234 (
    .A(\genblk1[3].u_ce.Ain12b [11]),
    .Y(\genblk1[3].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert233 (
    .A(\genblk1[3].u_ce.Ain12b [11]),
    .Y(\genblk1[3].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert232 (
    .A(\genblk1[3].u_ce.Ain12b [11]),
    .Y(\genblk1[3].u_ce.Ain12b_11_bF$buf4 )
);

BUFX2 BUFX2_insert231 (
    .A(_4480_),
    .Y(_4480__bF$buf0)
);

BUFX2 BUFX2_insert230 (
    .A(_4480_),
    .Y(_4480__bF$buf1)
);

BUFX2 BUFX2_insert229 (
    .A(_4480_),
    .Y(_4480__bF$buf2)
);

BUFX2 BUFX2_insert228 (
    .A(_4480_),
    .Y(_4480__bF$buf3)
);

BUFX2 BUFX2_insert227 (
    .A(_4480_),
    .Y(_4480__bF$buf4)
);

BUFX2 BUFX2_insert226 (
    .A(\genblk1[2].u_ce.Ain12b [11]),
    .Y(\genblk1[2].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert225 (
    .A(\genblk1[2].u_ce.Ain12b [11]),
    .Y(\genblk1[2].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert224 (
    .A(\genblk1[2].u_ce.Ain12b [11]),
    .Y(\genblk1[2].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert223 (
    .A(\genblk1[2].u_ce.Ain12b [11]),
    .Y(\genblk1[2].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert222 (
    .A(\genblk1[2].u_ce.Ain12b [11]),
    .Y(\genblk1[2].u_ce.Ain12b_11_bF$buf4 )
);

BUFX2 BUFX2_insert221 (
    .A(_5365_),
    .Y(_5365__bF$buf0)
);

BUFX2 BUFX2_insert220 (
    .A(_5365_),
    .Y(_5365__bF$buf1)
);

BUFX2 BUFX2_insert219 (
    .A(_5365_),
    .Y(_5365__bF$buf2)
);

BUFX2 BUFX2_insert218 (
    .A(_5365_),
    .Y(_5365__bF$buf3)
);

BUFX2 BUFX2_insert217 (
    .A(_5365_),
    .Y(_5365__bF$buf4)
);

BUFX2 BUFX2_insert216 (
    .A(_5365_),
    .Y(_5365__bF$buf5)
);

BUFX2 BUFX2_insert215 (
    .A(_3622_),
    .Y(_3622__bF$buf0)
);

BUFX2 BUFX2_insert214 (
    .A(_3622_),
    .Y(_3622__bF$buf1)
);

BUFX2 BUFX2_insert213 (
    .A(_3622_),
    .Y(_3622__bF$buf2)
);

BUFX2 BUFX2_insert212 (
    .A(_3622_),
    .Y(_3622__bF$buf3)
);

BUFX2 BUFX2_insert211 (
    .A(_3622_),
    .Y(_3622__bF$buf4)
);

BUFX2 BUFX2_insert210 (
    .A(_1896_),
    .Y(_1896__bF$buf0)
);

BUFX2 BUFX2_insert209 (
    .A(_1896_),
    .Y(_1896__bF$buf1)
);

BUFX2 BUFX2_insert208 (
    .A(_1896_),
    .Y(_1896__bF$buf2)
);

BUFX2 BUFX2_insert207 (
    .A(_1896_),
    .Y(_1896__bF$buf3)
);

BUFX2 BUFX2_insert206 (
    .A(_1896_),
    .Y(_1896__bF$buf4)
);

BUFX2 BUFX2_insert205 (
    .A(_158_),
    .Y(_158__bF$buf0)
);

BUFX2 BUFX2_insert204 (
    .A(_158_),
    .Y(_158__bF$buf1)
);

BUFX2 BUFX2_insert203 (
    .A(_158_),
    .Y(_158__bF$buf2)
);

BUFX2 BUFX2_insert202 (
    .A(_158_),
    .Y(_158__bF$buf3)
);

BUFX2 BUFX2_insert201 (
    .A(_158_),
    .Y(_158__bF$buf4)
);

BUFX2 BUFX2_insert200 (
    .A(\genblk1[3].u_ce.Vld ),
    .Y(\genblk1[3].u_ce.Vld_bF$buf0 )
);

BUFX2 BUFX2_insert199 (
    .A(\genblk1[3].u_ce.Vld ),
    .Y(\genblk1[3].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert198 (
    .A(\genblk1[3].u_ce.Vld ),
    .Y(\genblk1[3].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert197 (
    .A(\genblk1[3].u_ce.Vld ),
    .Y(\genblk1[3].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert196 (
    .A(\genblk1[3].u_ce.Vld ),
    .Y(\genblk1[3].u_ce.Vld_bF$buf4 )
);

BUFX2 BUFX2_insert195 (
    .A(_4507_),
    .Y(_4507__bF$buf0)
);

BUFX2 BUFX2_insert194 (
    .A(_4507_),
    .Y(_4507__bF$buf1)
);

BUFX2 BUFX2_insert193 (
    .A(_4507_),
    .Y(_4507__bF$buf2)
);

BUFX2 BUFX2_insert192 (
    .A(_4507_),
    .Y(_4507__bF$buf3)
);

BUFX2 BUFX2_insert191 (
    .A(_164_),
    .Y(_164__bF$buf0)
);

BUFX2 BUFX2_insert190 (
    .A(_164_),
    .Y(_164__bF$buf1)
);

BUFX2 BUFX2_insert189 (
    .A(_164_),
    .Y(_164__bF$buf2)
);

BUFX2 BUFX2_insert188 (
    .A(_164_),
    .Y(_164__bF$buf3)
);

BUFX2 BUFX2_insert187 (
    .A(_164_),
    .Y(_164__bF$buf4)
);

BUFX2 BUFX2_insert186 (
    .A(_1024_),
    .Y(_1024__bF$buf0)
);

BUFX2 BUFX2_insert185 (
    .A(_1024_),
    .Y(_1024__bF$buf1)
);

BUFX2 BUFX2_insert184 (
    .A(_1024_),
    .Y(_1024__bF$buf2)
);

BUFX2 BUFX2_insert183 (
    .A(_1024_),
    .Y(_1024__bF$buf3)
);

BUFX2 BUFX2_insert182 (
    .A(_1024_),
    .Y(_1024__bF$buf4)
);

BUFX2 BUFX2_insert181 (
    .A(_1923_),
    .Y(_1923__bF$buf0)
);

BUFX2 BUFX2_insert180 (
    .A(_1923_),
    .Y(_1923__bF$buf1)
);

BUFX2 BUFX2_insert179 (
    .A(_1923_),
    .Y(_1923__bF$buf2)
);

BUFX2 BUFX2_insert178 (
    .A(_1923_),
    .Y(_1923__bF$buf3)
);

BUFX2 BUFX2_insert177 (
    .A(_3628_),
    .Y(_3628__bF$buf0)
);

BUFX2 BUFX2_insert176 (
    .A(_3628_),
    .Y(_3628__bF$buf1)
);

BUFX2 BUFX2_insert175 (
    .A(_3628_),
    .Y(_3628__bF$buf2)
);

BUFX2 BUFX2_insert174 (
    .A(_3628_),
    .Y(_3628__bF$buf3)
);

BUFX2 BUFX2_insert173 (
    .A(_3628_),
    .Y(_3628__bF$buf4)
);

BUFX2 BUFX2_insert172 (
    .A(\genblk1[6].u_ce.LoadCtl [0]),
    .Y(\genblk1[6].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert171 (
    .A(\genblk1[6].u_ce.LoadCtl [0]),
    .Y(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert170 (
    .A(\genblk1[6].u_ce.LoadCtl [0]),
    .Y(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert169 (
    .A(\genblk1[6].u_ce.LoadCtl [0]),
    .Y(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert168 (
    .A(_1030_),
    .Y(_1030__bF$buf0)
);

BUFX2 BUFX2_insert167 (
    .A(_1030_),
    .Y(_1030__bF$buf1)
);

BUFX2 BUFX2_insert166 (
    .A(_1030_),
    .Y(_1030__bF$buf2)
);

BUFX2 BUFX2_insert165 (
    .A(_1030_),
    .Y(_1030__bF$buf3)
);

BUFX2 BUFX2_insert164 (
    .A(_1030_),
    .Y(_1030__bF$buf4)
);

BUFX2 BUFX2_insert163 (
    .A(\genblk1[5].u_ce.LoadCtl [0]),
    .Y(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert162 (
    .A(\genblk1[5].u_ce.LoadCtl [0]),
    .Y(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert161 (
    .A(\genblk1[5].u_ce.LoadCtl [0]),
    .Y(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert160 (
    .A(\genblk1[5].u_ce.LoadCtl [0]),
    .Y(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert159 (
    .A(\genblk1[5].u_ce.LoadCtl [0]),
    .Y(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 )
);

BUFX2 BUFX2_insert158 (
    .A(\genblk1[5].u_ce.Vld ),
    .Y(\genblk1[5].u_ce.Vld_bF$buf0 )
);

BUFX2 BUFX2_insert157 (
    .A(\genblk1[5].u_ce.Vld ),
    .Y(\genblk1[5].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert156 (
    .A(\genblk1[5].u_ce.Vld ),
    .Y(\genblk1[5].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert155 (
    .A(\genblk1[5].u_ce.Vld ),
    .Y(\genblk1[5].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert154 (
    .A(_6133_),
    .Y(_6133__bF$buf0)
);

BUFX2 BUFX2_insert153 (
    .A(_6133_),
    .Y(_6133__bF$buf1)
);

BUFX2 BUFX2_insert152 (
    .A(_6133_),
    .Y(_6133__bF$buf2)
);

BUFX2 BUFX2_insert151 (
    .A(_6133_),
    .Y(_6133__bF$buf3)
);

BUFX2 BUFX2_insert150 (
    .A(\genblk1[1].u_ce.LoadCtl [0]),
    .Y(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 )
);

BUFX2 BUFX2_insert149 (
    .A(\genblk1[1].u_ce.LoadCtl [0]),
    .Y(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 )
);

BUFX2 BUFX2_insert148 (
    .A(\genblk1[1].u_ce.LoadCtl [0]),
    .Y(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 )
);

BUFX2 BUFX2_insert147 (
    .A(\genblk1[1].u_ce.LoadCtl [0]),
    .Y(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 )
);

BUFX2 BUFX2_insert146 (
    .A(\genblk1[1].u_ce.LoadCtl [0]),
    .Y(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 )
);

BUFX2 BUFX2_insert145 (
    .A(\genblk1[0].u_ce.Vld ),
    .Y(\genblk1[0].u_ce.Vld_bF$buf0 )
);

BUFX2 BUFX2_insert144 (
    .A(\genblk1[0].u_ce.Vld ),
    .Y(\genblk1[0].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert143 (
    .A(\genblk1[0].u_ce.Vld ),
    .Y(\genblk1[0].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert142 (
    .A(\genblk1[0].u_ce.Vld ),
    .Y(\genblk1[0].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert141 (
    .A(\genblk1[0].u_ce.Vld ),
    .Y(\genblk1[0].u_ce.Vld_bF$buf4 )
);

BUFX2 BUFX2_insert140 (
    .A(selXY),
    .Y(selXY_bF$buf0)
);

BUFX2 BUFX2_insert139 (
    .A(selXY),
    .Y(selXY_bF$buf1)
);

BUFX2 BUFX2_insert138 (
    .A(selXY),
    .Y(selXY_bF$buf2)
);

BUFX2 BUFX2_insert137 (
    .A(selXY),
    .Y(selXY_bF$buf3)
);

BUFX2 BUFX2_insert136 (
    .A(\genblk1[6].u_ce.Ain12b [11]),
    .Y(\genblk1[6].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert135 (
    .A(\genblk1[6].u_ce.Ain12b [11]),
    .Y(\genblk1[6].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert134 (
    .A(\genblk1[6].u_ce.Ain12b [11]),
    .Y(\genblk1[6].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert133 (
    .A(\genblk1[6].u_ce.Ain12b [11]),
    .Y(\genblk1[6].u_ce.Ain12b_11_bF$buf3 )
);

CLKBUF1 CLKBUF1_insert132 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert131 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert130 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert129 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert128 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert127 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert126 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert125 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert124 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf8)
);

CLKBUF1 CLKBUF1_insert123 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf9)
);

CLKBUF1 CLKBUF1_insert122 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf10)
);

CLKBUF1 CLKBUF1_insert121 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf11)
);

CLKBUF1 CLKBUF1_insert120 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf12)
);

CLKBUF1 CLKBUF1_insert119 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf13)
);

CLKBUF1 CLKBUF1_insert118 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf14)
);

CLKBUF1 CLKBUF1_insert117 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf15)
);

CLKBUF1 CLKBUF1_insert116 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf16)
);

CLKBUF1 CLKBUF1_insert115 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf17)
);

CLKBUF1 CLKBUF1_insert114 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf18)
);

CLKBUF1 CLKBUF1_insert113 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf19)
);

CLKBUF1 CLKBUF1_insert112 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf20)
);

CLKBUF1 CLKBUF1_insert111 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf21)
);

CLKBUF1 CLKBUF1_insert110 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf22)
);

CLKBUF1 CLKBUF1_insert109 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf23)
);

CLKBUF1 CLKBUF1_insert108 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf24)
);

CLKBUF1 CLKBUF1_insert107 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf25)
);

CLKBUF1 CLKBUF1_insert106 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf26)
);

CLKBUF1 CLKBUF1_insert105 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf27)
);

CLKBUF1 CLKBUF1_insert104 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf28)
);

CLKBUF1 CLKBUF1_insert103 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf29)
);

CLKBUF1 CLKBUF1_insert102 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf30)
);

CLKBUF1 CLKBUF1_insert101 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf31)
);

CLKBUF1 CLKBUF1_insert100 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf32)
);

CLKBUF1 CLKBUF1_insert99 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf33)
);

CLKBUF1 CLKBUF1_insert98 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf34)
);

CLKBUF1 CLKBUF1_insert97 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf35)
);

CLKBUF1 CLKBUF1_insert96 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf36)
);

CLKBUF1 CLKBUF1_insert95 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf37)
);

CLKBUF1 CLKBUF1_insert94 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf38)
);

CLKBUF1 CLKBUF1_insert93 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf39)
);

CLKBUF1 CLKBUF1_insert92 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf40)
);

CLKBUF1 CLKBUF1_insert91 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf41)
);

CLKBUF1 CLKBUF1_insert90 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf42)
);

CLKBUF1 CLKBUF1_insert89 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf43)
);

CLKBUF1 CLKBUF1_insert88 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf44)
);

CLKBUF1 CLKBUF1_insert87 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf45)
);

CLKBUF1 CLKBUF1_insert86 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf46)
);

CLKBUF1 CLKBUF1_insert85 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf47)
);

CLKBUF1 CLKBUF1_insert84 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf48)
);

CLKBUF1 CLKBUF1_insert83 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf49)
);

CLKBUF1 CLKBUF1_insert82 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf50)
);

CLKBUF1 CLKBUF1_insert81 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf51)
);

CLKBUF1 CLKBUF1_insert80 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf52)
);

CLKBUF1 CLKBUF1_insert79 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf53)
);

CLKBUF1 CLKBUF1_insert78 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf54)
);

CLKBUF1 CLKBUF1_insert77 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf55)
);

CLKBUF1 CLKBUF1_insert76 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf56)
);

CLKBUF1 CLKBUF1_insert75 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf57)
);

CLKBUF1 CLKBUF1_insert74 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf58)
);

CLKBUF1 CLKBUF1_insert73 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf59)
);

CLKBUF1 CLKBUF1_insert72 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf60)
);

CLKBUF1 CLKBUF1_insert71 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf61)
);

CLKBUF1 CLKBUF1_insert70 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf62)
);

CLKBUF1 CLKBUF1_insert69 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf63)
);

CLKBUF1 CLKBUF1_insert68 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf64)
);

CLKBUF1 CLKBUF1_insert67 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf65)
);

CLKBUF1 CLKBUF1_insert66 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf66)
);

CLKBUF1 CLKBUF1_insert65 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf67)
);

CLKBUF1 CLKBUF1_insert64 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf68)
);

CLKBUF1 CLKBUF1_insert63 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf69)
);

CLKBUF1 CLKBUF1_insert62 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf70)
);

CLKBUF1 CLKBUF1_insert61 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf71)
);

CLKBUF1 CLKBUF1_insert60 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf72)
);

CLKBUF1 CLKBUF1_insert59 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf73)
);

CLKBUF1 CLKBUF1_insert58 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf74)
);

CLKBUF1 CLKBUF1_insert57 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf75)
);

BUFX2 BUFX2_insert56 (
    .A(_4569_),
    .Y(_4569__bF$buf0)
);

BUFX2 BUFX2_insert55 (
    .A(_4569_),
    .Y(_4569__bF$buf1)
);

BUFX2 BUFX2_insert54 (
    .A(_4569_),
    .Y(_4569__bF$buf2)
);

BUFX2 BUFX2_insert53 (
    .A(_4569_),
    .Y(_4569__bF$buf3)
);

BUFX2 BUFX2_insert52 (
    .A(_4569_),
    .Y(_4569__bF$buf4)
);

BUFX2 BUFX2_insert51 (
    .A(_4569_),
    .Y(_4569__bF$buf5)
);

BUFX2 BUFX2_insert50 (
    .A(\genblk1[5].u_ce.Ain12b [11]),
    .Y(\genblk1[5].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert49 (
    .A(\genblk1[5].u_ce.Ain12b [11]),
    .Y(\genblk1[5].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert48 (
    .A(\genblk1[5].u_ce.Ain12b [11]),
    .Y(\genblk1[5].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert47 (
    .A(\genblk1[5].u_ce.Ain12b [11]),
    .Y(\genblk1[5].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert46 (
    .A(\genblk1[5].u_ce.Ain12b [11]),
    .Y(\genblk1[5].u_ce.Ain12b_11_bF$buf4 )
);

BUFX2 BUFX2_insert45 (
    .A(_1985_),
    .Y(_1985__bF$buf0)
);

BUFX2 BUFX2_insert44 (
    .A(_1985_),
    .Y(_1985__bF$buf1)
);

BUFX2 BUFX2_insert43 (
    .A(_1985_),
    .Y(_1985__bF$buf2)
);

BUFX2 BUFX2_insert42 (
    .A(_1985_),
    .Y(_1985__bF$buf3)
);

BUFX2 BUFX2_insert41 (
    .A(_1985_),
    .Y(_1985__bF$buf4)
);

BUFX2 BUFX2_insert40 (
    .A(_1985_),
    .Y(_1985__bF$buf5)
);

BUFX2 BUFX2_insert39 (
    .A(_191_),
    .Y(_191__bF$buf0)
);

BUFX2 BUFX2_insert38 (
    .A(_191_),
    .Y(_191__bF$buf1)
);

BUFX2 BUFX2_insert37 (
    .A(_191_),
    .Y(_191__bF$buf2)
);

BUFX2 BUFX2_insert36 (
    .A(_191_),
    .Y(_191__bF$buf3)
);

BUFX2 BUFX2_insert35 (
    .A(_3655_),
    .Y(_3655__bF$buf0)
);

BUFX2 BUFX2_insert34 (
    .A(_3655_),
    .Y(_3655__bF$buf1)
);

BUFX2 BUFX2_insert33 (
    .A(_3655_),
    .Y(_3655__bF$buf2)
);

BUFX2 BUFX2_insert32 (
    .A(_3655_),
    .Y(_3655__bF$buf3)
);

BUFX2 BUFX2_insert31 (
    .A(\genblk1[2].u_ce.Vld ),
    .Y(\genblk1[2].u_ce.Vld_bF$buf0 )
);

BUFX2 BUFX2_insert30 (
    .A(\genblk1[2].u_ce.Vld ),
    .Y(\genblk1[2].u_ce.Vld_bF$buf1 )
);

BUFX2 BUFX2_insert29 (
    .A(\genblk1[2].u_ce.Vld ),
    .Y(\genblk1[2].u_ce.Vld_bF$buf2 )
);

BUFX2 BUFX2_insert28 (
    .A(\genblk1[2].u_ce.Vld ),
    .Y(\genblk1[2].u_ce.Vld_bF$buf3 )
);

BUFX2 BUFX2_insert27 (
    .A(\genblk1[2].u_ce.Vld ),
    .Y(\genblk1[2].u_ce.Vld_bF$buf4 )
);

BUFX2 BUFX2_insert26 (
    .A(_253_),
    .Y(_253__bF$buf0)
);

BUFX2 BUFX2_insert25 (
    .A(_253_),
    .Y(_253__bF$buf1)
);

BUFX2 BUFX2_insert24 (
    .A(_253_),
    .Y(_253__bF$buf2)
);

BUFX2 BUFX2_insert23 (
    .A(_253_),
    .Y(_253__bF$buf3)
);

BUFX2 BUFX2_insert22 (
    .A(_253_),
    .Y(_253__bF$buf4)
);

BUFX2 BUFX2_insert21 (
    .A(_253_),
    .Y(_253__bF$buf5)
);

BUFX2 BUFX2_insert20 (
    .A(\genblk1[1].u_ce.Ain12b [11]),
    .Y(\genblk1[1].u_ce.Ain12b_11_bF$buf0 )
);

BUFX2 BUFX2_insert19 (
    .A(\genblk1[1].u_ce.Ain12b [11]),
    .Y(\genblk1[1].u_ce.Ain12b_11_bF$buf1 )
);

BUFX2 BUFX2_insert18 (
    .A(\genblk1[1].u_ce.Ain12b [11]),
    .Y(\genblk1[1].u_ce.Ain12b_11_bF$buf2 )
);

BUFX2 BUFX2_insert17 (
    .A(\genblk1[1].u_ce.Ain12b [11]),
    .Y(\genblk1[1].u_ce.Ain12b_11_bF$buf3 )
);

BUFX2 BUFX2_insert16 (
    .A(\genblk1[1].u_ce.Ain12b [11]),
    .Y(\genblk1[1].u_ce.Ain12b_11_bF$buf4 )
);

BUFX2 BUFX2_insert15 (
    .A(_3717_),
    .Y(_3717__bF$buf0)
);

BUFX2 BUFX2_insert14 (
    .A(_3717_),
    .Y(_3717__bF$buf1)
);

BUFX2 BUFX2_insert13 (
    .A(_3717_),
    .Y(_3717__bF$buf2)
);

BUFX2 BUFX2_insert12 (
    .A(_3717_),
    .Y(_3717__bF$buf3)
);

BUFX2 BUFX2_insert11 (
    .A(_3717_),
    .Y(_3717__bF$buf4)
);

BUFX2 BUFX2_insert10 (
    .A(_3717_),
    .Y(_3717__bF$buf5)
);

BUFX2 BUFX2_insert9 (
    .A(_1057_),
    .Y(_1057__bF$buf0)
);

BUFX2 BUFX2_insert8 (
    .A(_1057_),
    .Y(_1057__bF$buf1)
);

BUFX2 BUFX2_insert7 (
    .A(_1057_),
    .Y(_1057__bF$buf2)
);

BUFX2 BUFX2_insert6 (
    .A(_1057_),
    .Y(_1057__bF$buf3)
);

BUFX2 BUFX2_insert5 (
    .A(_1119_),
    .Y(_1119__bF$buf0)
);

BUFX2 BUFX2_insert4 (
    .A(_1119_),
    .Y(_1119__bF$buf1)
);

BUFX2 BUFX2_insert3 (
    .A(_1119_),
    .Y(_1119__bF$buf2)
);

BUFX2 BUFX2_insert2 (
    .A(_1119_),
    .Y(_1119__bF$buf3)
);

BUFX2 BUFX2_insert1 (
    .A(_1119_),
    .Y(_1119__bF$buf4)
);

BUFX2 BUFX2_insert0 (
    .A(_1119_),
    .Y(_1119__bF$buf5)
);

NOR2X1 _10000_ (
    .A(_3425_),
    .B(_3419_),
    .Y(_3426_)
);

NAND2X1 _10001_ (
    .A(_3425_),
    .B(_3419_),
    .Y(_3427_)
);

NAND2X1 _10002_ (
    .A(\genblk1[3].u_ce.Vld_bF$buf4 ),
    .B(_3427_),
    .Y(_3428_)
);

OAI21X1 _10003_ (
    .A(_3426_),
    .B(_3428_),
    .C(_3418_),
    .Y(_2633_)
);

AOI21X1 _10004_ (
    .A(_3419_),
    .B(_3421_),
    .C(_3422_),
    .Y(_3429_)
);

INVX1 _10005_ (
    .A(\genblk1[3].u_ce.Ain12b [10]),
    .Y(_3430_)
);

NAND2X1 _10006_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf4 ),
    .B(_3430_),
    .Y(_3431_)
);

NAND2X1 _10007_ (
    .A(\genblk1[3].u_ce.Ain12b [10]),
    .B(_2851__bF$buf5),
    .Y(_3432_)
);

NAND2X1 _10008_ (
    .A(_3431_),
    .B(_3432_),
    .Y(_3433_)
);

AND2X2 _10009_ (
    .A(_3429_),
    .B(_3433_),
    .Y(_3434_)
);

OAI21X1 _10010_ (
    .A(_3433_),
    .B(_3429_),
    .C(\genblk1[3].u_ce.Vld_bF$buf3 ),
    .Y(_3435_)
);

OAI22X1 _10011_ (
    .A(_2691_),
    .B(\genblk1[3].u_ce.Vld_bF$buf2 ),
    .C(_3435_),
    .D(_3434_),
    .Y(_2634_)
);

NAND2X1 _10012_ (
    .A(\genblk1[3].u_ce.Acalc [11]),
    .B(_2756__bF$buf4),
    .Y(_3436_)
);

OAI21X1 _10013_ (
    .A(_3433_),
    .B(_3429_),
    .C(_3432_),
    .Y(_3437_)
);

OAI21X1 _10014_ (
    .A(_2756__bF$buf3),
    .B(_3437_),
    .C(_3436_),
    .Y(_2635_)
);

INVX1 _10015_ (
    .A(_2690_),
    .Y(_3438_)
);

NAND3X1 _10016_ (
    .A(_2743_),
    .B(\genblk1[3].u_ce.LoadCtl [5]),
    .C(_2701_),
    .Y(_3439_)
);

NOR2X1 _10017_ (
    .A(_3438_),
    .B(_3439_),
    .Y(_3440_)
);

NAND2X1 _10018_ (
    .A(\genblk1[2].u_ce.X_ [0]),
    .B(_3440_),
    .Y(_3441_)
);

OAI21X1 _10019_ (
    .A(_2885_),
    .B(_3440_),
    .C(_3441_),
    .Y(_2636_)
);

NAND2X1 _10020_ (
    .A(\genblk1[2].u_ce.X_ [1]),
    .B(_3440_),
    .Y(_3442_)
);

OAI21X1 _10021_ (
    .A(_2910_),
    .B(_3440_),
    .C(_3442_),
    .Y(_2637_)
);

INVX1 _10022_ (
    .A(\genblk1[2].u_ce.X_ [0]),
    .Y(_3443_)
);

NAND3X1 _10023_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(_2690_),
    .C(_2701_),
    .Y(_3444_)
);

NAND2X1 _10024_ (
    .A(\genblk1[3].u_ce.Xin12b [8]),
    .B(_3444_),
    .Y(_3445_)
);

OAI21X1 _10025_ (
    .A(_3443_),
    .B(_3444_),
    .C(_3445_),
    .Y(_2638_)
);

INVX1 _10026_ (
    .A(\genblk1[2].u_ce.X_ [1]),
    .Y(_3446_)
);

NAND2X1 _10027_ (
    .A(\genblk1[3].u_ce.Xin12b [9]),
    .B(_3444_),
    .Y(_3447_)
);

OAI21X1 _10028_ (
    .A(_3446_),
    .B(_3444_),
    .C(_3447_),
    .Y(_2639_)
);

NAND2X1 _10029_ (
    .A(_2701_),
    .B(_2697_),
    .Y(_3448_)
);

OAI21X1 _10030_ (
    .A(_2702_),
    .B(_2710_),
    .C(\genblk1[3].u_ce.Xin12b [6]),
    .Y(_3449_)
);

OAI21X1 _10031_ (
    .A(_3443_),
    .B(_3448_),
    .C(_3449_),
    .Y(_2640_)
);

OAI21X1 _10032_ (
    .A(_2702_),
    .B(_2710_),
    .C(\genblk1[3].u_ce.Xin12b [7]),
    .Y(_3450_)
);

OAI21X1 _10033_ (
    .A(_3446_),
    .B(_3448_),
    .C(_3450_),
    .Y(_2641_)
);

NOR2X1 _10034_ (
    .A(_2694_),
    .B(_2702_),
    .Y(_3451_)
);

NAND2X1 _10035_ (
    .A(\genblk1[2].u_ce.X_ [0]),
    .B(_3451_),
    .Y(_3452_)
);

OAI21X1 _10036_ (
    .A(_2795_),
    .B(_3451_),
    .C(_3452_),
    .Y(_2642_)
);

NAND2X1 _10037_ (
    .A(\genblk1[2].u_ce.X_ [1]),
    .B(_3451_),
    .Y(_3453_)
);

OAI21X1 _10038_ (
    .A(_2803_),
    .B(_3451_),
    .C(_3453_),
    .Y(_2643_)
);

OAI21X1 _10039_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_2703_),
    .C(\genblk1[3].u_ce.Xin1 [0]),
    .Y(_3454_)
);

OAI21X1 _10040_ (
    .A(_3443_),
    .B(_2732_),
    .C(_3454_),
    .Y(_2644_)
);

OAI21X1 _10041_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_2703_),
    .C(\genblk1[3].u_ce.Xin1 [1]),
    .Y(_3455_)
);

OAI21X1 _10042_ (
    .A(_3446_),
    .B(_2732_),
    .C(_3455_),
    .Y(_2645_)
);

NAND2X1 _10043_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[2].u_ce.X_ [0]),
    .Y(_3456_)
);

OAI21X1 _10044_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_2818_),
    .C(_3456_),
    .Y(_2646_)
);

NAND2X1 _10045_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[2].u_ce.X_ [1]),
    .Y(_3457_)
);

OAI21X1 _10046_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_2798_),
    .C(_3457_),
    .Y(_2647_)
);

NAND2X1 _10047_ (
    .A(\genblk1[2].u_ce.Y_ [0]),
    .B(_3440_),
    .Y(_3458_)
);

OAI21X1 _10048_ (
    .A(_3018_),
    .B(_3440_),
    .C(_3458_),
    .Y(_2648_)
);

NAND2X1 _10049_ (
    .A(\genblk1[2].u_ce.Y_ [1]),
    .B(_3440_),
    .Y(_3459_)
);

OAI21X1 _10050_ (
    .A(_3042_),
    .B(_3440_),
    .C(_3459_),
    .Y(_2649_)
);

INVX1 _10051_ (
    .A(\genblk1[2].u_ce.Y_ [0]),
    .Y(_3460_)
);

NAND2X1 _10052_ (
    .A(\genblk1[3].u_ce.Yin12b [8]),
    .B(_3444_),
    .Y(_3461_)
);

OAI21X1 _10053_ (
    .A(_3460_),
    .B(_3444_),
    .C(_3461_),
    .Y(_2650_)
);

INVX1 _10054_ (
    .A(\genblk1[2].u_ce.Y_ [1]),
    .Y(_3462_)
);

NAND2X1 _10055_ (
    .A(\genblk1[3].u_ce.Yin12b [9]),
    .B(_3444_),
    .Y(_3463_)
);

OAI21X1 _10056_ (
    .A(_3462_),
    .B(_3444_),
    .C(_3463_),
    .Y(_2651_)
);

OAI21X1 _10057_ (
    .A(_2702_),
    .B(_2710_),
    .C(\genblk1[3].u_ce.Yin12b [6]),
    .Y(_2670_)
);

OAI21X1 _10058_ (
    .A(_3460_),
    .B(_3448_),
    .C(_2670_),
    .Y(_2652_)
);

OAI21X1 _10059_ (
    .A(_2702_),
    .B(_2710_),
    .C(\genblk1[3].u_ce.Yin12b [7]),
    .Y(_2671_)
);

OAI21X1 _10060_ (
    .A(_3462_),
    .B(_3448_),
    .C(_2671_),
    .Y(_2653_)
);

NAND2X1 _10061_ (
    .A(\genblk1[2].u_ce.Y_ [0]),
    .B(_3451_),
    .Y(_2672_)
);

OAI21X1 _10062_ (
    .A(_2883_),
    .B(_3451_),
    .C(_2672_),
    .Y(_2654_)
);

NAND2X1 _10063_ (
    .A(\genblk1[2].u_ce.Y_ [1]),
    .B(_3451_),
    .Y(_2673_)
);

OAI21X1 _10064_ (
    .A(_2908_),
    .B(_3451_),
    .C(_2673_),
    .Y(_2655_)
);

OAI21X1 _10065_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_2703_),
    .C(\genblk1[3].u_ce.Yin1 [0]),
    .Y(_2674_)
);

OAI21X1 _10066_ (
    .A(_3460_),
    .B(_2732_),
    .C(_2674_),
    .Y(_2656_)
);

OAI21X1 _10067_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_2703_),
    .C(\genblk1[3].u_ce.Yin1 [1]),
    .Y(_2675_)
);

OAI21X1 _10068_ (
    .A(_3462_),
    .B(_2732_),
    .C(_2675_),
    .Y(_2657_)
);

NAND2X1 _10069_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[2].u_ce.Y_ [0]),
    .Y(_2676_)
);

OAI21X1 _10070_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_3055_),
    .C(_2676_),
    .Y(_2658_)
);

NAND2X1 _10071_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[2].u_ce.Y_ [1]),
    .Y(_2677_)
);

OAI21X1 _10072_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_2840_),
    .C(_2677_),
    .Y(_2659_)
);

NAND2X1 _10073_ (
    .A(\a[3] [0]),
    .B(_3440_),
    .Y(_2678_)
);

OAI21X1 _10074_ (
    .A(_3430_),
    .B(_3440_),
    .C(_2678_),
    .Y(_2660_)
);

NAND2X1 _10075_ (
    .A(\a[3] [1]),
    .B(_3440_),
    .Y(_2679_)
);

OAI21X1 _10076_ (
    .A(_2851__bF$buf4),
    .B(_3440_),
    .C(_2679_),
    .Y(_2661_)
);

INVX1 _10077_ (
    .A(\a[3] [0]),
    .Y(_2680_)
);

NAND2X1 _10078_ (
    .A(\genblk1[3].u_ce.Ain12b [8]),
    .B(_3444_),
    .Y(_2681_)
);

OAI21X1 _10079_ (
    .A(_2680_),
    .B(_3444_),
    .C(_2681_),
    .Y(_2662_)
);

INVX1 _10080_ (
    .A(\a[3] [1]),
    .Y(_2682_)
);

NAND2X1 _10081_ (
    .A(\genblk1[3].u_ce.Ain12b [9]),
    .B(_3444_),
    .Y(_2683_)
);

OAI21X1 _10082_ (
    .A(_2682_),
    .B(_3444_),
    .C(_2683_),
    .Y(_2663_)
);

OAI21X1 _10083_ (
    .A(_2702_),
    .B(_2710_),
    .C(\genblk1[3].u_ce.Ain12b [6]),
    .Y(_2684_)
);

OAI21X1 _10084_ (
    .A(_2680_),
    .B(_3448_),
    .C(_2684_),
    .Y(_2664_)
);

OAI21X1 _10085_ (
    .A(_2702_),
    .B(_2710_),
    .C(\genblk1[3].u_ce.Ain12b [7]),
    .Y(_2685_)
);

OAI21X1 _10086_ (
    .A(_2682_),
    .B(_3448_),
    .C(_2685_),
    .Y(_2665_)
);

NAND2X1 _10087_ (
    .A(\a[3] [0]),
    .B(_3451_),
    .Y(_2686_)
);

OAI21X1 _10088_ (
    .A(_3354_),
    .B(_3451_),
    .C(_2686_),
    .Y(_2666_)
);

NAND2X1 _10089_ (
    .A(\a[3] [1]),
    .B(_3451_),
    .Y(_2687_)
);

OAI21X1 _10090_ (
    .A(_3368_),
    .B(_3451_),
    .C(_2687_),
    .Y(_2667_)
);

OAI21X1 _10091_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_2703_),
    .C(\genblk1[3].u_ce.Ain1 [0]),
    .Y(_2688_)
);

OAI21X1 _10092_ (
    .A(_2680_),
    .B(_2732_),
    .C(_2688_),
    .Y(_2668_)
);

OAI21X1 _10093_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_2703_),
    .C(\genblk1[3].u_ce.Ain1 [1]),
    .Y(_2689_)
);

OAI21X1 _10094_ (
    .A(_2682_),
    .B(_2732_),
    .C(_2689_),
    .Y(_2669_)
);

DFFPOSX1 _10095_ (
    .CLK(clk_bF$buf75),
    .D(_2598_),
    .Q(\genblk1[3].u_ce.Ain0 [0])
);

DFFPOSX1 _10096_ (
    .CLK(clk_bF$buf74),
    .D(_2599_),
    .Q(\genblk1[3].u_ce.Ain0 [1])
);

DFFPOSX1 _10097_ (
    .CLK(clk_bF$buf73),
    .D(_2600_),
    .Q(\genblk1[3].u_ce.Ycalc [2])
);

DFFPOSX1 _10098_ (
    .CLK(clk_bF$buf72),
    .D(_2601_),
    .Q(\genblk1[3].u_ce.Ycalc [3])
);

DFFPOSX1 _10099_ (
    .CLK(clk_bF$buf71),
    .D(_2602_),
    .Q(\genblk1[3].u_ce.Ycalc [4])
);

DFFPOSX1 _10100_ (
    .CLK(clk_bF$buf70),
    .D(_2603_),
    .Q(\genblk1[3].u_ce.Ycalc [5])
);

DFFPOSX1 _10101_ (
    .CLK(clk_bF$buf69),
    .D(_2604_),
    .Q(\genblk1[3].u_ce.Ycalc [6])
);

DFFPOSX1 _10102_ (
    .CLK(clk_bF$buf68),
    .D(_2605_),
    .Q(\genblk1[3].u_ce.Ycalc [7])
);

DFFPOSX1 _10103_ (
    .CLK(clk_bF$buf67),
    .D(_2606_),
    .Q(\genblk1[3].u_ce.Ycalc [8])
);

DFFPOSX1 _10104_ (
    .CLK(clk_bF$buf66),
    .D(_2607_),
    .Q(\genblk1[3].u_ce.Ycalc [9])
);

DFFPOSX1 _10105_ (
    .CLK(clk_bF$buf65),
    .D(_2608_),
    .Q(\genblk1[3].u_ce.Ycalc [10])
);

DFFPOSX1 _10106_ (
    .CLK(clk_bF$buf64),
    .D(_2609_),
    .Q(\genblk1[3].u_ce.Ycalc [11])
);

DFFPOSX1 _10107_ (
    .CLK(clk_bF$buf63),
    .D(_2610_),
    .Q(\genblk1[3].u_ce.Ycalc [0])
);

DFFPOSX1 _10108_ (
    .CLK(clk_bF$buf62),
    .D(_2611_),
    .Q(\genblk1[3].u_ce.Ycalc [1])
);

DFFPOSX1 _10109_ (
    .CLK(clk_bF$buf61),
    .D(_2612_),
    .Q(\genblk1[3].u_ce.Xcalc [0])
);

DFFPOSX1 _10110_ (
    .CLK(clk_bF$buf60),
    .D(_2613_),
    .Q(\genblk1[3].u_ce.Xcalc [1])
);

DFFPOSX1 _10111_ (
    .CLK(clk_bF$buf59),
    .D(_2614_),
    .Q(\genblk1[3].u_ce.Xcalc [2])
);

DFFPOSX1 _10112_ (
    .CLK(clk_bF$buf58),
    .D(_2615_),
    .Q(\genblk1[3].u_ce.Xcalc [3])
);

DFFPOSX1 _10113_ (
    .CLK(clk_bF$buf57),
    .D(_2616_),
    .Q(\genblk1[3].u_ce.Xcalc [4])
);

DFFPOSX1 _10114_ (
    .CLK(clk_bF$buf56),
    .D(_2617_),
    .Q(\genblk1[3].u_ce.Xcalc [5])
);

DFFPOSX1 _10115_ (
    .CLK(clk_bF$buf55),
    .D(_2618_),
    .Q(\genblk1[3].u_ce.Xcalc [6])
);

DFFPOSX1 _10116_ (
    .CLK(clk_bF$buf54),
    .D(_2619_),
    .Q(\genblk1[3].u_ce.Xcalc [7])
);

DFFPOSX1 _10117_ (
    .CLK(clk_bF$buf53),
    .D(_2620_),
    .Q(\genblk1[3].u_ce.Xcalc [8])
);

DFFPOSX1 _10118_ (
    .CLK(clk_bF$buf52),
    .D(_2621_),
    .Q(\genblk1[3].u_ce.Xcalc [9])
);

DFFPOSX1 _10119_ (
    .CLK(clk_bF$buf51),
    .D(_2622_),
    .Q(\genblk1[3].u_ce.Xcalc [10])
);

DFFPOSX1 _10120_ (
    .CLK(clk_bF$buf50),
    .D(_2623_),
    .Q(\genblk1[3].u_ce.Xcalc [11])
);

DFFPOSX1 _10121_ (
    .CLK(clk_bF$buf49),
    .D(_2624_),
    .Q(\genblk1[3].u_ce.Acalc [0])
);

DFFPOSX1 _10122_ (
    .CLK(clk_bF$buf48),
    .D(_2625_),
    .Q(\genblk1[3].u_ce.Acalc [1])
);

DFFPOSX1 _10123_ (
    .CLK(clk_bF$buf47),
    .D(_2626_),
    .Q(\genblk1[3].u_ce.Acalc [2])
);

DFFPOSX1 _10124_ (
    .CLK(clk_bF$buf46),
    .D(_2627_),
    .Q(\genblk1[3].u_ce.Acalc [3])
);

DFFPOSX1 _10125_ (
    .CLK(clk_bF$buf45),
    .D(_2628_),
    .Q(\genblk1[3].u_ce.Acalc [4])
);

DFFPOSX1 _10126_ (
    .CLK(clk_bF$buf44),
    .D(_2629_),
    .Q(\genblk1[3].u_ce.Acalc [5])
);

DFFPOSX1 _10127_ (
    .CLK(clk_bF$buf43),
    .D(_2630_),
    .Q(\genblk1[3].u_ce.Acalc [6])
);

DFFPOSX1 _10128_ (
    .CLK(clk_bF$buf42),
    .D(_2631_),
    .Q(\genblk1[3].u_ce.Acalc [7])
);

DFFPOSX1 _10129_ (
    .CLK(clk_bF$buf41),
    .D(_2632_),
    .Q(\genblk1[3].u_ce.Acalc [8])
);

DFFPOSX1 _10130_ (
    .CLK(clk_bF$buf40),
    .D(_2633_),
    .Q(\genblk1[3].u_ce.Acalc [9])
);

DFFPOSX1 _10131_ (
    .CLK(clk_bF$buf39),
    .D(_2634_),
    .Q(\genblk1[3].u_ce.Acalc [10])
);

DFFPOSX1 _10132_ (
    .CLK(clk_bF$buf38),
    .D(_2635_),
    .Q(\genblk1[3].u_ce.Acalc [11])
);

DFFPOSX1 _10133_ (
    .CLK(clk_bF$buf37),
    .D(_2636_),
    .Q(\genblk1[3].u_ce.Xin12b [10])
);

DFFPOSX1 _10134_ (
    .CLK(clk_bF$buf36),
    .D(_2637_),
    .Q(\genblk1[3].u_ce.Xin12b [11])
);

DFFPOSX1 _10135_ (
    .CLK(clk_bF$buf35),
    .D(_2638_),
    .Q(\genblk1[3].u_ce.Xin12b [8])
);

DFFPOSX1 _10136_ (
    .CLK(clk_bF$buf34),
    .D(_2639_),
    .Q(\genblk1[3].u_ce.Xin12b [9])
);

DFFPOSX1 _10137_ (
    .CLK(clk_bF$buf33),
    .D(_2640_),
    .Q(\genblk1[3].u_ce.Xin12b [6])
);

DFFPOSX1 _10138_ (
    .CLK(clk_bF$buf32),
    .D(_2641_),
    .Q(\genblk1[3].u_ce.Xin12b [7])
);

DFFPOSX1 _10139_ (
    .CLK(clk_bF$buf31),
    .D(_2642_),
    .Q(\genblk1[3].u_ce.Xin12b [4])
);

DFFPOSX1 _10140_ (
    .CLK(clk_bF$buf30),
    .D(_2643_),
    .Q(\genblk1[3].u_ce.Xin12b [5])
);

DFFPOSX1 _10141_ (
    .CLK(clk_bF$buf29),
    .D(_2644_),
    .Q(\genblk1[3].u_ce.Xin1 [0])
);

DFFPOSX1 _10142_ (
    .CLK(clk_bF$buf28),
    .D(_2645_),
    .Q(\genblk1[3].u_ce.Xin1 [1])
);

DFFPOSX1 _10143_ (
    .CLK(clk_bF$buf27),
    .D(_2646_),
    .Q(\genblk1[3].u_ce.Xin0 [0])
);

DFFPOSX1 _10144_ (
    .CLK(clk_bF$buf26),
    .D(_2647_),
    .Q(\genblk1[3].u_ce.Xin0 [1])
);

DFFPOSX1 _10145_ (
    .CLK(clk_bF$buf25),
    .D(_2648_),
    .Q(\genblk1[3].u_ce.Yin12b [10])
);

DFFPOSX1 _10146_ (
    .CLK(clk_bF$buf24),
    .D(_2649_),
    .Q(\genblk1[3].u_ce.Yin12b [11])
);

DFFPOSX1 _10147_ (
    .CLK(clk_bF$buf23),
    .D(_2650_),
    .Q(\genblk1[3].u_ce.Yin12b [8])
);

DFFPOSX1 _10148_ (
    .CLK(clk_bF$buf22),
    .D(_2651_),
    .Q(\genblk1[3].u_ce.Yin12b [9])
);

DFFPOSX1 _10149_ (
    .CLK(clk_bF$buf21),
    .D(_2652_),
    .Q(\genblk1[3].u_ce.Yin12b [6])
);

DFFPOSX1 _10150_ (
    .CLK(clk_bF$buf20),
    .D(_2653_),
    .Q(\genblk1[3].u_ce.Yin12b [7])
);

DFFPOSX1 _10151_ (
    .CLK(clk_bF$buf19),
    .D(_2654_),
    .Q(\genblk1[3].u_ce.Yin12b [4])
);

DFFPOSX1 _10152_ (
    .CLK(clk_bF$buf18),
    .D(_2655_),
    .Q(\genblk1[3].u_ce.Yin12b [5])
);

DFFPOSX1 _10153_ (
    .CLK(clk_bF$buf17),
    .D(_2656_),
    .Q(\genblk1[3].u_ce.Yin1 [0])
);

DFFPOSX1 _10154_ (
    .CLK(clk_bF$buf16),
    .D(_2657_),
    .Q(\genblk1[3].u_ce.Yin1 [1])
);

DFFPOSX1 _10155_ (
    .CLK(clk_bF$buf15),
    .D(_2658_),
    .Q(\genblk1[3].u_ce.Yin0 [0])
);

DFFPOSX1 _10156_ (
    .CLK(clk_bF$buf14),
    .D(_2659_),
    .Q(\genblk1[3].u_ce.Yin0 [1])
);

DFFPOSX1 _10157_ (
    .CLK(clk_bF$buf13),
    .D(_2660_),
    .Q(\genblk1[3].u_ce.Ain12b [10])
);

DFFPOSX1 _10158_ (
    .CLK(clk_bF$buf12),
    .D(_2661_),
    .Q(\genblk1[3].u_ce.Ain12b [11])
);

DFFPOSX1 _10159_ (
    .CLK(clk_bF$buf11),
    .D(_2662_),
    .Q(\genblk1[3].u_ce.Ain12b [8])
);

DFFPOSX1 _10160_ (
    .CLK(clk_bF$buf10),
    .D(_2663_),
    .Q(\genblk1[3].u_ce.Ain12b [9])
);

DFFPOSX1 _10161_ (
    .CLK(clk_bF$buf9),
    .D(_2664_),
    .Q(\genblk1[3].u_ce.Ain12b [6])
);

DFFPOSX1 _10162_ (
    .CLK(clk_bF$buf8),
    .D(_2665_),
    .Q(\genblk1[3].u_ce.Ain12b [7])
);

DFFPOSX1 _10163_ (
    .CLK(clk_bF$buf7),
    .D(_2666_),
    .Q(\genblk1[3].u_ce.Ain12b [4])
);

DFFPOSX1 _10164_ (
    .CLK(clk_bF$buf6),
    .D(_2667_),
    .Q(\genblk1[3].u_ce.Ain12b [5])
);

DFFPOSX1 _10165_ (
    .CLK(clk_bF$buf5),
    .D(_2668_),
    .Q(\genblk1[3].u_ce.Ain1 [0])
);

DFFPOSX1 _10166_ (
    .CLK(clk_bF$buf4),
    .D(_2669_),
    .Q(\genblk1[3].u_ce.Ain1 [1])
);

DFFPOSX1 _10167_ (
    .CLK(clk_bF$buf3),
    .D(\genblk1[2].u_ce.ISout ),
    .Q(\genblk1[3].u_ce.ISpipe [0])
);

DFFPOSX1 _10168_ (
    .CLK(clk_bF$buf2),
    .D(\genblk1[3].u_ce.ISpipe [0]),
    .Q(\genblk1[3].u_ce.ISpipe [1])
);

DFFPOSX1 _10169_ (
    .CLK(clk_bF$buf1),
    .D(\genblk1[3].u_ce.ISpipe [1]),
    .Q(\genblk1[3].u_ce.ISpipe [2])
);

DFFPOSX1 _10170_ (
    .CLK(clk_bF$buf0),
    .D(\genblk1[3].u_ce.ISpipe [2]),
    .Q(\genblk1[3].u_ce.ISpipe [3])
);

DFFPOSX1 _10171_ (
    .CLK(clk_bF$buf75),
    .D(\genblk1[3].u_ce.ISpipe [3]),
    .Q(\genblk1[3].u_ce.ISpipe [4])
);

DFFPOSX1 _10172_ (
    .CLK(clk_bF$buf74),
    .D(\genblk1[3].u_ce.ISpipe [4]),
    .Q(\genblk1[3].u_ce.ISpipe [5])
);

DFFPOSX1 _10173_ (
    .CLK(clk_bF$buf73),
    .D(\genblk1[3].u_ce.ISpipe [5]),
    .Q(\genblk1[3].u_ce.ISout )
);

DFFPOSX1 _10174_ (
    .CLK(clk_bF$buf72),
    .D(\genblk1[2].u_ce.Vld_bF$buf4 ),
    .Q(\genblk1[3].u_ce.LoadCtl [0])
);

DFFPOSX1 _10175_ (
    .CLK(clk_bF$buf71),
    .D(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 ),
    .Q(\genblk1[3].u_ce.LoadCtl [1])
);

DFFPOSX1 _10176_ (
    .CLK(clk_bF$buf70),
    .D(\genblk1[3].u_ce.LoadCtl [1]),
    .Q(\genblk1[3].u_ce.LoadCtl [2])
);

DFFPOSX1 _10177_ (
    .CLK(clk_bF$buf69),
    .D(\genblk1[3].u_ce.LoadCtl [2]),
    .Q(\genblk1[3].u_ce.LoadCtl [3])
);

DFFPOSX1 _10178_ (
    .CLK(clk_bF$buf68),
    .D(\genblk1[3].u_ce.LoadCtl [3]),
    .Q(\genblk1[3].u_ce.LoadCtl [4])
);

DFFPOSX1 _10179_ (
    .CLK(clk_bF$buf67),
    .D(\genblk1[3].u_ce.LoadCtl [4]),
    .Q(\genblk1[3].u_ce.LoadCtl [5])
);

DFFPOSX1 _10180_ (
    .CLK(clk_bF$buf66),
    .D(\genblk1[3].u_ce.LoadCtl [5]),
    .Q(\genblk1[3].u_ce.Vld )
);

NOR2X1 _10181_ (
    .A(\genblk1[4].u_ce.LoadCtl [3]),
    .B(\genblk1[4].u_ce.LoadCtl [2]),
    .Y(_3556_)
);

INVX1 _10182_ (
    .A(\genblk1[4].u_ce.Acalc [10]),
    .Y(_3557_)
);

NAND2X1 _10183_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(\genblk1[4].u_ce.Acalc [8]),
    .Y(_3558_)
);

OAI21X1 _10184_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(_3557_),
    .C(_3558_),
    .Y(_3559_)
);

INVX2 _10185_ (
    .A(\genblk1[4].u_ce.LoadCtl [2]),
    .Y(_3560_)
);

INVX1 _10186_ (
    .A(\genblk1[4].u_ce.Acalc [4]),
    .Y(_3561_)
);

INVX1 _10187_ (
    .A(\genblk1[4].u_ce.LoadCtl [3]),
    .Y(_3562_)
);

NOR2X1 _10188_ (
    .A(\genblk1[4].u_ce.LoadCtl [2]),
    .B(_3562_),
    .Y(_3563_)
);

NAND2X1 _10189_ (
    .A(\genblk1[4].u_ce.Acalc [6]),
    .B(_3563_),
    .Y(_3564_)
);

OAI21X1 _10190_ (
    .A(_3560_),
    .B(_3561_),
    .C(_3564_),
    .Y(_3565_)
);

AOI21X1 _10191_ (
    .A(_3556_),
    .B(_3559_),
    .C(_3565_),
    .Y(_3566_)
);

NOR2X1 _10192_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[4].u_ce.LoadCtl [1]),
    .Y(_3567_)
);

INVX4 _10193_ (
    .A(_3567_),
    .Y(_3568_)
);

INVX2 _10194_ (
    .A(\genblk1[4].u_ce.LoadCtl [1]),
    .Y(_3569_)
);

NOR2X1 _10195_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_3569_),
    .Y(_3570_)
);

AOI22X1 _10196_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[4].u_ce.Acalc [0]),
    .C(_3570_),
    .D(\genblk1[4].u_ce.Acalc [2]),
    .Y(_3571_)
);

OAI21X1 _10197_ (
    .A(_3568_),
    .B(_3566_),
    .C(_3571_),
    .Y(\a[5] [0])
);

INVX1 _10198_ (
    .A(\genblk1[4].u_ce.Acalc [11]),
    .Y(_3572_)
);

NAND2X1 _10199_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(\genblk1[4].u_ce.Acalc [9]),
    .Y(_3573_)
);

OAI21X1 _10200_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(_3572_),
    .C(_3573_),
    .Y(_3574_)
);

INVX1 _10201_ (
    .A(\genblk1[4].u_ce.Acalc [7]),
    .Y(_3575_)
);

INVX4 _10202_ (
    .A(_3563_),
    .Y(_3576_)
);

NAND2X1 _10203_ (
    .A(\genblk1[4].u_ce.LoadCtl [2]),
    .B(\genblk1[4].u_ce.Acalc [5]),
    .Y(_3577_)
);

OAI21X1 _10204_ (
    .A(_3575_),
    .B(_3576_),
    .C(_3577_),
    .Y(_3578_)
);

AOI21X1 _10205_ (
    .A(_3556_),
    .B(_3574_),
    .C(_3578_),
    .Y(_3579_)
);

AOI22X1 _10206_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[4].u_ce.Acalc [1]),
    .C(_3570_),
    .D(\genblk1[4].u_ce.Acalc [3]),
    .Y(_3580_)
);

OAI21X1 _10207_ (
    .A(_3568_),
    .B(_3579_),
    .C(_3580_),
    .Y(\a[5] [1])
);

INVX1 _10208_ (
    .A(\genblk1[4].u_ce.Ycalc [10]),
    .Y(_3581_)
);

NAND2X1 _10209_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(\genblk1[4].u_ce.Ycalc [8]),
    .Y(_3582_)
);

OAI21X1 _10210_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(_3581_),
    .C(_3582_),
    .Y(_3583_)
);

INVX1 _10211_ (
    .A(\genblk1[4].u_ce.Ycalc [6]),
    .Y(_3584_)
);

INVX1 _10212_ (
    .A(\genblk1[4].u_ce.Ycalc [4]),
    .Y(_3585_)
);

OAI22X1 _10213_ (
    .A(_3560_),
    .B(_3585_),
    .C(_3584_),
    .D(_3576_),
    .Y(_3586_)
);

AOI21X1 _10214_ (
    .A(_3556_),
    .B(_3583_),
    .C(_3586_),
    .Y(_3587_)
);

AOI22X1 _10215_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[4].u_ce.Ycalc [0]),
    .C(_3570_),
    .D(\genblk1[4].u_ce.Ycalc [2]),
    .Y(_3588_)
);

OAI21X1 _10216_ (
    .A(_3568_),
    .B(_3587_),
    .C(_3588_),
    .Y(\genblk1[4].u_ce.Y_ [0])
);

INVX1 _10217_ (
    .A(\genblk1[4].u_ce.Ycalc [11]),
    .Y(_3589_)
);

NAND2X1 _10218_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(\genblk1[4].u_ce.Ycalc [9]),
    .Y(_3590_)
);

OAI21X1 _10219_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(_3589_),
    .C(_3590_),
    .Y(_3591_)
);

INVX1 _10220_ (
    .A(\genblk1[4].u_ce.Ycalc [7]),
    .Y(_3592_)
);

INVX1 _10221_ (
    .A(\genblk1[4].u_ce.Ycalc [5]),
    .Y(_3593_)
);

OAI22X1 _10222_ (
    .A(_3560_),
    .B(_3593_),
    .C(_3592_),
    .D(_3576_),
    .Y(_3594_)
);

AOI21X1 _10223_ (
    .A(_3556_),
    .B(_3591_),
    .C(_3594_),
    .Y(_3595_)
);

AOI22X1 _10224_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[4].u_ce.Ycalc [1]),
    .C(_3570_),
    .D(\genblk1[4].u_ce.Ycalc [3]),
    .Y(_3596_)
);

OAI21X1 _10225_ (
    .A(_3568_),
    .B(_3595_),
    .C(_3596_),
    .Y(\genblk1[4].u_ce.Y_ [1])
);

INVX1 _10226_ (
    .A(\genblk1[4].u_ce.Xcalc [2]),
    .Y(_3597_)
);

INVX2 _10227_ (
    .A(_3570_),
    .Y(_3598_)
);

INVX1 _10228_ (
    .A(\genblk1[4].u_ce.Xcalc [4]),
    .Y(_3599_)
);

INVX1 _10229_ (
    .A(\genblk1[4].u_ce.Xcalc [6]),
    .Y(_3600_)
);

NOR2X1 _10230_ (
    .A(_3562_),
    .B(_3600_),
    .Y(_3601_)
);

INVX1 _10231_ (
    .A(\genblk1[4].u_ce.Xcalc [8]),
    .Y(_3602_)
);

NAND2X1 _10232_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(_3602_),
    .Y(_3603_)
);

OAI21X1 _10233_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(\genblk1[4].u_ce.Xcalc [10]),
    .C(_3603_),
    .Y(_3604_)
);

NOR2X1 _10234_ (
    .A(\genblk1[4].u_ce.LoadCtl [3]),
    .B(_3604_),
    .Y(_3605_)
);

OAI21X1 _10235_ (
    .A(_3601_),
    .B(_3605_),
    .C(_3560_),
    .Y(_3606_)
);

OAI21X1 _10236_ (
    .A(_3560_),
    .B(_3599_),
    .C(_3606_),
    .Y(_3607_)
);

AOI22X1 _10237_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[4].u_ce.Xcalc [0]),
    .C(_3607_),
    .D(_3567_),
    .Y(_3608_)
);

OAI21X1 _10238_ (
    .A(_3597_),
    .B(_3598_),
    .C(_3608_),
    .Y(\genblk1[4].u_ce.X_ [0])
);

INVX1 _10239_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .Y(_3609_)
);

INVX1 _10240_ (
    .A(\genblk1[4].u_ce.Xcalc [9]),
    .Y(_3610_)
);

NAND2X1 _10241_ (
    .A(\genblk1[4].u_ce.Xcalc [11]),
    .B(_3609_),
    .Y(_3611_)
);

OAI21X1 _10242_ (
    .A(_3609_),
    .B(_3610_),
    .C(_3611_),
    .Y(_3612_)
);

INVX1 _10243_ (
    .A(\genblk1[4].u_ce.Xcalc [7]),
    .Y(_3613_)
);

INVX1 _10244_ (
    .A(\genblk1[4].u_ce.Xcalc [5]),
    .Y(_3614_)
);

OAI22X1 _10245_ (
    .A(_3560_),
    .B(_3614_),
    .C(_3613_),
    .D(_3576_),
    .Y(_3615_)
);

AOI21X1 _10246_ (
    .A(_3556_),
    .B(_3612_),
    .C(_3615_),
    .Y(_3616_)
);

AOI22X1 _10247_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[4].u_ce.Xcalc [1]),
    .C(_3570_),
    .D(\genblk1[4].u_ce.Xcalc [3]),
    .Y(_3617_)
);

OAI21X1 _10248_ (
    .A(_3568_),
    .B(_3616_),
    .C(_3617_),
    .Y(\genblk1[4].u_ce.X_ [1])
);

INVX1 _10249_ (
    .A(\genblk1[4].u_ce.Ain0 [0]),
    .Y(_3618_)
);

NAND2X1 _10250_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\a[4] [0]),
    .Y(_3619_)
);

OAI21X1 _10251_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_3618_),
    .C(_3619_),
    .Y(_3464_)
);

INVX1 _10252_ (
    .A(\genblk1[4].u_ce.Ain0 [1]),
    .Y(_3620_)
);

NAND2X1 _10253_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\a[4] [1]),
    .Y(_3621_)
);

OAI21X1 _10254_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_3620_),
    .C(_3621_),
    .Y(_3465_)
);

INVX8 _10255_ (
    .A(\genblk1[4].u_ce.Vld_bF$buf4 ),
    .Y(_3622_)
);

NAND2X1 _10256_ (
    .A(\genblk1[4].u_ce.Ycalc [2]),
    .B(_3622__bF$buf4),
    .Y(_3623_)
);

INVX2 _10257_ (
    .A(1'h0),
    .Y(_3624_)
);

NOR2X1 _10258_ (
    .A(1'h1),
    .B(1'h0),
    .Y(_3625_)
);

NAND2X1 _10259_ (
    .A(_3624_),
    .B(_3625_),
    .Y(_3626_)
);

INVX2 _10260_ (
    .A(_3626_),
    .Y(_3627_)
);

INVX8 _10261_ (
    .A(1'h0),
    .Y(_3628_)
);

MUX2X1 _10262_ (
    .A(\genblk1[4].u_ce.Xin12b [4]),
    .B(\genblk1[4].u_ce.Xin1 [1]),
    .S(1'h0),
    .Y(_3629_)
);

MUX2X1 _10263_ (
    .A(\genblk1[4].u_ce.Xin1 [0]),
    .B(\genblk1[4].u_ce.Xin0 [1]),
    .S(1'h0),
    .Y(_3630_)
);

MUX2X1 _10264_ (
    .A(_3630_),
    .B(_3629_),
    .S(_3628__bF$buf4),
    .Y(_3631_)
);

MUX2X1 _10265_ (
    .A(\genblk1[4].u_ce.Xin12b [8]),
    .B(\genblk1[4].u_ce.Xin12b [7]),
    .S(1'h0),
    .Y(_3632_)
);

MUX2X1 _10266_ (
    .A(\genblk1[4].u_ce.Xin12b [6]),
    .B(\genblk1[4].u_ce.Xin12b [5]),
    .S(1'h0),
    .Y(_3633_)
);

MUX2X1 _10267_ (
    .A(_3633_),
    .B(_3632_),
    .S(_3628__bF$buf3),
    .Y(_3634_)
);

MUX2X1 _10268_ (
    .A(_3634_),
    .B(_3631_),
    .S(1'h1),
    .Y(_3635_)
);

INVX1 _10269_ (
    .A(_3635_),
    .Y(_3636_)
);

MUX2X1 _10270_ (
    .A(\genblk1[4].u_ce.Xin1 [1]),
    .B(\genblk1[4].u_ce.Xin1 [0]),
    .S(1'h0),
    .Y(_3637_)
);

MUX2X1 _10271_ (
    .A(\genblk1[4].u_ce.Xin0 [1]),
    .B(\genblk1[4].u_ce.Xin0 [0]),
    .S(1'h0),
    .Y(_3638_)
);

MUX2X1 _10272_ (
    .A(_3638_),
    .B(_3637_),
    .S(_3628__bF$buf2),
    .Y(_3639_)
);

MUX2X1 _10273_ (
    .A(\genblk1[4].u_ce.Xin12b [7]),
    .B(\genblk1[4].u_ce.Xin12b [6]),
    .S(1'h0),
    .Y(_3640_)
);

MUX2X1 _10274_ (
    .A(\genblk1[4].u_ce.Xin12b [5]),
    .B(\genblk1[4].u_ce.Xin12b [4]),
    .S(1'h0),
    .Y(_3641_)
);

MUX2X1 _10275_ (
    .A(_3641_),
    .B(_3640_),
    .S(_3628__bF$buf1),
    .Y(_3642_)
);

MUX2X1 _10276_ (
    .A(_3642_),
    .B(_3639_),
    .S(1'h1),
    .Y(_3643_)
);

OAI21X1 _10277_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf4 ),
    .B(_3643_),
    .C(_3636_),
    .Y(_3644_)
);

NOR2X1 _10278_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3643_),
    .Y(_3645_)
);

NAND2X1 _10279_ (
    .A(_3635_),
    .B(_3645_),
    .Y(_3646_)
);

NAND3X1 _10280_ (
    .A(\genblk1[4].u_ce.Yin0 [1]),
    .B(_3644_),
    .C(_3646_),
    .Y(_3647_)
);

NOR2X1 _10281_ (
    .A(\genblk1[4].u_ce.Yin0 [0]),
    .B(_3643_),
    .Y(_3648_)
);

AOI21X1 _10282_ (
    .A(_3646_),
    .B(_3644_),
    .C(\genblk1[4].u_ce.Yin0 [1]),
    .Y(_3649_)
);

OAI21X1 _10283_ (
    .A(_3648_),
    .B(_3649_),
    .C(_3647_),
    .Y(_3650_)
);

INVX1 _10284_ (
    .A(\genblk1[4].u_ce.Yin1 [0]),
    .Y(_3651_)
);

MUX2X1 _10285_ (
    .A(\genblk1[4].u_ce.Xin12b [9]),
    .B(\genblk1[4].u_ce.Xin12b [8]),
    .S(1'h0),
    .Y(_3652_)
);

MUX2X1 _10286_ (
    .A(_3652_),
    .B(_3640_),
    .S(1'h0),
    .Y(_3653_)
);

AND2X2 _10287_ (
    .A(_3653_),
    .B(1'h1),
    .Y(_3654_)
);

INVX4 _10288_ (
    .A(1'h1),
    .Y(_3655_)
);

NAND2X1 _10289_ (
    .A(_3655__bF$buf3),
    .B(_3628__bF$buf0),
    .Y(_3656_)
);

NAND2X1 _10290_ (
    .A(1'h0),
    .B(_3655__bF$buf2),
    .Y(_3657_)
);

OAI22X1 _10291_ (
    .A(_3656_),
    .B(_3637_),
    .C(_3641_),
    .D(_3657_),
    .Y(_3658_)
);

INVX1 _10292_ (
    .A(\genblk1[4].u_ce.Xin1 [1]),
    .Y(_3659_)
);

NAND2X1 _10293_ (
    .A(_3624_),
    .B(_3659_),
    .Y(_3660_)
);

INVX1 _10294_ (
    .A(\genblk1[4].u_ce.Xin12b [4]),
    .Y(_3661_)
);

NAND2X1 _10295_ (
    .A(1'h0),
    .B(_3661_),
    .Y(_3662_)
);

NAND3X1 _10296_ (
    .A(1'h0),
    .B(_3662_),
    .C(_3660_),
    .Y(_3663_)
);

INVX1 _10297_ (
    .A(\genblk1[4].u_ce.Xin0 [1]),
    .Y(_3664_)
);

NAND2X1 _10298_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Xin1 [0]),
    .Y(_3665_)
);

OAI21X1 _10299_ (
    .A(1'h0),
    .B(_3664_),
    .C(_3665_),
    .Y(_3666_)
);

NAND2X1 _10300_ (
    .A(_3628__bF$buf4),
    .B(_3666_),
    .Y(_3667_)
);

NAND3X1 _10301_ (
    .A(_3655__bF$buf1),
    .B(_3663_),
    .C(_3667_),
    .Y(_3668_)
);

INVX1 _10302_ (
    .A(\genblk1[4].u_ce.Xin12b [5]),
    .Y(_3669_)
);

NAND2X1 _10303_ (
    .A(_3624_),
    .B(_3669_),
    .Y(_3670_)
);

INVX1 _10304_ (
    .A(\genblk1[4].u_ce.Xin12b [6]),
    .Y(_3671_)
);

NAND2X1 _10305_ (
    .A(1'h0),
    .B(_3671_),
    .Y(_3672_)
);

NAND3X1 _10306_ (
    .A(_3628__bF$buf3),
    .B(_3672_),
    .C(_3670_),
    .Y(_3673_)
);

INVX1 _10307_ (
    .A(\genblk1[4].u_ce.Xin12b [7]),
    .Y(_3674_)
);

NAND2X1 _10308_ (
    .A(_3624_),
    .B(_3674_),
    .Y(_3675_)
);

INVX1 _10309_ (
    .A(\genblk1[4].u_ce.Xin12b [8]),
    .Y(_3676_)
);

NAND2X1 _10310_ (
    .A(1'h0),
    .B(_3676_),
    .Y(_3677_)
);

NAND3X1 _10311_ (
    .A(1'h0),
    .B(_3677_),
    .C(_3675_),
    .Y(_3678_)
);

NAND3X1 _10312_ (
    .A(1'h1),
    .B(_3673_),
    .C(_3678_),
    .Y(_3679_)
);

INVX1 _10313_ (
    .A(\genblk1[4].u_ce.Xin1 [0]),
    .Y(_3680_)
);

NAND2X1 _10314_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Xin1 [1]),
    .Y(_3681_)
);

OAI21X1 _10315_ (
    .A(1'h0),
    .B(_3680_),
    .C(_3681_),
    .Y(_3682_)
);

NAND2X1 _10316_ (
    .A(1'h0),
    .B(_3682_),
    .Y(_3683_)
);

INVX1 _10317_ (
    .A(\genblk1[4].u_ce.Xin0 [0]),
    .Y(_3684_)
);

NAND2X1 _10318_ (
    .A(\genblk1[4].u_ce.Xin0 [1]),
    .B(1'h0),
    .Y(_3685_)
);

OAI21X1 _10319_ (
    .A(1'h0),
    .B(_3684_),
    .C(_3685_),
    .Y(_3686_)
);

NAND2X1 _10320_ (
    .A(_3628__bF$buf2),
    .B(_3686_),
    .Y(_3687_)
);

NAND3X1 _10321_ (
    .A(_3655__bF$buf0),
    .B(_3683_),
    .C(_3687_),
    .Y(_3688_)
);

NAND2X1 _10322_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Xin12b [5]),
    .Y(_3689_)
);

OAI21X1 _10323_ (
    .A(1'h0),
    .B(_3661_),
    .C(_3689_),
    .Y(_3690_)
);

NAND2X1 _10324_ (
    .A(_3628__bF$buf1),
    .B(_3690_),
    .Y(_3691_)
);

NAND2X1 _10325_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Xin12b [7]),
    .Y(_3692_)
);

OAI21X1 _10326_ (
    .A(1'h0),
    .B(_3671_),
    .C(_3692_),
    .Y(_3693_)
);

NAND2X1 _10327_ (
    .A(1'h0),
    .B(_3693_),
    .Y(_3694_)
);

NAND3X1 _10328_ (
    .A(1'h1),
    .B(_3691_),
    .C(_3694_),
    .Y(_3695_)
);

AOI22X1 _10329_ (
    .A(_3668_),
    .B(_3679_),
    .C(_3688_),
    .D(_3695_),
    .Y(_3696_)
);

NOR2X1 _10330_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3696_),
    .Y(_3697_)
);

OAI21X1 _10331_ (
    .A(_3654_),
    .B(_3658_),
    .C(_3697_),
    .Y(_3698_)
);

AOI21X1 _10332_ (
    .A(1'h1),
    .B(_3653_),
    .C(_3658_),
    .Y(_3699_)
);

OAI21X1 _10333_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .B(_3696_),
    .C(_3699_),
    .Y(_3700_)
);

NAND3X1 _10334_ (
    .A(_3651_),
    .B(_3700_),
    .C(_3698_),
    .Y(_3701_)
);

NAND2X1 _10335_ (
    .A(_3699_),
    .B(_3697_),
    .Y(_3702_)
);

OAI22X1 _10336_ (
    .A(_3654_),
    .B(_3658_),
    .C(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .D(_3696_),
    .Y(_3703_)
);

NAND3X1 _10337_ (
    .A(\genblk1[4].u_ce.Yin1 [0]),
    .B(_3703_),
    .C(_3702_),
    .Y(_3704_)
);

NAND3X1 _10338_ (
    .A(_3701_),
    .B(_3704_),
    .C(_3650_),
    .Y(_3705_)
);

INVX1 _10339_ (
    .A(\genblk1[4].u_ce.Yin0 [1]),
    .Y(_3706_)
);

NAND2X1 _10340_ (
    .A(_3636_),
    .B(_3645_),
    .Y(_3707_)
);

OAI21X1 _10341_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf4 ),
    .B(_3643_),
    .C(_3635_),
    .Y(_3708_)
);

AOI21X1 _10342_ (
    .A(_3707_),
    .B(_3708_),
    .C(_3706_),
    .Y(_3709_)
);

INVX1 _10343_ (
    .A(_3648_),
    .Y(_3710_)
);

NAND3X1 _10344_ (
    .A(_3706_),
    .B(_3708_),
    .C(_3707_),
    .Y(_3711_)
);

AOI21X1 _10345_ (
    .A(_3710_),
    .B(_3711_),
    .C(_3709_),
    .Y(_3712_)
);

AOI21X1 _10346_ (
    .A(_3702_),
    .B(_3703_),
    .C(\genblk1[4].u_ce.Yin1 [0]),
    .Y(_3713_)
);

AOI21X1 _10347_ (
    .A(_3698_),
    .B(_3700_),
    .C(_3651_),
    .Y(_3714_)
);

OAI21X1 _10348_ (
    .A(_3713_),
    .B(_3714_),
    .C(_3712_),
    .Y(_3715_)
);

AOI21X1 _10349_ (
    .A(_3705_),
    .B(_3715_),
    .C(_3627_),
    .Y(_3716_)
);

INVX8 _10350_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_3717_)
);

NAND3X1 _10351_ (
    .A(_3655__bF$buf3),
    .B(_3624_),
    .C(_3717__bF$buf5),
    .Y(_3718_)
);

OAI21X1 _10352_ (
    .A(1'h0),
    .B(_3718_),
    .C(\genblk1[4].u_ce.Vld_bF$buf3 ),
    .Y(_3719_)
);

OAI21X1 _10353_ (
    .A(_3719_),
    .B(_3716_),
    .C(_3623_),
    .Y(_3466_)
);

INVX1 _10354_ (
    .A(\genblk1[4].u_ce.Ycalc [3]),
    .Y(_3720_)
);

INVX1 _10355_ (
    .A(\genblk1[4].u_ce.Xin12b [9]),
    .Y(_3721_)
);

NAND2X1 _10356_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Xin12b [10]),
    .Y(_3722_)
);

OAI21X1 _10357_ (
    .A(1'h0),
    .B(_3721_),
    .C(_3722_),
    .Y(_3723_)
);

NAND2X1 _10358_ (
    .A(1'h0),
    .B(_3723_),
    .Y(_3724_)
);

OAI21X1 _10359_ (
    .A(1'h0),
    .B(_3632_),
    .C(_3724_),
    .Y(_3725_)
);

OAI22X1 _10360_ (
    .A(_3656_),
    .B(_3629_),
    .C(_3633_),
    .D(_3657_),
    .Y(_3726_)
);

AOI21X1 _10361_ (
    .A(_3725_),
    .B(1'h1),
    .C(_3726_),
    .Y(_3727_)
);

NAND3X1 _10362_ (
    .A(_3699_),
    .B(_3635_),
    .C(_3643_),
    .Y(_3728_)
);

INVX1 _10363_ (
    .A(_3728_),
    .Y(_3729_)
);

NOR2X1 _10364_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3729_),
    .Y(_3730_)
);

NAND2X1 _10365_ (
    .A(_3727_),
    .B(_3730_),
    .Y(_3731_)
);

INVX1 _10366_ (
    .A(_3727_),
    .Y(_3732_)
);

OAI21X1 _10367_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .B(_3729_),
    .C(_3732_),
    .Y(_3733_)
);

AOI21X1 _10368_ (
    .A(_3731_),
    .B(_3733_),
    .C(\genblk1[4].u_ce.Yin1 [1]),
    .Y(_3734_)
);

AOI21X1 _10369_ (
    .A(_3650_),
    .B(_3701_),
    .C(_3714_),
    .Y(_3735_)
);

NAND3X1 _10370_ (
    .A(\genblk1[4].u_ce.Yin1 [1]),
    .B(_3733_),
    .C(_3731_),
    .Y(_3736_)
);

NAND2X1 _10371_ (
    .A(_3736_),
    .B(_3735_),
    .Y(_3737_)
);

OAI21X1 _10372_ (
    .A(_3713_),
    .B(_3712_),
    .C(_3704_),
    .Y(_3738_)
);

INVX1 _10373_ (
    .A(\genblk1[4].u_ce.Yin1 [1]),
    .Y(_3739_)
);

NAND2X1 _10374_ (
    .A(_3732_),
    .B(_3730_),
    .Y(_3740_)
);

OAI21X1 _10375_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .B(_3729_),
    .C(_3727_),
    .Y(_3741_)
);

AOI21X1 _10376_ (
    .A(_3740_),
    .B(_3741_),
    .C(_3739_),
    .Y(_3742_)
);

OAI21X1 _10377_ (
    .A(_3734_),
    .B(_3742_),
    .C(_3738_),
    .Y(_3743_)
);

OAI21X1 _10378_ (
    .A(_3734_),
    .B(_3737_),
    .C(_3743_),
    .Y(_3744_)
);

OAI21X1 _10379_ (
    .A(_3717__bF$buf4),
    .B(_3626_),
    .C(\genblk1[4].u_ce.Vld_bF$buf2 ),
    .Y(_3745_)
);

INVX1 _10380_ (
    .A(_3745_),
    .Y(_3746_)
);

OAI21X1 _10381_ (
    .A(_3627_),
    .B(_3744_),
    .C(_3746_),
    .Y(_3747_)
);

OAI21X1 _10382_ (
    .A(_3720_),
    .B(\genblk1[4].u_ce.Vld_bF$buf1 ),
    .C(_3747_),
    .Y(_3467_)
);

INVX1 _10383_ (
    .A(_3719_),
    .Y(_3748_)
);

INVX1 _10384_ (
    .A(\genblk1[4].u_ce.Yin12b [4]),
    .Y(_3749_)
);

NAND3X1 _10385_ (
    .A(_3699_),
    .B(_3727_),
    .C(_3696_),
    .Y(_3750_)
);

INVX1 _10386_ (
    .A(\genblk1[4].u_ce.Xin12b [10]),
    .Y(_3751_)
);

NAND2X1 _10387_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Xin12b [11]),
    .Y(_3752_)
);

OAI21X1 _10388_ (
    .A(1'h0),
    .B(_3751_),
    .C(_3752_),
    .Y(_3753_)
);

NAND2X1 _10389_ (
    .A(_3628__bF$buf0),
    .B(_3652_),
    .Y(_3754_)
);

OAI21X1 _10390_ (
    .A(_3628__bF$buf4),
    .B(_3753_),
    .C(_3754_),
    .Y(_3755_)
);

NAND2X1 _10391_ (
    .A(_3655__bF$buf2),
    .B(_3642_),
    .Y(_3756_)
);

OAI21X1 _10392_ (
    .A(_3655__bF$buf1),
    .B(_3755_),
    .C(_3756_),
    .Y(_3757_)
);

INVX1 _10393_ (
    .A(_3757_),
    .Y(_3758_)
);

NAND3X1 _10394_ (
    .A(_3717__bF$buf3),
    .B(_3758_),
    .C(_3750_),
    .Y(_3759_)
);

INVX1 _10395_ (
    .A(_3759_),
    .Y(_3760_)
);

AOI21X1 _10396_ (
    .A(_3750_),
    .B(_3717__bF$buf2),
    .C(_3758_),
    .Y(_3761_)
);

OAI21X1 _10397_ (
    .A(_3761_),
    .B(_3760_),
    .C(_3749_),
    .Y(_3762_)
);

OAI21X1 _10398_ (
    .A(_3728_),
    .B(_3732_),
    .C(_3717__bF$buf1),
    .Y(_3763_)
);

NAND2X1 _10399_ (
    .A(_3757_),
    .B(_3763_),
    .Y(_3764_)
);

NAND3X1 _10400_ (
    .A(\genblk1[4].u_ce.Yin12b [4]),
    .B(_3759_),
    .C(_3764_),
    .Y(_3765_)
);

NAND2X1 _10401_ (
    .A(_3765_),
    .B(_3762_),
    .Y(_3766_)
);

INVX1 _10402_ (
    .A(_3734_),
    .Y(_3767_)
);

OAI21X1 _10403_ (
    .A(_3742_),
    .B(_3738_),
    .C(_3767_),
    .Y(_3768_)
);

AOI21X1 _10404_ (
    .A(_3768_),
    .B(_3766_),
    .C(_3627_),
    .Y(_3769_)
);

OAI21X1 _10405_ (
    .A(_3766_),
    .B(_3768_),
    .C(_3769_),
    .Y(_3770_)
);

AOI22X1 _10406_ (
    .A(_3585_),
    .B(_3622__bF$buf3),
    .C(_3770_),
    .D(_3748_),
    .Y(_3468_)
);

INVX1 _10407_ (
    .A(_3765_),
    .Y(_3771_)
);

AOI21X1 _10408_ (
    .A(_3735_),
    .B(_3736_),
    .C(_3734_),
    .Y(_3772_)
);

AOI21X1 _10409_ (
    .A(_3772_),
    .B(_3762_),
    .C(_3771_),
    .Y(_3773_)
);

INVX1 _10410_ (
    .A(\genblk1[4].u_ce.Yin12b [5]),
    .Y(_3774_)
);

NAND3X1 _10411_ (
    .A(_3727_),
    .B(_3758_),
    .C(_3729_),
    .Y(_3775_)
);

INVX1 _10412_ (
    .A(\genblk1[4].u_ce.Xin12b [11]),
    .Y(_3776_)
);

NOR2X1 _10413_ (
    .A(_3628__bF$buf3),
    .B(_3776_),
    .Y(_3777_)
);

AOI21X1 _10414_ (
    .A(_3628__bF$buf2),
    .B(_3723_),
    .C(_3777_),
    .Y(_3778_)
);

NAND2X1 _10415_ (
    .A(_3655__bF$buf0),
    .B(_3634_),
    .Y(_3779_)
);

OAI21X1 _10416_ (
    .A(_3655__bF$buf3),
    .B(_3778_),
    .C(_3779_),
    .Y(_3780_)
);

NAND3X1 _10417_ (
    .A(_3717__bF$buf0),
    .B(_3780_),
    .C(_3775_),
    .Y(_3781_)
);

INVX1 _10418_ (
    .A(_3780_),
    .Y(_3782_)
);

OAI21X1 _10419_ (
    .A(_3757_),
    .B(_3750_),
    .C(_3717__bF$buf5),
    .Y(_3783_)
);

NAND2X1 _10420_ (
    .A(_3782_),
    .B(_3783_),
    .Y(_3784_)
);

NAND3X1 _10421_ (
    .A(_3774_),
    .B(_3784_),
    .C(_3781_),
    .Y(_3785_)
);

NAND3X1 _10422_ (
    .A(_3717__bF$buf4),
    .B(_3782_),
    .C(_3775_),
    .Y(_3786_)
);

NAND2X1 _10423_ (
    .A(_3780_),
    .B(_3783_),
    .Y(_3787_)
);

NAND3X1 _10424_ (
    .A(\genblk1[4].u_ce.Yin12b [5]),
    .B(_3787_),
    .C(_3786_),
    .Y(_3788_)
);

NAND2X1 _10425_ (
    .A(_3785_),
    .B(_3788_),
    .Y(_3789_)
);

INVX1 _10426_ (
    .A(_3789_),
    .Y(_3790_)
);

NOR2X1 _10427_ (
    .A(_3790_),
    .B(_3773_),
    .Y(_3791_)
);

OAI21X1 _10428_ (
    .A(_3766_),
    .B(_3768_),
    .C(_3765_),
    .Y(_3792_)
);

OAI21X1 _10429_ (
    .A(_3789_),
    .B(_3792_),
    .C(_3626_),
    .Y(_3793_)
);

OAI21X1 _10430_ (
    .A(_3793_),
    .B(_3791_),
    .C(_3748_),
    .Y(_3794_)
);

OAI21X1 _10431_ (
    .A(_3593_),
    .B(\genblk1[4].u_ce.Vld_bF$buf0 ),
    .C(_3794_),
    .Y(_3469_)
);

NOR2X1 _10432_ (
    .A(_3766_),
    .B(_3789_),
    .Y(_3795_)
);

OAI21X1 _10433_ (
    .A(_3765_),
    .B(_3789_),
    .C(_3788_),
    .Y(_3796_)
);

AOI21X1 _10434_ (
    .A(_3795_),
    .B(_3772_),
    .C(_3796_),
    .Y(_3797_)
);

INVX1 _10435_ (
    .A(\genblk1[4].u_ce.Yin12b [6]),
    .Y(_3798_)
);

NOR2X1 _10436_ (
    .A(_3757_),
    .B(_3750_),
    .Y(_3799_)
);

NAND2X1 _10437_ (
    .A(_3782_),
    .B(_3799_),
    .Y(_3800_)
);

AOI21X1 _10438_ (
    .A(_3628__bF$buf1),
    .B(_3753_),
    .C(_3777_),
    .Y(_3801_)
);

NAND2X1 _10439_ (
    .A(_3655__bF$buf2),
    .B(_3653_),
    .Y(_3802_)
);

OAI21X1 _10440_ (
    .A(_3655__bF$buf1),
    .B(_3801_),
    .C(_3802_),
    .Y(_3803_)
);

NAND3X1 _10441_ (
    .A(_3717__bF$buf3),
    .B(_3803_),
    .C(_3800_),
    .Y(_3804_)
);

NOR3X1 _10442_ (
    .A(_3757_),
    .B(_3780_),
    .C(_3750_),
    .Y(_3805_)
);

INVX1 _10443_ (
    .A(_3803_),
    .Y(_3806_)
);

OAI21X1 _10444_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf4 ),
    .B(_3805_),
    .C(_3806_),
    .Y(_3807_)
);

NAND3X1 _10445_ (
    .A(_3798_),
    .B(_3807_),
    .C(_3804_),
    .Y(_3808_)
);

NAND3X1 _10446_ (
    .A(_3717__bF$buf2),
    .B(_3806_),
    .C(_3800_),
    .Y(_3809_)
);

OAI21X1 _10447_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3805_),
    .C(_3803_),
    .Y(_3810_)
);

NAND3X1 _10448_ (
    .A(\genblk1[4].u_ce.Yin12b [6]),
    .B(_3810_),
    .C(_3809_),
    .Y(_3811_)
);

AND2X2 _10449_ (
    .A(_3808_),
    .B(_3811_),
    .Y(_3812_)
);

INVX1 _10450_ (
    .A(_3812_),
    .Y(_3813_)
);

AOI21X1 _10451_ (
    .A(_3797_),
    .B(_3813_),
    .C(_3627_),
    .Y(_3814_)
);

OAI21X1 _10452_ (
    .A(_3797_),
    .B(_3813_),
    .C(_3814_),
    .Y(_3815_)
);

AOI22X1 _10453_ (
    .A(_3584_),
    .B(_3622__bF$buf2),
    .C(_3815_),
    .D(_3748_),
    .Y(_3470_)
);

AND2X2 _10454_ (
    .A(_3762_),
    .B(_3765_),
    .Y(_3816_)
);

NAND3X1 _10455_ (
    .A(_3785_),
    .B(_3788_),
    .C(_3816_),
    .Y(_3817_)
);

INVX1 _10456_ (
    .A(_3788_),
    .Y(_3818_)
);

AOI21X1 _10457_ (
    .A(_3771_),
    .B(_3785_),
    .C(_3818_),
    .Y(_3819_)
);

OAI21X1 _10458_ (
    .A(_3768_),
    .B(_3817_),
    .C(_3819_),
    .Y(_3820_)
);

INVX1 _10459_ (
    .A(_3811_),
    .Y(_3821_)
);

AOI21X1 _10460_ (
    .A(_3820_),
    .B(_3808_),
    .C(_3821_),
    .Y(_3822_)
);

INVX1 _10461_ (
    .A(\genblk1[4].u_ce.Yin12b [7]),
    .Y(_3823_)
);

NAND2X1 _10462_ (
    .A(_3806_),
    .B(_3805_),
    .Y(_3824_)
);

NOR2X1 _10463_ (
    .A(_3655__bF$buf0),
    .B(_3776_),
    .Y(_3825_)
);

AOI21X1 _10464_ (
    .A(_3725_),
    .B(_3655__bF$buf3),
    .C(_3825_),
    .Y(_3826_)
);

INVX1 _10465_ (
    .A(_3826_),
    .Y(_3827_)
);

NAND3X1 _10466_ (
    .A(_3717__bF$buf1),
    .B(_3827_),
    .C(_3824_),
    .Y(_3828_)
);

AND2X2 _10467_ (
    .A(_3805_),
    .B(_3806_),
    .Y(_3829_)
);

OAI21X1 _10468_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3829_),
    .C(_3826_),
    .Y(_3830_)
);

NAND3X1 _10469_ (
    .A(_3823_),
    .B(_3828_),
    .C(_3830_),
    .Y(_3831_)
);

NAND3X1 _10470_ (
    .A(_3717__bF$buf0),
    .B(_3826_),
    .C(_3824_),
    .Y(_3832_)
);

OAI21X1 _10471_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .B(_3829_),
    .C(_3827_),
    .Y(_3833_)
);

NAND3X1 _10472_ (
    .A(\genblk1[4].u_ce.Yin12b [7]),
    .B(_3832_),
    .C(_3833_),
    .Y(_3834_)
);

AND2X2 _10473_ (
    .A(_3831_),
    .B(_3834_),
    .Y(_3835_)
);

NOR2X1 _10474_ (
    .A(_3835_),
    .B(_3822_),
    .Y(_3836_)
);

NAND2X1 _10475_ (
    .A(_3624_),
    .B(_3628__bF$buf0),
    .Y(_3837_)
);

NAND2X1 _10476_ (
    .A(_3835_),
    .B(_3822_),
    .Y(_3838_)
);

OAI21X1 _10477_ (
    .A(1'h1),
    .B(_3837_),
    .C(_3838_),
    .Y(_3839_)
);

OAI21X1 _10478_ (
    .A(_3836_),
    .B(_3839_),
    .C(_3746_),
    .Y(_3840_)
);

OAI21X1 _10479_ (
    .A(_3592_),
    .B(\genblk1[4].u_ce.Vld_bF$buf4 ),
    .C(_3840_),
    .Y(_3471_)
);

INVX1 _10480_ (
    .A(\genblk1[4].u_ce.Ycalc [8]),
    .Y(_3841_)
);

AOI21X1 _10481_ (
    .A(_3830_),
    .B(_3828_),
    .C(_3823_),
    .Y(_3842_)
);

OAI21X1 _10482_ (
    .A(_3821_),
    .B(_3842_),
    .C(_3831_),
    .Y(_3843_)
);

NAND3X1 _10483_ (
    .A(_3812_),
    .B(_3835_),
    .C(_3820_),
    .Y(_3844_)
);

INVX1 _10484_ (
    .A(\genblk1[4].u_ce.Yin12b [8]),
    .Y(_3845_)
);

NAND3X1 _10485_ (
    .A(_3806_),
    .B(_3826_),
    .C(_3805_),
    .Y(_3846_)
);

INVX1 _10486_ (
    .A(_3825_),
    .Y(_3847_)
);

OAI21X1 _10487_ (
    .A(1'h1),
    .B(_3755_),
    .C(_3847_),
    .Y(_3848_)
);

NAND3X1 _10488_ (
    .A(_3717__bF$buf5),
    .B(_3848_),
    .C(_3846_),
    .Y(_3849_)
);

INVX1 _10489_ (
    .A(_3848_),
    .Y(_3850_)
);

NAND2X1 _10490_ (
    .A(_3717__bF$buf4),
    .B(_3846_),
    .Y(_3851_)
);

NAND2X1 _10491_ (
    .A(_3850_),
    .B(_3851_),
    .Y(_3852_)
);

NAND3X1 _10492_ (
    .A(_3845_),
    .B(_3849_),
    .C(_3852_),
    .Y(_3853_)
);

NAND3X1 _10493_ (
    .A(_3717__bF$buf3),
    .B(_3850_),
    .C(_3846_),
    .Y(_3854_)
);

NAND2X1 _10494_ (
    .A(_3848_),
    .B(_3851_),
    .Y(_3855_)
);

NAND3X1 _10495_ (
    .A(\genblk1[4].u_ce.Yin12b [8]),
    .B(_3854_),
    .C(_3855_),
    .Y(_3856_)
);

AND2X2 _10496_ (
    .A(_3853_),
    .B(_3856_),
    .Y(_3857_)
);

INVX1 _10497_ (
    .A(_3857_),
    .Y(_3858_)
);

AOI21X1 _10498_ (
    .A(_3844_),
    .B(_3843_),
    .C(_3858_),
    .Y(_3859_)
);

NAND3X1 _10499_ (
    .A(_3831_),
    .B(_3834_),
    .C(_3812_),
    .Y(_3860_)
);

OAI21X1 _10500_ (
    .A(_3860_),
    .B(_3797_),
    .C(_3843_),
    .Y(_3861_)
);

OAI21X1 _10501_ (
    .A(_3857_),
    .B(_3861_),
    .C(_3626_),
    .Y(_3862_)
);

OR2X2 _10502_ (
    .A(_3862_),
    .B(_3859_),
    .Y(_3863_)
);

AOI22X1 _10503_ (
    .A(_3841_),
    .B(_3622__bF$buf1),
    .C(_3863_),
    .D(_3746_),
    .Y(_3472_)
);

INVX1 _10504_ (
    .A(\genblk1[4].u_ce.Ycalc [9]),
    .Y(_3864_)
);

INVX1 _10505_ (
    .A(_3856_),
    .Y(_3865_)
);

NOR2X1 _10506_ (
    .A(_3865_),
    .B(_3859_),
    .Y(_3866_)
);

INVX1 _10507_ (
    .A(\genblk1[4].u_ce.Yin12b [9]),
    .Y(_3867_)
);

OAI21X1 _10508_ (
    .A(1'h1),
    .B(_3778_),
    .C(_3847_),
    .Y(_3868_)
);

INVX1 _10509_ (
    .A(_3868_),
    .Y(_3869_)
);

OAI21X1 _10510_ (
    .A(_3848_),
    .B(_3846_),
    .C(_3717__bF$buf2),
    .Y(_3870_)
);

NAND2X1 _10511_ (
    .A(_3869_),
    .B(_3870_),
    .Y(_3871_)
);

NAND3X1 _10512_ (
    .A(_3826_),
    .B(_3850_),
    .C(_3829_),
    .Y(_3872_)
);

NAND3X1 _10513_ (
    .A(_3717__bF$buf1),
    .B(_3868_),
    .C(_3872_),
    .Y(_3873_)
);

NAND3X1 _10514_ (
    .A(_3867_),
    .B(_3871_),
    .C(_3873_),
    .Y(_3874_)
);

AND2X2 _10515_ (
    .A(_3870_),
    .B(_3869_),
    .Y(_3875_)
);

NOR2X1 _10516_ (
    .A(_3869_),
    .B(_3870_),
    .Y(_3876_)
);

OAI21X1 _10517_ (
    .A(_3876_),
    .B(_3875_),
    .C(\genblk1[4].u_ce.Yin12b [9]),
    .Y(_3877_)
);

NAND2X1 _10518_ (
    .A(_3874_),
    .B(_3877_),
    .Y(_3878_)
);

AOI21X1 _10519_ (
    .A(_3866_),
    .B(_3878_),
    .C(_3627_),
    .Y(_3879_)
);

OAI21X1 _10520_ (
    .A(_3866_),
    .B(_3878_),
    .C(_3879_),
    .Y(_3880_)
);

AOI22X1 _10521_ (
    .A(_3864_),
    .B(_3622__bF$buf0),
    .C(_3880_),
    .D(_3746_),
    .Y(_3473_)
);

OAI21X1 _10522_ (
    .A(_3856_),
    .B(_3878_),
    .C(_3877_),
    .Y(_3881_)
);

NAND3X1 _10523_ (
    .A(_3874_),
    .B(_3877_),
    .C(_3857_),
    .Y(_3882_)
);

AOI21X1 _10524_ (
    .A(_3843_),
    .B(_3844_),
    .C(_3882_),
    .Y(_3883_)
);

INVX1 _10525_ (
    .A(\genblk1[4].u_ce.Yin12b [10]),
    .Y(_3884_)
);

OAI21X1 _10526_ (
    .A(1'h1),
    .B(_3801_),
    .C(_3847_),
    .Y(_3885_)
);

INVX1 _10527_ (
    .A(_3885_),
    .Y(_3886_)
);

OAI21X1 _10528_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .B(_3869_),
    .C(_3870_),
    .Y(_3887_)
);

NAND2X1 _10529_ (
    .A(_3886_),
    .B(_3887_),
    .Y(_3888_)
);

OAI21X1 _10530_ (
    .A(_3868_),
    .B(_3872_),
    .C(_3717__bF$buf0),
    .Y(_3889_)
);

NAND2X1 _10531_ (
    .A(_3885_),
    .B(_3889_),
    .Y(_3890_)
);

NAND2X1 _10532_ (
    .A(_3888_),
    .B(_3890_),
    .Y(_3891_)
);

NAND2X1 _10533_ (
    .A(_3884_),
    .B(_3891_),
    .Y(_3892_)
);

NAND3X1 _10534_ (
    .A(\genblk1[4].u_ce.Yin12b [10]),
    .B(_3888_),
    .C(_3890_),
    .Y(_3893_)
);

AND2X2 _10535_ (
    .A(_3892_),
    .B(_3893_),
    .Y(_3894_)
);

OAI21X1 _10536_ (
    .A(_3881_),
    .B(_3883_),
    .C(_3894_),
    .Y(_3895_)
);

INVX1 _10537_ (
    .A(_3877_),
    .Y(_3896_)
);

AOI21X1 _10538_ (
    .A(_3865_),
    .B(_3874_),
    .C(_3896_),
    .Y(_3897_)
);

AND2X2 _10539_ (
    .A(_3877_),
    .B(_3874_),
    .Y(_3898_)
);

NAND3X1 _10540_ (
    .A(_3857_),
    .B(_3898_),
    .C(_3861_),
    .Y(_3899_)
);

NAND2X1 _10541_ (
    .A(_3893_),
    .B(_3892_),
    .Y(_3900_)
);

NAND3X1 _10542_ (
    .A(_3897_),
    .B(_3900_),
    .C(_3899_),
    .Y(_3901_)
);

NAND3X1 _10543_ (
    .A(_3626_),
    .B(_3901_),
    .C(_3895_),
    .Y(_3902_)
);

AOI22X1 _10544_ (
    .A(_3581_),
    .B(_3622__bF$buf4),
    .C(_3902_),
    .D(_3748_),
    .Y(_3474_)
);

INVX1 _10545_ (
    .A(_3893_),
    .Y(_3903_)
);

AOI21X1 _10546_ (
    .A(_3899_),
    .B(_3897_),
    .C(_3900_),
    .Y(_3904_)
);

OAI21X1 _10547_ (
    .A(_3885_),
    .B(_3887_),
    .C(_3717__bF$buf5),
    .Y(_3905_)
);

INVX1 _10548_ (
    .A(_3905_),
    .Y(_3906_)
);

NAND2X1 _10549_ (
    .A(\genblk1[4].u_ce.Yin12b [11]),
    .B(_3776_),
    .Y(_3907_)
);

INVX1 _10550_ (
    .A(\genblk1[4].u_ce.Yin12b [11]),
    .Y(_3908_)
);

NAND2X1 _10551_ (
    .A(\genblk1[4].u_ce.Xin12b [11]),
    .B(_3908_),
    .Y(_3909_)
);

NAND2X1 _10552_ (
    .A(_3907_),
    .B(_3909_),
    .Y(_3910_)
);

OR2X2 _10553_ (
    .A(_3906_),
    .B(_3910_),
    .Y(_3911_)
);

NAND2X1 _10554_ (
    .A(_3910_),
    .B(_3906_),
    .Y(_3912_)
);

NAND2X1 _10555_ (
    .A(_3912_),
    .B(_3911_),
    .Y(_3913_)
);

OAI21X1 _10556_ (
    .A(_3903_),
    .B(_3904_),
    .C(_3913_),
    .Y(_3914_)
);

INVX1 _10557_ (
    .A(_3913_),
    .Y(_3915_)
);

NAND3X1 _10558_ (
    .A(_3893_),
    .B(_3915_),
    .C(_3895_),
    .Y(_3916_)
);

NAND3X1 _10559_ (
    .A(_3626_),
    .B(_3916_),
    .C(_3914_),
    .Y(_3917_)
);

AOI22X1 _10560_ (
    .A(_3589_),
    .B(_3622__bF$buf3),
    .C(_3917_),
    .D(_3746_),
    .Y(_3475_)
);

INVX1 _10561_ (
    .A(\genblk1[4].u_ce.Ycalc [0]),
    .Y(_3918_)
);

OAI21X1 _10562_ (
    .A(1'h1),
    .B(_3837_),
    .C(\genblk1[4].u_ce.Vld_bF$buf3 ),
    .Y(_3919_)
);

INVX2 _10563_ (
    .A(_3919_),
    .Y(_3920_)
);

INVX1 _10564_ (
    .A(\genblk1[4].u_ce.Yin0 [0]),
    .Y(_3921_)
);

AOI21X1 _10565_ (
    .A(_3688_),
    .B(_3695_),
    .C(_3921_),
    .Y(_3922_)
);

OAI21X1 _10566_ (
    .A(_3922_),
    .B(_3648_),
    .C(_3920_),
    .Y(_3923_)
);

OAI21X1 _10567_ (
    .A(_3918_),
    .B(\genblk1[4].u_ce.Vld_bF$buf2 ),
    .C(_3923_),
    .Y(_3476_)
);

NAND2X1 _10568_ (
    .A(\genblk1[4].u_ce.Ycalc [1]),
    .B(_3622__bF$buf2),
    .Y(_3924_)
);

NAND3X1 _10569_ (
    .A(_3710_),
    .B(_3647_),
    .C(_3711_),
    .Y(_3925_)
);

OAI21X1 _10570_ (
    .A(_3709_),
    .B(_3649_),
    .C(_3648_),
    .Y(_3926_)
);

AOI21X1 _10571_ (
    .A(_3926_),
    .B(_3925_),
    .C(_3627_),
    .Y(_3927_)
);

OAI21X1 _10572_ (
    .A(_3622__bF$buf1),
    .B(_3927_),
    .C(_3924_),
    .Y(_3477_)
);

NAND2X1 _10573_ (
    .A(\genblk1[4].u_ce.Xcalc [0]),
    .B(_3622__bF$buf0),
    .Y(_3928_)
);

MUX2X1 _10574_ (
    .A(\genblk1[4].u_ce.Yin12b [7]),
    .B(\genblk1[4].u_ce.Yin12b [6]),
    .S(1'h0),
    .Y(_3929_)
);

NAND2X1 _10575_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin12b [5]),
    .Y(_3930_)
);

OAI21X1 _10576_ (
    .A(1'h0),
    .B(_3749_),
    .C(_3930_),
    .Y(_3931_)
);

NAND2X1 _10577_ (
    .A(_3628__bF$buf4),
    .B(_3931_),
    .Y(_3932_)
);

OAI21X1 _10578_ (
    .A(_3628__bF$buf3),
    .B(_3929_),
    .C(_3932_),
    .Y(_3933_)
);

NAND2X1 _10579_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin1 [1]),
    .Y(_3934_)
);

OAI21X1 _10580_ (
    .A(1'h0),
    .B(_3651_),
    .C(_3934_),
    .Y(_3935_)
);

NAND2X1 _10581_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin0 [1]),
    .Y(_3936_)
);

OAI21X1 _10582_ (
    .A(1'h0),
    .B(_3921_),
    .C(_3936_),
    .Y(_3937_)
);

MUX2X1 _10583_ (
    .A(_3937_),
    .B(_3935_),
    .S(_3628__bF$buf2),
    .Y(_3938_)
);

NAND2X1 _10584_ (
    .A(_3655__bF$buf2),
    .B(_3938_),
    .Y(_3939_)
);

OAI21X1 _10585_ (
    .A(_3655__bF$buf1),
    .B(_3933_),
    .C(_3939_),
    .Y(_3940_)
);

INVX1 _10586_ (
    .A(_3940_),
    .Y(_3941_)
);

NOR2X1 _10587_ (
    .A(\genblk1[4].u_ce.Xin0 [0]),
    .B(_3941_),
    .Y(_3942_)
);

OAI21X1 _10588_ (
    .A(_3684_),
    .B(_3940_),
    .C(_3920_),
    .Y(_3943_)
);

OAI21X1 _10589_ (
    .A(_3943_),
    .B(_3942_),
    .C(_3928_),
    .Y(_3478_)
);

NAND2X1 _10590_ (
    .A(\genblk1[4].u_ce.Xcalc [1]),
    .B(_3622__bF$buf4),
    .Y(_3944_)
);

NOR2X1 _10591_ (
    .A(_3684_),
    .B(_3940_),
    .Y(_3945_)
);

NAND2X1 _10592_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin12b [4]),
    .Y(_3946_)
);

OAI21X1 _10593_ (
    .A(1'h0),
    .B(_3739_),
    .C(_3946_),
    .Y(_3947_)
);

NAND2X1 _10594_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin1 [0]),
    .Y(_3948_)
);

OAI21X1 _10595_ (
    .A(1'h0),
    .B(_3706_),
    .C(_3948_),
    .Y(_3949_)
);

MUX2X1 _10596_ (
    .A(_3949_),
    .B(_3947_),
    .S(_3628__bF$buf1),
    .Y(_3950_)
);

NAND2X1 _10597_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin12b [8]),
    .Y(_3951_)
);

OAI21X1 _10598_ (
    .A(1'h0),
    .B(_3823_),
    .C(_3951_),
    .Y(_3952_)
);

NAND2X1 _10599_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin12b [6]),
    .Y(_3953_)
);

OAI21X1 _10600_ (
    .A(1'h0),
    .B(_3774_),
    .C(_3953_),
    .Y(_3954_)
);

MUX2X1 _10601_ (
    .A(_3954_),
    .B(_3952_),
    .S(_3628__bF$buf0),
    .Y(_3955_)
);

MUX2X1 _10602_ (
    .A(_3955_),
    .B(_3950_),
    .S(1'h1),
    .Y(_3956_)
);

NOR2X1 _10603_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf4 ),
    .B(_3940_),
    .Y(_3957_)
);

NAND2X1 _10604_ (
    .A(_3956_),
    .B(_3957_),
    .Y(_3958_)
);

NAND2X1 _10605_ (
    .A(_3655__bF$buf0),
    .B(_3950_),
    .Y(_3959_)
);

NAND2X1 _10606_ (
    .A(1'h1),
    .B(_3955_),
    .Y(_3960_)
);

NAND2X1 _10607_ (
    .A(_3959_),
    .B(_3960_),
    .Y(_3961_)
);

OAI21X1 _10608_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3940_),
    .C(_3961_),
    .Y(_3962_)
);

NAND3X1 _10609_ (
    .A(\genblk1[4].u_ce.Xin0 [1]),
    .B(_3962_),
    .C(_3958_),
    .Y(_3963_)
);

OAI21X1 _10610_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3940_),
    .C(_3956_),
    .Y(_3964_)
);

NAND2X1 _10611_ (
    .A(_3961_),
    .B(_3957_),
    .Y(_3965_)
);

NAND3X1 _10612_ (
    .A(_3664_),
    .B(_3964_),
    .C(_3965_),
    .Y(_3966_)
);

NAND3X1 _10613_ (
    .A(_3945_),
    .B(_3963_),
    .C(_3966_),
    .Y(_3967_)
);

INVX1 _10614_ (
    .A(_3945_),
    .Y(_3968_)
);

AOI21X1 _10615_ (
    .A(_3965_),
    .B(_3964_),
    .C(_3664_),
    .Y(_3969_)
);

AOI21X1 _10616_ (
    .A(_3958_),
    .B(_3962_),
    .C(\genblk1[4].u_ce.Xin0 [1]),
    .Y(_3970_)
);

OAI21X1 _10617_ (
    .A(_3969_),
    .B(_3970_),
    .C(_3968_),
    .Y(_3971_)
);

AOI21X1 _10618_ (
    .A(_3971_),
    .B(_3967_),
    .C(_3627_),
    .Y(_3972_)
);

OAI21X1 _10619_ (
    .A(_3622__bF$buf3),
    .B(_3972_),
    .C(_3944_),
    .Y(_3479_)
);

OAI21X1 _10620_ (
    .A(_3968_),
    .B(_3970_),
    .C(_3963_),
    .Y(_3973_)
);

MUX2X1 _10621_ (
    .A(\genblk1[4].u_ce.Yin12b [9]),
    .B(\genblk1[4].u_ce.Yin12b [8]),
    .S(1'h0),
    .Y(_3974_)
);

MUX2X1 _10622_ (
    .A(_3974_),
    .B(_3929_),
    .S(1'h0),
    .Y(_3975_)
);

NOR2X1 _10623_ (
    .A(1'h1),
    .B(_3628__bF$buf4),
    .Y(_3976_)
);

NAND2X1 _10624_ (
    .A(_3931_),
    .B(_3976_),
    .Y(_3977_)
);

NAND2X1 _10625_ (
    .A(_3625_),
    .B(_3935_),
    .Y(_3978_)
);

NAND2X1 _10626_ (
    .A(_3978_),
    .B(_3977_),
    .Y(_3979_)
);

AOI21X1 _10627_ (
    .A(1'h1),
    .B(_3975_),
    .C(_3979_),
    .Y(_3980_)
);

NAND2X1 _10628_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin12b [7]),
    .Y(_3981_)
);

OAI21X1 _10629_ (
    .A(1'h0),
    .B(_3798_),
    .C(_3981_),
    .Y(_3982_)
);

MUX2X1 _10630_ (
    .A(_3931_),
    .B(_3982_),
    .S(_3628__bF$buf3),
    .Y(_3983_)
);

NAND2X1 _10631_ (
    .A(1'h1),
    .B(_3983_),
    .Y(_3984_)
);

AOI21X1 _10632_ (
    .A(_3939_),
    .B(_3984_),
    .C(_3956_),
    .Y(_3985_)
);

NOR2X1 _10633_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .B(_3985_),
    .Y(_3986_)
);

NAND2X1 _10634_ (
    .A(_3980_),
    .B(_3986_),
    .Y(_3987_)
);

INVX1 _10635_ (
    .A(_3980_),
    .Y(_3988_)
);

OAI21X1 _10636_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .B(_3985_),
    .C(_3988_),
    .Y(_3989_)
);

AOI21X1 _10637_ (
    .A(_3987_),
    .B(_3989_),
    .C(_3680_),
    .Y(_3990_)
);

NAND3X1 _10638_ (
    .A(_3680_),
    .B(_3989_),
    .C(_3987_),
    .Y(_3991_)
);

INVX1 _10639_ (
    .A(_3991_),
    .Y(_3992_)
);

NOR2X1 _10640_ (
    .A(_3990_),
    .B(_3992_),
    .Y(_3993_)
);

NOR2X1 _10641_ (
    .A(_3973_),
    .B(_3993_),
    .Y(_3994_)
);

AOI21X1 _10642_ (
    .A(_3945_),
    .B(_3966_),
    .C(_3969_),
    .Y(_3995_)
);

INVX1 _10643_ (
    .A(_3993_),
    .Y(_3996_)
);

OAI21X1 _10644_ (
    .A(_3995_),
    .B(_3996_),
    .C(_3920_),
    .Y(_3997_)
);

OAI22X1 _10645_ (
    .A(_3597_),
    .B(\genblk1[4].u_ce.Vld_bF$buf1 ),
    .C(_3994_),
    .D(_3997_),
    .Y(_3480_)
);

NAND2X1 _10646_ (
    .A(\genblk1[4].u_ce.Xcalc [3]),
    .B(_3622__bF$buf2),
    .Y(_3998_)
);

AOI21X1 _10647_ (
    .A(_3973_),
    .B(_3991_),
    .C(_3990_),
    .Y(_3999_)
);

NAND2X1 _10648_ (
    .A(1'h0),
    .B(_3884_),
    .Y(_4000_)
);

OAI21X1 _10649_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin12b [9]),
    .C(_4000_),
    .Y(_4001_)
);

NAND2X1 _10650_ (
    .A(_3628__bF$buf2),
    .B(_3952_),
    .Y(_4002_)
);

OAI21X1 _10651_ (
    .A(_3628__bF$buf1),
    .B(_4001_),
    .C(_4002_),
    .Y(_4003_)
);

NAND2X1 _10652_ (
    .A(_3954_),
    .B(_3976_),
    .Y(_4004_)
);

NAND2X1 _10653_ (
    .A(_3625_),
    .B(_3947_),
    .Y(_4005_)
);

NAND2X1 _10654_ (
    .A(_4005_),
    .B(_4004_),
    .Y(_4006_)
);

AOI21X1 _10655_ (
    .A(_4003_),
    .B(1'h1),
    .C(_4006_),
    .Y(_4007_)
);

NAND3X1 _10656_ (
    .A(_3980_),
    .B(_3961_),
    .C(_3940_),
    .Y(_4008_)
);

NAND2X1 _10657_ (
    .A(_3717__bF$buf4),
    .B(_4008_),
    .Y(_4009_)
);

OR2X2 _10658_ (
    .A(_4009_),
    .B(_4007_),
    .Y(_4010_)
);

INVX1 _10659_ (
    .A(_4008_),
    .Y(_4011_)
);

OAI21X1 _10660_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf4 ),
    .B(_4011_),
    .C(_4007_),
    .Y(_4012_)
);

NAND3X1 _10661_ (
    .A(\genblk1[4].u_ce.Xin1 [1]),
    .B(_4012_),
    .C(_4010_),
    .Y(_4013_)
);

INVX1 _10662_ (
    .A(_4007_),
    .Y(_4014_)
);

OR2X2 _10663_ (
    .A(_4009_),
    .B(_4014_),
    .Y(_4015_)
);

OAI21X1 _10664_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4011_),
    .C(_4014_),
    .Y(_4016_)
);

NAND3X1 _10665_ (
    .A(_3659_),
    .B(_4016_),
    .C(_4015_),
    .Y(_4017_)
);

NAND2X1 _10666_ (
    .A(_4013_),
    .B(_4017_),
    .Y(_4018_)
);

OR2X2 _10667_ (
    .A(_3999_),
    .B(_4018_),
    .Y(_4019_)
);

NAND2X1 _10668_ (
    .A(_4018_),
    .B(_3999_),
    .Y(_4020_)
);

AOI21X1 _10669_ (
    .A(_4019_),
    .B(_4020_),
    .C(_3627_),
    .Y(_4021_)
);

OAI21X1 _10670_ (
    .A(_3622__bF$buf1),
    .B(_4021_),
    .C(_3998_),
    .Y(_3481_)
);

OAI21X1 _10671_ (
    .A(_4018_),
    .B(_3999_),
    .C(_4013_),
    .Y(_4022_)
);

NAND2X1 _10672_ (
    .A(1'h0),
    .B(\genblk1[4].u_ce.Yin12b [11]),
    .Y(_4023_)
);

OAI21X1 _10673_ (
    .A(1'h0),
    .B(_3884_),
    .C(_4023_),
    .Y(_4024_)
);

NAND2X1 _10674_ (
    .A(1'h0),
    .B(_4024_),
    .Y(_4025_)
);

OAI21X1 _10675_ (
    .A(1'h0),
    .B(_3974_),
    .C(_4025_),
    .Y(_4026_)
);

NAND2X1 _10676_ (
    .A(1'h1),
    .B(_4026_),
    .Y(_4027_)
);

OAI21X1 _10677_ (
    .A(1'h1),
    .B(_3983_),
    .C(_4027_),
    .Y(_4028_)
);

INVX1 _10678_ (
    .A(_4028_),
    .Y(_4029_)
);

OAI21X1 _10679_ (
    .A(_4014_),
    .B(_4008_),
    .C(_3717__bF$buf3),
    .Y(_4030_)
);

OR2X2 _10680_ (
    .A(_4030_),
    .B(_4029_),
    .Y(_4031_)
);

NAND2X1 _10681_ (
    .A(_4029_),
    .B(_4030_),
    .Y(_4032_)
);

NAND3X1 _10682_ (
    .A(\genblk1[4].u_ce.Xin12b [4]),
    .B(_4032_),
    .C(_4031_),
    .Y(_4033_)
);

OR2X2 _10683_ (
    .A(_4030_),
    .B(_4028_),
    .Y(_4034_)
);

NAND2X1 _10684_ (
    .A(_4028_),
    .B(_4030_),
    .Y(_4035_)
);

NAND3X1 _10685_ (
    .A(_3661_),
    .B(_4035_),
    .C(_4034_),
    .Y(_4036_)
);

AND2X2 _10686_ (
    .A(_4033_),
    .B(_4036_),
    .Y(_4037_)
);

NAND2X1 _10687_ (
    .A(_4037_),
    .B(_4022_),
    .Y(_4038_)
);

INVX1 _10688_ (
    .A(_3990_),
    .Y(_4039_)
);

OAI21X1 _10689_ (
    .A(_3992_),
    .B(_3995_),
    .C(_4039_),
    .Y(_4040_)
);

INVX1 _10690_ (
    .A(_4013_),
    .Y(_4041_)
);

AOI21X1 _10691_ (
    .A(_4040_),
    .B(_4017_),
    .C(_4041_),
    .Y(_4042_)
);

NAND2X1 _10692_ (
    .A(_4036_),
    .B(_4033_),
    .Y(_4043_)
);

NAND2X1 _10693_ (
    .A(_4043_),
    .B(_4042_),
    .Y(_4044_)
);

NAND2X1 _10694_ (
    .A(_4038_),
    .B(_4044_),
    .Y(_4045_)
);

AOI22X1 _10695_ (
    .A(_3599_),
    .B(_3622__bF$buf0),
    .C(_4045_),
    .D(_3920_),
    .Y(_3482_)
);

NAND3X1 _10696_ (
    .A(_4007_),
    .B(_4029_),
    .C(_4011_),
    .Y(_4046_)
);

NOR2X1 _10697_ (
    .A(1'h0),
    .B(_4001_),
    .Y(_4047_)
);

NOR2X1 _10698_ (
    .A(_3628__bF$buf0),
    .B(_3908_),
    .Y(_4048_)
);

OAI21X1 _10699_ (
    .A(_4048_),
    .B(_4047_),
    .C(1'h1),
    .Y(_4049_)
);

OAI21X1 _10700_ (
    .A(1'h1),
    .B(_3955_),
    .C(_4049_),
    .Y(_4050_)
);

NAND3X1 _10701_ (
    .A(_3717__bF$buf2),
    .B(_4050_),
    .C(_4046_),
    .Y(_4051_)
);

INVX1 _10702_ (
    .A(_4050_),
    .Y(_4052_)
);

NAND3X1 _10703_ (
    .A(_3980_),
    .B(_4007_),
    .C(_3985_),
    .Y(_4053_)
);

OAI21X1 _10704_ (
    .A(_4028_),
    .B(_4053_),
    .C(_3717__bF$buf1),
    .Y(_4054_)
);

NAND2X1 _10705_ (
    .A(_4052_),
    .B(_4054_),
    .Y(_4055_)
);

NAND3X1 _10706_ (
    .A(\genblk1[4].u_ce.Xin12b [5]),
    .B(_4055_),
    .C(_4051_),
    .Y(_4056_)
);

NAND3X1 _10707_ (
    .A(_3717__bF$buf0),
    .B(_4052_),
    .C(_4046_),
    .Y(_4057_)
);

NAND2X1 _10708_ (
    .A(_4050_),
    .B(_4054_),
    .Y(_4058_)
);

NAND3X1 _10709_ (
    .A(_3669_),
    .B(_4058_),
    .C(_4057_),
    .Y(_4059_)
);

NAND2X1 _10710_ (
    .A(_4056_),
    .B(_4059_),
    .Y(_4060_)
);

AOI21X1 _10711_ (
    .A(_4038_),
    .B(_4033_),
    .C(_4060_),
    .Y(_4061_)
);

OAI21X1 _10712_ (
    .A(_4043_),
    .B(_4042_),
    .C(_4033_),
    .Y(_4062_)
);

AND2X2 _10713_ (
    .A(_4056_),
    .B(_4059_),
    .Y(_4063_)
);

OAI21X1 _10714_ (
    .A(_4063_),
    .B(_4062_),
    .C(_3920_),
    .Y(_4064_)
);

OAI22X1 _10715_ (
    .A(_3614_),
    .B(\genblk1[4].u_ce.Vld_bF$buf0 ),
    .C(_4061_),
    .D(_4064_),
    .Y(_3483_)
);

NOR2X1 _10716_ (
    .A(_4028_),
    .B(_4053_),
    .Y(_4065_)
);

NAND2X1 _10717_ (
    .A(_4052_),
    .B(_4065_),
    .Y(_4066_)
);

AOI21X1 _10718_ (
    .A(_3628__bF$buf4),
    .B(_4024_),
    .C(_4048_),
    .Y(_4067_)
);

NAND2X1 _10719_ (
    .A(_3655__bF$buf3),
    .B(_3975_),
    .Y(_4068_)
);

OAI21X1 _10720_ (
    .A(_3655__bF$buf2),
    .B(_4067_),
    .C(_4068_),
    .Y(_4069_)
);

NAND3X1 _10721_ (
    .A(_3717__bF$buf5),
    .B(_4069_),
    .C(_4066_),
    .Y(_4070_)
);

NOR3X1 _10722_ (
    .A(_4028_),
    .B(_4050_),
    .C(_4053_),
    .Y(_4071_)
);

INVX1 _10723_ (
    .A(_4069_),
    .Y(_4072_)
);

OAI21X1 _10724_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4071_),
    .C(_4072_),
    .Y(_4073_)
);

NAND3X1 _10725_ (
    .A(\genblk1[4].u_ce.Xin12b [6]),
    .B(_4073_),
    .C(_4070_),
    .Y(_4074_)
);

NAND3X1 _10726_ (
    .A(_3717__bF$buf4),
    .B(_4072_),
    .C(_4066_),
    .Y(_4075_)
);

OAI21X1 _10727_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .B(_4071_),
    .C(_4069_),
    .Y(_4076_)
);

NAND3X1 _10728_ (
    .A(_3671_),
    .B(_4076_),
    .C(_4075_),
    .Y(_4077_)
);

AND2X2 _10729_ (
    .A(_4074_),
    .B(_4077_),
    .Y(_4078_)
);

NAND2X1 _10730_ (
    .A(_4037_),
    .B(_4063_),
    .Y(_4079_)
);

INVX1 _10731_ (
    .A(_4033_),
    .Y(_4080_)
);

INVX1 _10732_ (
    .A(_4056_),
    .Y(_4081_)
);

AOI21X1 _10733_ (
    .A(_4080_),
    .B(_4059_),
    .C(_4081_),
    .Y(_4082_)
);

OAI21X1 _10734_ (
    .A(_4042_),
    .B(_4079_),
    .C(_4082_),
    .Y(_4083_)
);

AND2X2 _10735_ (
    .A(_4083_),
    .B(_4078_),
    .Y(_4084_)
);

NOR2X1 _10736_ (
    .A(_4078_),
    .B(_4083_),
    .Y(_4085_)
);

OAI21X1 _10737_ (
    .A(_4085_),
    .B(_4084_),
    .C(_3626_),
    .Y(_4086_)
);

NAND2X1 _10738_ (
    .A(\genblk1[4].u_ce.Vld_bF$buf4 ),
    .B(_4086_),
    .Y(_4087_)
);

OAI21X1 _10739_ (
    .A(_3600_),
    .B(\genblk1[4].u_ce.Vld_bF$buf3 ),
    .C(_4087_),
    .Y(_3484_)
);

INVX1 _10740_ (
    .A(_4074_),
    .Y(_4088_)
);

NOR2X1 _10741_ (
    .A(_4088_),
    .B(_4084_),
    .Y(_4089_)
);

NAND2X1 _10742_ (
    .A(_4072_),
    .B(_4071_),
    .Y(_4090_)
);

NOR2X1 _10743_ (
    .A(_3655__bF$buf1),
    .B(_3908_),
    .Y(_4091_)
);

AOI21X1 _10744_ (
    .A(_4003_),
    .B(_3655__bF$buf0),
    .C(_4091_),
    .Y(_4092_)
);

NAND3X1 _10745_ (
    .A(_3717__bF$buf3),
    .B(_4092_),
    .C(_4090_),
    .Y(_4093_)
);

INVX1 _10746_ (
    .A(_4093_),
    .Y(_4094_)
);

AOI21X1 _10747_ (
    .A(_4090_),
    .B(_3717__bF$buf2),
    .C(_4092_),
    .Y(_4095_)
);

OAI21X1 _10748_ (
    .A(_4095_),
    .B(_4094_),
    .C(\genblk1[4].u_ce.Xin12b [7]),
    .Y(_4096_)
);

INVX1 _10749_ (
    .A(_4095_),
    .Y(_4097_)
);

NAND3X1 _10750_ (
    .A(_3674_),
    .B(_4093_),
    .C(_4097_),
    .Y(_4098_)
);

AND2X2 _10751_ (
    .A(_4098_),
    .B(_4096_),
    .Y(_4099_)
);

OR2X2 _10752_ (
    .A(_4089_),
    .B(_4099_),
    .Y(_4100_)
);

AOI21X1 _10753_ (
    .A(_4089_),
    .B(_4099_),
    .C(_3919_),
    .Y(_4101_)
);

AOI22X1 _10754_ (
    .A(_3613_),
    .B(_3622__bF$buf4),
    .C(_4100_),
    .D(_4101_),
    .Y(_3485_)
);

NOR2X1 _10755_ (
    .A(_4043_),
    .B(_4060_),
    .Y(_4102_)
);

OAI21X1 _10756_ (
    .A(_4033_),
    .B(_4060_),
    .C(_4056_),
    .Y(_4103_)
);

AOI21X1 _10757_ (
    .A(_4102_),
    .B(_4022_),
    .C(_4103_),
    .Y(_4104_)
);

AOI21X1 _10758_ (
    .A(_4097_),
    .B(_4093_),
    .C(_3674_),
    .Y(_4105_)
);

AOI21X1 _10759_ (
    .A(_4088_),
    .B(_4098_),
    .C(_4105_),
    .Y(_4106_)
);

NAND3X1 _10760_ (
    .A(_4078_),
    .B(_4096_),
    .C(_4098_),
    .Y(_4107_)
);

OAI21X1 _10761_ (
    .A(_4107_),
    .B(_4104_),
    .C(_4106_),
    .Y(_4108_)
);

NAND3X1 _10762_ (
    .A(_4072_),
    .B(_4092_),
    .C(_4071_),
    .Y(_4109_)
);

INVX1 _10763_ (
    .A(_4026_),
    .Y(_4110_)
);

INVX1 _10764_ (
    .A(_4091_),
    .Y(_4111_)
);

OAI21X1 _10765_ (
    .A(1'h1),
    .B(_4110_),
    .C(_4111_),
    .Y(_4112_)
);

INVX1 _10766_ (
    .A(_4112_),
    .Y(_4113_)
);

NAND3X1 _10767_ (
    .A(_3717__bF$buf1),
    .B(_4113_),
    .C(_4109_),
    .Y(_4114_)
);

INVX1 _10768_ (
    .A(_4114_),
    .Y(_4115_)
);

AOI21X1 _10769_ (
    .A(_4109_),
    .B(_3717__bF$buf0),
    .C(_4113_),
    .Y(_4116_)
);

OAI21X1 _10770_ (
    .A(_4116_),
    .B(_4115_),
    .C(\genblk1[4].u_ce.Xin12b [8]),
    .Y(_4117_)
);

INVX1 _10771_ (
    .A(_4116_),
    .Y(_4118_)
);

NAND3X1 _10772_ (
    .A(_3676_),
    .B(_4114_),
    .C(_4118_),
    .Y(_4119_)
);

AND2X2 _10773_ (
    .A(_4119_),
    .B(_4117_),
    .Y(_4120_)
);

OR2X2 _10774_ (
    .A(_4108_),
    .B(_4120_),
    .Y(_4121_)
);

INVX1 _10775_ (
    .A(_4121_),
    .Y(_4122_)
);

NAND2X1 _10776_ (
    .A(_4120_),
    .B(_4108_),
    .Y(_4123_)
);

NAND2X1 _10777_ (
    .A(_3920_),
    .B(_4123_),
    .Y(_4124_)
);

OAI22X1 _10778_ (
    .A(_3602_),
    .B(\genblk1[4].u_ce.Vld_bF$buf2 ),
    .C(_4124_),
    .D(_4122_),
    .Y(_3486_)
);

NOR3X1 _10779_ (
    .A(_4050_),
    .B(_4069_),
    .C(_4046_),
    .Y(_4125_)
);

NAND3X1 _10780_ (
    .A(_4092_),
    .B(_4113_),
    .C(_4125_),
    .Y(_4126_)
);

OR2X2 _10781_ (
    .A(_4047_),
    .B(_4048_),
    .Y(_4127_)
);

AOI21X1 _10782_ (
    .A(_4127_),
    .B(_3655__bF$buf3),
    .C(_4091_),
    .Y(_4128_)
);

INVX1 _10783_ (
    .A(_4128_),
    .Y(_4129_)
);

NAND3X1 _10784_ (
    .A(_3717__bF$buf5),
    .B(_4129_),
    .C(_4126_),
    .Y(_4130_)
);

OAI21X1 _10785_ (
    .A(_4112_),
    .B(_4109_),
    .C(_3717__bF$buf4),
    .Y(_4131_)
);

NAND2X1 _10786_ (
    .A(_4128_),
    .B(_4131_),
    .Y(_4132_)
);

NAND3X1 _10787_ (
    .A(\genblk1[4].u_ce.Xin12b [9]),
    .B(_4132_),
    .C(_4130_),
    .Y(_4133_)
);

NAND3X1 _10788_ (
    .A(_3717__bF$buf3),
    .B(_4128_),
    .C(_4126_),
    .Y(_4134_)
);

NAND2X1 _10789_ (
    .A(_4129_),
    .B(_4131_),
    .Y(_4135_)
);

NAND3X1 _10790_ (
    .A(_3721_),
    .B(_4135_),
    .C(_4134_),
    .Y(_4136_)
);

NAND2X1 _10791_ (
    .A(_4133_),
    .B(_4136_),
    .Y(_4137_)
);

AOI21X1 _10792_ (
    .A(_4123_),
    .B(_4117_),
    .C(_4137_),
    .Y(_4138_)
);

NAND3X1 _10793_ (
    .A(_4117_),
    .B(_4137_),
    .C(_4123_),
    .Y(_4139_)
);

NAND2X1 _10794_ (
    .A(_3920_),
    .B(_4139_),
    .Y(_4140_)
);

OAI22X1 _10795_ (
    .A(_3610_),
    .B(\genblk1[4].u_ce.Vld_bF$buf1 ),
    .C(_4138_),
    .D(_4140_),
    .Y(_3487_)
);

NAND2X1 _10796_ (
    .A(\genblk1[4].u_ce.Xcalc [10]),
    .B(_3622__bF$buf3),
    .Y(_4141_)
);

OAI21X1 _10797_ (
    .A(1'h1),
    .B(_4067_),
    .C(_4111_),
    .Y(_4142_)
);

OAI21X1 _10798_ (
    .A(_4129_),
    .B(_4126_),
    .C(_3717__bF$buf2),
    .Y(_4143_)
);

NOR2X1 _10799_ (
    .A(_4142_),
    .B(_4143_),
    .Y(_4144_)
);

NAND2X1 _10800_ (
    .A(_4142_),
    .B(_4143_),
    .Y(_4145_)
);

INVX1 _10801_ (
    .A(_4145_),
    .Y(_4146_)
);

OAI21X1 _10802_ (
    .A(_4144_),
    .B(_4146_),
    .C(\genblk1[4].u_ce.Xin12b [10]),
    .Y(_4147_)
);

INVX1 _10803_ (
    .A(_4144_),
    .Y(_4148_)
);

NAND3X1 _10804_ (
    .A(_3751_),
    .B(_4145_),
    .C(_4148_),
    .Y(_4149_)
);

AND2X2 _10805_ (
    .A(_4149_),
    .B(_4147_),
    .Y(_4150_)
);

OAI21X1 _10806_ (
    .A(_4117_),
    .B(_4137_),
    .C(_4133_),
    .Y(_4151_)
);

NAND3X1 _10807_ (
    .A(_4078_),
    .B(_4083_),
    .C(_4099_),
    .Y(_4152_)
);

NAND3X1 _10808_ (
    .A(_4133_),
    .B(_4136_),
    .C(_4120_),
    .Y(_4153_)
);

AOI21X1 _10809_ (
    .A(_4152_),
    .B(_4106_),
    .C(_4153_),
    .Y(_4154_)
);

OAI21X1 _10810_ (
    .A(_4151_),
    .B(_4154_),
    .C(_4150_),
    .Y(_4155_)
);

NAND2X1 _10811_ (
    .A(_4147_),
    .B(_4149_),
    .Y(_4156_)
);

NAND2X1 _10812_ (
    .A(_4117_),
    .B(_4119_),
    .Y(_4157_)
);

NOR2X1 _10813_ (
    .A(_4157_),
    .B(_4137_),
    .Y(_4158_)
);

AOI21X1 _10814_ (
    .A(_4108_),
    .B(_4158_),
    .C(_4151_),
    .Y(_4159_)
);

NAND2X1 _10815_ (
    .A(_4156_),
    .B(_4159_),
    .Y(_4160_)
);

AOI21X1 _10816_ (
    .A(_4155_),
    .B(_4160_),
    .C(_3627_),
    .Y(_4161_)
);

OAI21X1 _10817_ (
    .A(_3622__bF$buf2),
    .B(_4161_),
    .C(_4141_),
    .Y(_3488_)
);

NAND2X1 _10818_ (
    .A(\genblk1[4].u_ce.Xcalc [11]),
    .B(_3622__bF$buf1),
    .Y(_4162_)
);

OR2X2 _10819_ (
    .A(_4126_),
    .B(_4129_),
    .Y(_4163_)
);

OAI21X1 _10820_ (
    .A(_4142_),
    .B(_4163_),
    .C(_3717__bF$buf1),
    .Y(_4164_)
);

OR2X2 _10821_ (
    .A(_4164_),
    .B(_3910_),
    .Y(_4165_)
);

NAND2X1 _10822_ (
    .A(_3910_),
    .B(_4164_),
    .Y(_4166_)
);

AOI22X1 _10823_ (
    .A(_4165_),
    .B(_4166_),
    .C(_4155_),
    .D(_4147_),
    .Y(_4167_)
);

OAI21X1 _10824_ (
    .A(_4156_),
    .B(_4159_),
    .C(_4147_),
    .Y(_4168_)
);

NAND2X1 _10825_ (
    .A(_4166_),
    .B(_4165_),
    .Y(_4169_)
);

OAI21X1 _10826_ (
    .A(_4169_),
    .B(_4168_),
    .C(_3920_),
    .Y(_4170_)
);

OAI21X1 _10827_ (
    .A(_4167_),
    .B(_4170_),
    .C(_4162_),
    .Y(_3489_)
);

NAND2X1 _10828_ (
    .A(1'h0),
    .B(1'h0),
    .Y(_4171_)
);

OAI21X1 _10829_ (
    .A(_3655__bF$buf2),
    .B(_3837_),
    .C(_4171_),
    .Y(_4172_)
);

NOR2X1 _10830_ (
    .A(_3618_),
    .B(_4172_),
    .Y(_4173_)
);

AND2X2 _10831_ (
    .A(_4172_),
    .B(_3618_),
    .Y(_4174_)
);

OR2X2 _10832_ (
    .A(_4174_),
    .B(_4173_),
    .Y(_4175_)
);

NAND2X1 _10833_ (
    .A(\genblk1[4].u_ce.Acalc [0]),
    .B(_3622__bF$buf0),
    .Y(_4176_)
);

OAI21X1 _10834_ (
    .A(_3622__bF$buf4),
    .B(_4175_),
    .C(_4176_),
    .Y(_3490_)
);

NAND2X1 _10835_ (
    .A(\genblk1[4].u_ce.Acalc [1]),
    .B(_3622__bF$buf3),
    .Y(_4177_)
);

OAI21X1 _10836_ (
    .A(1'h0),
    .B(_3624_),
    .C(1'h1),
    .Y(_4178_)
);

OAI21X1 _10837_ (
    .A(1'h1),
    .B(_3624_),
    .C(_4178_),
    .Y(_4179_)
);

OAI21X1 _10838_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .B(_4172_),
    .C(_4179_),
    .Y(_4180_)
);

OAI21X1 _10839_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf4 ),
    .B(_4179_),
    .C(_4180_),
    .Y(_4181_)
);

OR2X2 _10840_ (
    .A(_4181_),
    .B(\genblk1[4].u_ce.Ain0 [1]),
    .Y(_4182_)
);

NAND2X1 _10841_ (
    .A(\genblk1[4].u_ce.Ain0 [1]),
    .B(_4181_),
    .Y(_4183_)
);

NAND2X1 _10842_ (
    .A(_4183_),
    .B(_4182_),
    .Y(_4184_)
);

NOR2X1 _10843_ (
    .A(_4173_),
    .B(_4184_),
    .Y(_4185_)
);

NAND2X1 _10844_ (
    .A(_4173_),
    .B(_4184_),
    .Y(_4186_)
);

NAND2X1 _10845_ (
    .A(\genblk1[4].u_ce.Vld_bF$buf0 ),
    .B(_4186_),
    .Y(_4187_)
);

OAI21X1 _10846_ (
    .A(_4185_),
    .B(_4187_),
    .C(_4177_),
    .Y(_3491_)
);

NAND2X1 _10847_ (
    .A(\genblk1[4].u_ce.Acalc [2]),
    .B(_3622__bF$buf2),
    .Y(_4188_)
);

OAI21X1 _10848_ (
    .A(_3620_),
    .B(_4181_),
    .C(_4186_),
    .Y(_4189_)
);

OAI21X1 _10849_ (
    .A(_3624_),
    .B(_3628__bF$buf3),
    .C(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_4190_)
);

NAND3X1 _10850_ (
    .A(1'h1),
    .B(_3837_),
    .C(_4190_),
    .Y(_4191_)
);

OAI21X1 _10851_ (
    .A(1'h1),
    .B(_4190_),
    .C(_4191_),
    .Y(_4192_)
);

NAND2X1 _10852_ (
    .A(\genblk1[4].u_ce.Ain1 [0]),
    .B(_4192_),
    .Y(_4193_)
);

OR2X2 _10853_ (
    .A(_4192_),
    .B(\genblk1[4].u_ce.Ain1 [0]),
    .Y(_4194_)
);

NAND2X1 _10854_ (
    .A(_4193_),
    .B(_4194_),
    .Y(_4195_)
);

INVX1 _10855_ (
    .A(_4195_),
    .Y(_4196_)
);

NOR2X1 _10856_ (
    .A(_4196_),
    .B(_4189_),
    .Y(_4197_)
);

NAND2X1 _10857_ (
    .A(_4196_),
    .B(_4189_),
    .Y(_4198_)
);

NAND2X1 _10858_ (
    .A(\genblk1[4].u_ce.Vld_bF$buf4 ),
    .B(_4198_),
    .Y(_4199_)
);

OAI21X1 _10859_ (
    .A(_4197_),
    .B(_4199_),
    .C(_4188_),
    .Y(_3492_)
);

NAND2X1 _10860_ (
    .A(_4193_),
    .B(_4198_),
    .Y(_4200_)
);

INVX1 _10861_ (
    .A(_4200_),
    .Y(_4201_)
);

INVX1 _10862_ (
    .A(\genblk1[4].u_ce.Ain1 [1]),
    .Y(_4202_)
);

OAI21X1 _10863_ (
    .A(1'h0),
    .B(_3628__bF$buf2),
    .C(1'h1),
    .Y(_4203_)
);

NAND2X1 _10864_ (
    .A(_3717__bF$buf0),
    .B(_4203_),
    .Y(_4204_)
);

OAI21X1 _10865_ (
    .A(1'h1),
    .B(1'h0),
    .C(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .Y(_4205_)
);

OAI21X1 _10866_ (
    .A(_3624_),
    .B(_4205_),
    .C(_4204_),
    .Y(_4206_)
);

NOR2X1 _10867_ (
    .A(_4202_),
    .B(_4206_),
    .Y(_4207_)
);

NAND2X1 _10868_ (
    .A(_4202_),
    .B(_4206_),
    .Y(_4208_)
);

INVX1 _10869_ (
    .A(_4208_),
    .Y(_4209_)
);

OAI21X1 _10870_ (
    .A(_4207_),
    .B(_4209_),
    .C(_4201_),
    .Y(_4210_)
);

INVX1 _10871_ (
    .A(_4207_),
    .Y(_4211_)
);

NAND3X1 _10872_ (
    .A(_4211_),
    .B(_4208_),
    .C(_4200_),
    .Y(_4212_)
);

NAND2X1 _10873_ (
    .A(_4212_),
    .B(_4210_),
    .Y(_4213_)
);

NAND2X1 _10874_ (
    .A(\genblk1[4].u_ce.Acalc [3]),
    .B(_3622__bF$buf1),
    .Y(_4214_)
);

OAI21X1 _10875_ (
    .A(_3622__bF$buf0),
    .B(_4213_),
    .C(_4214_),
    .Y(_3493_)
);

NOR2X1 _10876_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf1 ),
    .B(_4179_),
    .Y(_4215_)
);

NAND3X1 _10877_ (
    .A(1'h0),
    .B(_3655__bF$buf1),
    .C(_3628__bF$buf1),
    .Y(_4216_)
);

AOI21X1 _10878_ (
    .A(_4178_),
    .B(_4216_),
    .C(_3717__bF$buf5),
    .Y(_4217_)
);

NOR2X1 _10879_ (
    .A(_4217_),
    .B(_4215_),
    .Y(_4218_)
);

NAND2X1 _10880_ (
    .A(\genblk1[4].u_ce.Ain12b [4]),
    .B(_4218_),
    .Y(_4219_)
);

INVX1 _10881_ (
    .A(\genblk1[4].u_ce.Ain12b [4]),
    .Y(_4220_)
);

OAI21X1 _10882_ (
    .A(_4217_),
    .B(_4215_),
    .C(_4220_),
    .Y(_4221_)
);

NAND2X1 _10883_ (
    .A(_4221_),
    .B(_4219_),
    .Y(_4222_)
);

AOI21X1 _10884_ (
    .A(_4200_),
    .B(_4208_),
    .C(_4207_),
    .Y(_4223_)
);

AND2X2 _10885_ (
    .A(_4223_),
    .B(_4222_),
    .Y(_4224_)
);

OAI21X1 _10886_ (
    .A(_4222_),
    .B(_4223_),
    .C(\genblk1[4].u_ce.Vld_bF$buf3 ),
    .Y(_4225_)
);

OAI22X1 _10887_ (
    .A(_3561_),
    .B(\genblk1[4].u_ce.Vld_bF$buf2 ),
    .C(_4225_),
    .D(_4224_),
    .Y(_3494_)
);

NAND2X1 _10888_ (
    .A(\genblk1[4].u_ce.Acalc [5]),
    .B(_3622__bF$buf4),
    .Y(_4226_)
);

OAI21X1 _10889_ (
    .A(_4222_),
    .B(_4223_),
    .C(_4219_),
    .Y(_4227_)
);

OAI21X1 _10890_ (
    .A(1'h0),
    .B(1'h0),
    .C(_3656_),
    .Y(_4228_)
);

NAND2X1 _10891_ (
    .A(_3717__bF$buf4),
    .B(_4228_),
    .Y(_4229_)
);

INVX1 _10892_ (
    .A(_4229_),
    .Y(_4230_)
);

NOR2X1 _10893_ (
    .A(_3717__bF$buf3),
    .B(_4228_),
    .Y(_4231_)
);

NOR2X1 _10894_ (
    .A(_4231_),
    .B(_4230_),
    .Y(_4232_)
);

NAND2X1 _10895_ (
    .A(\genblk1[4].u_ce.Ain12b [5]),
    .B(_4232_),
    .Y(_4233_)
);

INVX1 _10896_ (
    .A(\genblk1[4].u_ce.Ain12b [5]),
    .Y(_4234_)
);

OAI21X1 _10897_ (
    .A(_4231_),
    .B(_4230_),
    .C(_4234_),
    .Y(_4235_)
);

NAND2X1 _10898_ (
    .A(_4235_),
    .B(_4233_),
    .Y(_4236_)
);

INVX1 _10899_ (
    .A(_4236_),
    .Y(_4237_)
);

NOR2X1 _10900_ (
    .A(_4237_),
    .B(_4227_),
    .Y(_4238_)
);

NAND2X1 _10901_ (
    .A(_4237_),
    .B(_4227_),
    .Y(_4239_)
);

NAND2X1 _10902_ (
    .A(\genblk1[4].u_ce.Vld_bF$buf1 ),
    .B(_4239_),
    .Y(_4240_)
);

OAI21X1 _10903_ (
    .A(_4238_),
    .B(_4240_),
    .C(_4226_),
    .Y(_3495_)
);

NAND2X1 _10904_ (
    .A(\genblk1[4].u_ce.Acalc [6]),
    .B(_3622__bF$buf3),
    .Y(_4241_)
);

INVX1 _10905_ (
    .A(_4223_),
    .Y(_4242_)
);

NOR2X1 _10906_ (
    .A(_4222_),
    .B(_4236_),
    .Y(_4243_)
);

OAI21X1 _10907_ (
    .A(_4219_),
    .B(_4236_),
    .C(_4233_),
    .Y(_4244_)
);

AOI21X1 _10908_ (
    .A(_4242_),
    .B(_4243_),
    .C(_4244_),
    .Y(_4245_)
);

OAI21X1 _10909_ (
    .A(1'h1),
    .B(_4171_),
    .C(_3626_),
    .Y(_4246_)
);

NOR2X1 _10910_ (
    .A(_3717__bF$buf2),
    .B(_4246_),
    .Y(_4247_)
);

NAND2X1 _10911_ (
    .A(_3717__bF$buf1),
    .B(_4246_),
    .Y(_4248_)
);

INVX1 _10912_ (
    .A(_4248_),
    .Y(_4249_)
);

NOR2X1 _10913_ (
    .A(_4247_),
    .B(_4249_),
    .Y(_4250_)
);

NAND2X1 _10914_ (
    .A(\genblk1[4].u_ce.Ain12b [6]),
    .B(_4250_),
    .Y(_4251_)
);

OR2X2 _10915_ (
    .A(_4250_),
    .B(\genblk1[4].u_ce.Ain12b [6]),
    .Y(_4252_)
);

AND2X2 _10916_ (
    .A(_4252_),
    .B(_4251_),
    .Y(_4253_)
);

INVX1 _10917_ (
    .A(_4253_),
    .Y(_4254_)
);

AND2X2 _10918_ (
    .A(_4245_),
    .B(_4254_),
    .Y(_4255_)
);

OAI21X1 _10919_ (
    .A(_4254_),
    .B(_4245_),
    .C(\genblk1[4].u_ce.Vld_bF$buf0 ),
    .Y(_4256_)
);

OAI21X1 _10920_ (
    .A(_4256_),
    .B(_4255_),
    .C(_4241_),
    .Y(_3496_)
);

OAI21X1 _10921_ (
    .A(_4254_),
    .B(_4245_),
    .C(_4251_),
    .Y(_4257_)
);

OAI21X1 _10922_ (
    .A(1'h1),
    .B(1'h0),
    .C(\genblk1[4].u_ce.Ain12b_11_bF$buf0 ),
    .Y(_4258_)
);

NAND2X1 _10923_ (
    .A(_4258_),
    .B(_3718_),
    .Y(_4259_)
);

INVX1 _10924_ (
    .A(_4259_),
    .Y(_4260_)
);

NAND2X1 _10925_ (
    .A(\genblk1[4].u_ce.Ain12b [7]),
    .B(_4260_),
    .Y(_4261_)
);

INVX1 _10926_ (
    .A(_4261_),
    .Y(_4262_)
);

NOR2X1 _10927_ (
    .A(\genblk1[4].u_ce.Ain12b [7]),
    .B(_4260_),
    .Y(_4263_)
);

NOR2X1 _10928_ (
    .A(_4263_),
    .B(_4262_),
    .Y(_4264_)
);

INVX1 _10929_ (
    .A(_4264_),
    .Y(_4265_)
);

OR2X2 _10930_ (
    .A(_4257_),
    .B(_4265_),
    .Y(_4266_)
);

AOI21X1 _10931_ (
    .A(_4257_),
    .B(_4265_),
    .C(_3622__bF$buf2),
    .Y(_4267_)
);

AOI22X1 _10932_ (
    .A(_3575_),
    .B(_3622__bF$buf1),
    .C(_4266_),
    .D(_4267_),
    .Y(_3497_)
);

NAND2X1 _10933_ (
    .A(\genblk1[4].u_ce.Acalc [8]),
    .B(_3622__bF$buf0),
    .Y(_4268_)
);

OAI21X1 _10934_ (
    .A(_4263_),
    .B(_4251_),
    .C(_4261_),
    .Y(_4269_)
);

NAND2X1 _10935_ (
    .A(_4264_),
    .B(_4253_),
    .Y(_4270_)
);

INVX1 _10936_ (
    .A(_4270_),
    .Y(_4271_)
);

AOI21X1 _10937_ (
    .A(_4271_),
    .B(_4244_),
    .C(_4269_),
    .Y(_4272_)
);

NAND2X1 _10938_ (
    .A(_4243_),
    .B(_4271_),
    .Y(_4273_)
);

OAI21X1 _10939_ (
    .A(_4273_),
    .B(_4223_),
    .C(_4272_),
    .Y(_4274_)
);

INVX1 _10940_ (
    .A(\genblk1[4].u_ce.Ain12b [8]),
    .Y(_4275_)
);

NAND2X1 _10941_ (
    .A(_3717__bF$buf0),
    .B(_3625_),
    .Y(_4276_)
);

NAND2X1 _10942_ (
    .A(_4205_),
    .B(_4276_),
    .Y(_4277_)
);

OR2X2 _10943_ (
    .A(_4277_),
    .B(_4275_),
    .Y(_4278_)
);

NAND2X1 _10944_ (
    .A(_4275_),
    .B(_4277_),
    .Y(_4279_)
);

AND2X2 _10945_ (
    .A(_4278_),
    .B(_4279_),
    .Y(_4280_)
);

NOR2X1 _10946_ (
    .A(_4280_),
    .B(_4274_),
    .Y(_4281_)
);

NAND2X1 _10947_ (
    .A(_4280_),
    .B(_4274_),
    .Y(_4282_)
);

NAND2X1 _10948_ (
    .A(\genblk1[4].u_ce.Vld_bF$buf4 ),
    .B(_4282_),
    .Y(_4283_)
);

OAI21X1 _10949_ (
    .A(_4281_),
    .B(_4283_),
    .C(_4268_),
    .Y(_3498_)
);

NAND2X1 _10950_ (
    .A(\genblk1[4].u_ce.Acalc [9]),
    .B(_3622__bF$buf4),
    .Y(_4284_)
);

OAI21X1 _10951_ (
    .A(_4275_),
    .B(_4277_),
    .C(_4282_),
    .Y(_4285_)
);

INVX1 _10952_ (
    .A(\genblk1[4].u_ce.Ain12b [9]),
    .Y(_4286_)
);

NAND2X1 _10953_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf4 ),
    .B(_4286_),
    .Y(_4287_)
);

NOR2X1 _10954_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4286_),
    .Y(_4288_)
);

INVX1 _10955_ (
    .A(_4288_),
    .Y(_4289_)
);

NAND2X1 _10956_ (
    .A(_4287_),
    .B(_4289_),
    .Y(_4290_)
);

INVX1 _10957_ (
    .A(_4290_),
    .Y(_4291_)
);

NOR2X1 _10958_ (
    .A(_4291_),
    .B(_4285_),
    .Y(_4292_)
);

NAND2X1 _10959_ (
    .A(_4291_),
    .B(_4285_),
    .Y(_4293_)
);

NAND2X1 _10960_ (
    .A(\genblk1[4].u_ce.Vld_bF$buf3 ),
    .B(_4293_),
    .Y(_4294_)
);

OAI21X1 _10961_ (
    .A(_4292_),
    .B(_4294_),
    .C(_4284_),
    .Y(_3499_)
);

AOI21X1 _10962_ (
    .A(_4285_),
    .B(_4287_),
    .C(_4288_),
    .Y(_4295_)
);

INVX1 _10963_ (
    .A(\genblk1[4].u_ce.Ain12b [10]),
    .Y(_4296_)
);

NAND2X1 _10964_ (
    .A(\genblk1[4].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4296_),
    .Y(_4297_)
);

NAND2X1 _10965_ (
    .A(\genblk1[4].u_ce.Ain12b [10]),
    .B(_3717__bF$buf5),
    .Y(_4298_)
);

NAND2X1 _10966_ (
    .A(_4297_),
    .B(_4298_),
    .Y(_4299_)
);

AND2X2 _10967_ (
    .A(_4295_),
    .B(_4299_),
    .Y(_4300_)
);

OAI21X1 _10968_ (
    .A(_4299_),
    .B(_4295_),
    .C(\genblk1[4].u_ce.Vld_bF$buf2 ),
    .Y(_4301_)
);

OAI22X1 _10969_ (
    .A(_3557_),
    .B(\genblk1[4].u_ce.Vld_bF$buf1 ),
    .C(_4301_),
    .D(_4300_),
    .Y(_3500_)
);

NAND2X1 _10970_ (
    .A(\genblk1[4].u_ce.Acalc [11]),
    .B(_3622__bF$buf3),
    .Y(_4302_)
);

OAI21X1 _10971_ (
    .A(_4299_),
    .B(_4295_),
    .C(_4298_),
    .Y(_4303_)
);

OAI21X1 _10972_ (
    .A(_3622__bF$buf2),
    .B(_4303_),
    .C(_4302_),
    .Y(_3501_)
);

INVX1 _10973_ (
    .A(_3556_),
    .Y(_4304_)
);

NAND3X1 _10974_ (
    .A(_3609_),
    .B(\genblk1[4].u_ce.LoadCtl [5]),
    .C(_3567_),
    .Y(_4305_)
);

NOR2X1 _10975_ (
    .A(_4304_),
    .B(_4305_),
    .Y(_4306_)
);

NAND2X1 _10976_ (
    .A(\genblk1[3].u_ce.X_ [0]),
    .B(_4306_),
    .Y(_4307_)
);

OAI21X1 _10977_ (
    .A(_3751_),
    .B(_4306_),
    .C(_4307_),
    .Y(_3502_)
);

NAND2X1 _10978_ (
    .A(\genblk1[3].u_ce.X_ [1]),
    .B(_4306_),
    .Y(_4308_)
);

OAI21X1 _10979_ (
    .A(_3776_),
    .B(_4306_),
    .C(_4308_),
    .Y(_3503_)
);

INVX1 _10980_ (
    .A(\genblk1[3].u_ce.X_ [0]),
    .Y(_4309_)
);

NAND3X1 _10981_ (
    .A(\genblk1[4].u_ce.LoadCtl [4]),
    .B(_3556_),
    .C(_3567_),
    .Y(_4310_)
);

NAND2X1 _10982_ (
    .A(\genblk1[4].u_ce.Xin12b [8]),
    .B(_4310_),
    .Y(_4311_)
);

OAI21X1 _10983_ (
    .A(_4309_),
    .B(_4310_),
    .C(_4311_),
    .Y(_3504_)
);

INVX1 _10984_ (
    .A(\genblk1[3].u_ce.X_ [1]),
    .Y(_4312_)
);

NAND2X1 _10985_ (
    .A(\genblk1[4].u_ce.Xin12b [9]),
    .B(_4310_),
    .Y(_4313_)
);

OAI21X1 _10986_ (
    .A(_4312_),
    .B(_4310_),
    .C(_4313_),
    .Y(_3505_)
);

NAND2X1 _10987_ (
    .A(_3567_),
    .B(_3563_),
    .Y(_4314_)
);

OAI21X1 _10988_ (
    .A(_3568_),
    .B(_3576_),
    .C(\genblk1[4].u_ce.Xin12b [6]),
    .Y(_4315_)
);

OAI21X1 _10989_ (
    .A(_4309_),
    .B(_4314_),
    .C(_4315_),
    .Y(_3506_)
);

OAI21X1 _10990_ (
    .A(_3568_),
    .B(_3576_),
    .C(\genblk1[4].u_ce.Xin12b [7]),
    .Y(_4316_)
);

OAI21X1 _10991_ (
    .A(_4312_),
    .B(_4314_),
    .C(_4316_),
    .Y(_3507_)
);

NOR2X1 _10992_ (
    .A(_3560_),
    .B(_3568_),
    .Y(_4317_)
);

NAND2X1 _10993_ (
    .A(\genblk1[3].u_ce.X_ [0]),
    .B(_4317_),
    .Y(_4318_)
);

OAI21X1 _10994_ (
    .A(_3661_),
    .B(_4317_),
    .C(_4318_),
    .Y(_3508_)
);

NAND2X1 _10995_ (
    .A(\genblk1[3].u_ce.X_ [1]),
    .B(_4317_),
    .Y(_4319_)
);

OAI21X1 _10996_ (
    .A(_3669_),
    .B(_4317_),
    .C(_4319_),
    .Y(_3509_)
);

OAI21X1 _10997_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_3569_),
    .C(\genblk1[4].u_ce.Xin1 [0]),
    .Y(_4320_)
);

OAI21X1 _10998_ (
    .A(_4309_),
    .B(_3598_),
    .C(_4320_),
    .Y(_3510_)
);

OAI21X1 _10999_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_3569_),
    .C(\genblk1[4].u_ce.Xin1 [1]),
    .Y(_4321_)
);

OAI21X1 _11000_ (
    .A(_4312_),
    .B(_3598_),
    .C(_4321_),
    .Y(_3511_)
);

NAND2X1 _11001_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[3].u_ce.X_ [0]),
    .Y(_4322_)
);

OAI21X1 _11002_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_3684_),
    .C(_4322_),
    .Y(_3512_)
);

NAND2X1 _11003_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[3].u_ce.X_ [1]),
    .Y(_4323_)
);

OAI21X1 _11004_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_3664_),
    .C(_4323_),
    .Y(_3513_)
);

NAND2X1 _11005_ (
    .A(\genblk1[3].u_ce.Y_ [0]),
    .B(_4306_),
    .Y(_4324_)
);

OAI21X1 _11006_ (
    .A(_3884_),
    .B(_4306_),
    .C(_4324_),
    .Y(_3514_)
);

NAND2X1 _11007_ (
    .A(\genblk1[3].u_ce.Y_ [1]),
    .B(_4306_),
    .Y(_4325_)
);

OAI21X1 _11008_ (
    .A(_3908_),
    .B(_4306_),
    .C(_4325_),
    .Y(_3515_)
);

INVX1 _11009_ (
    .A(\genblk1[3].u_ce.Y_ [0]),
    .Y(_4326_)
);

NAND2X1 _11010_ (
    .A(\genblk1[4].u_ce.Yin12b [8]),
    .B(_4310_),
    .Y(_4327_)
);

OAI21X1 _11011_ (
    .A(_4326_),
    .B(_4310_),
    .C(_4327_),
    .Y(_3516_)
);

INVX1 _11012_ (
    .A(\genblk1[3].u_ce.Y_ [1]),
    .Y(_4328_)
);

NAND2X1 _11013_ (
    .A(\genblk1[4].u_ce.Yin12b [9]),
    .B(_4310_),
    .Y(_4329_)
);

OAI21X1 _11014_ (
    .A(_4328_),
    .B(_4310_),
    .C(_4329_),
    .Y(_3517_)
);

OAI21X1 _11015_ (
    .A(_3568_),
    .B(_3576_),
    .C(\genblk1[4].u_ce.Yin12b [6]),
    .Y(_3536_)
);

OAI21X1 _11016_ (
    .A(_4326_),
    .B(_4314_),
    .C(_3536_),
    .Y(_3518_)
);

OAI21X1 _11017_ (
    .A(_3568_),
    .B(_3576_),
    .C(\genblk1[4].u_ce.Yin12b [7]),
    .Y(_3537_)
);

OAI21X1 _11018_ (
    .A(_4328_),
    .B(_4314_),
    .C(_3537_),
    .Y(_3519_)
);

NAND2X1 _11019_ (
    .A(\genblk1[3].u_ce.Y_ [0]),
    .B(_4317_),
    .Y(_3538_)
);

OAI21X1 _11020_ (
    .A(_3749_),
    .B(_4317_),
    .C(_3538_),
    .Y(_3520_)
);

NAND2X1 _11021_ (
    .A(\genblk1[3].u_ce.Y_ [1]),
    .B(_4317_),
    .Y(_3539_)
);

OAI21X1 _11022_ (
    .A(_3774_),
    .B(_4317_),
    .C(_3539_),
    .Y(_3521_)
);

OAI21X1 _11023_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_3569_),
    .C(\genblk1[4].u_ce.Yin1 [0]),
    .Y(_3540_)
);

OAI21X1 _11024_ (
    .A(_4326_),
    .B(_3598_),
    .C(_3540_),
    .Y(_3522_)
);

OAI21X1 _11025_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_3569_),
    .C(\genblk1[4].u_ce.Yin1 [1]),
    .Y(_3541_)
);

OAI21X1 _11026_ (
    .A(_4328_),
    .B(_3598_),
    .C(_3541_),
    .Y(_3523_)
);

NAND2X1 _11027_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[3].u_ce.Y_ [0]),
    .Y(_3542_)
);

OAI21X1 _11028_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_3921_),
    .C(_3542_),
    .Y(_3524_)
);

NAND2X1 _11029_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[3].u_ce.Y_ [1]),
    .Y(_3543_)
);

OAI21X1 _11030_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_3706_),
    .C(_3543_),
    .Y(_3525_)
);

NAND2X1 _11031_ (
    .A(\a[4] [0]),
    .B(_4306_),
    .Y(_3544_)
);

OAI21X1 _11032_ (
    .A(_4296_),
    .B(_4306_),
    .C(_3544_),
    .Y(_3526_)
);

NAND2X1 _11033_ (
    .A(\a[4] [1]),
    .B(_4306_),
    .Y(_3545_)
);

OAI21X1 _11034_ (
    .A(_3717__bF$buf4),
    .B(_4306_),
    .C(_3545_),
    .Y(_3527_)
);

INVX1 _11035_ (
    .A(\a[4] [0]),
    .Y(_3546_)
);

NAND2X1 _11036_ (
    .A(\genblk1[4].u_ce.Ain12b [8]),
    .B(_4310_),
    .Y(_3547_)
);

OAI21X1 _11037_ (
    .A(_3546_),
    .B(_4310_),
    .C(_3547_),
    .Y(_3528_)
);

INVX1 _11038_ (
    .A(\a[4] [1]),
    .Y(_3548_)
);

NAND2X1 _11039_ (
    .A(\genblk1[4].u_ce.Ain12b [9]),
    .B(_4310_),
    .Y(_3549_)
);

OAI21X1 _11040_ (
    .A(_3548_),
    .B(_4310_),
    .C(_3549_),
    .Y(_3529_)
);

OAI21X1 _11041_ (
    .A(_3568_),
    .B(_3576_),
    .C(\genblk1[4].u_ce.Ain12b [6]),
    .Y(_3550_)
);

OAI21X1 _11042_ (
    .A(_3546_),
    .B(_4314_),
    .C(_3550_),
    .Y(_3530_)
);

OAI21X1 _11043_ (
    .A(_3568_),
    .B(_3576_),
    .C(\genblk1[4].u_ce.Ain12b [7]),
    .Y(_3551_)
);

OAI21X1 _11044_ (
    .A(_3548_),
    .B(_4314_),
    .C(_3551_),
    .Y(_3531_)
);

NAND2X1 _11045_ (
    .A(\a[4] [0]),
    .B(_4317_),
    .Y(_3552_)
);

OAI21X1 _11046_ (
    .A(_4220_),
    .B(_4317_),
    .C(_3552_),
    .Y(_3532_)
);

NAND2X1 _11047_ (
    .A(\a[4] [1]),
    .B(_4317_),
    .Y(_3553_)
);

OAI21X1 _11048_ (
    .A(_4234_),
    .B(_4317_),
    .C(_3553_),
    .Y(_3533_)
);

OAI21X1 _11049_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_3569_),
    .C(\genblk1[4].u_ce.Ain1 [0]),
    .Y(_3554_)
);

OAI21X1 _11050_ (
    .A(_3546_),
    .B(_3598_),
    .C(_3554_),
    .Y(_3534_)
);

OAI21X1 _11051_ (
    .A(\genblk1[4].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_3569_),
    .C(\genblk1[4].u_ce.Ain1 [1]),
    .Y(_3555_)
);

OAI21X1 _11052_ (
    .A(_3548_),
    .B(_3598_),
    .C(_3555_),
    .Y(_3535_)
);

DFFPOSX1 _11053_ (
    .CLK(clk_bF$buf65),
    .D(_3464_),
    .Q(\genblk1[4].u_ce.Ain0 [0])
);

DFFPOSX1 _11054_ (
    .CLK(clk_bF$buf64),
    .D(_3465_),
    .Q(\genblk1[4].u_ce.Ain0 [1])
);

DFFPOSX1 _11055_ (
    .CLK(clk_bF$buf63),
    .D(_3466_),
    .Q(\genblk1[4].u_ce.Ycalc [2])
);

DFFPOSX1 _11056_ (
    .CLK(clk_bF$buf62),
    .D(_3467_),
    .Q(\genblk1[4].u_ce.Ycalc [3])
);

DFFPOSX1 _11057_ (
    .CLK(clk_bF$buf61),
    .D(_3468_),
    .Q(\genblk1[4].u_ce.Ycalc [4])
);

DFFPOSX1 _11058_ (
    .CLK(clk_bF$buf60),
    .D(_3469_),
    .Q(\genblk1[4].u_ce.Ycalc [5])
);

DFFPOSX1 _11059_ (
    .CLK(clk_bF$buf59),
    .D(_3470_),
    .Q(\genblk1[4].u_ce.Ycalc [6])
);

DFFPOSX1 _11060_ (
    .CLK(clk_bF$buf58),
    .D(_3471_),
    .Q(\genblk1[4].u_ce.Ycalc [7])
);

DFFPOSX1 _11061_ (
    .CLK(clk_bF$buf57),
    .D(_3472_),
    .Q(\genblk1[4].u_ce.Ycalc [8])
);

DFFPOSX1 _11062_ (
    .CLK(clk_bF$buf56),
    .D(_3473_),
    .Q(\genblk1[4].u_ce.Ycalc [9])
);

DFFPOSX1 _11063_ (
    .CLK(clk_bF$buf55),
    .D(_3474_),
    .Q(\genblk1[4].u_ce.Ycalc [10])
);

DFFPOSX1 _11064_ (
    .CLK(clk_bF$buf54),
    .D(_3475_),
    .Q(\genblk1[4].u_ce.Ycalc [11])
);

DFFPOSX1 _11065_ (
    .CLK(clk_bF$buf53),
    .D(_3476_),
    .Q(\genblk1[4].u_ce.Ycalc [0])
);

DFFPOSX1 _11066_ (
    .CLK(clk_bF$buf52),
    .D(_3477_),
    .Q(\genblk1[4].u_ce.Ycalc [1])
);

DFFPOSX1 _11067_ (
    .CLK(clk_bF$buf51),
    .D(_3478_),
    .Q(\genblk1[4].u_ce.Xcalc [0])
);

DFFPOSX1 _11068_ (
    .CLK(clk_bF$buf50),
    .D(_3479_),
    .Q(\genblk1[4].u_ce.Xcalc [1])
);

DFFPOSX1 _11069_ (
    .CLK(clk_bF$buf49),
    .D(_3480_),
    .Q(\genblk1[4].u_ce.Xcalc [2])
);

DFFPOSX1 _11070_ (
    .CLK(clk_bF$buf48),
    .D(_3481_),
    .Q(\genblk1[4].u_ce.Xcalc [3])
);

DFFPOSX1 _11071_ (
    .CLK(clk_bF$buf47),
    .D(_3482_),
    .Q(\genblk1[4].u_ce.Xcalc [4])
);

DFFPOSX1 _11072_ (
    .CLK(clk_bF$buf46),
    .D(_3483_),
    .Q(\genblk1[4].u_ce.Xcalc [5])
);

DFFPOSX1 _11073_ (
    .CLK(clk_bF$buf45),
    .D(_3484_),
    .Q(\genblk1[4].u_ce.Xcalc [6])
);

DFFPOSX1 _11074_ (
    .CLK(clk_bF$buf44),
    .D(_3485_),
    .Q(\genblk1[4].u_ce.Xcalc [7])
);

DFFPOSX1 _11075_ (
    .CLK(clk_bF$buf43),
    .D(_3486_),
    .Q(\genblk1[4].u_ce.Xcalc [8])
);

DFFPOSX1 _11076_ (
    .CLK(clk_bF$buf42),
    .D(_3487_),
    .Q(\genblk1[4].u_ce.Xcalc [9])
);

DFFPOSX1 _11077_ (
    .CLK(clk_bF$buf41),
    .D(_3488_),
    .Q(\genblk1[4].u_ce.Xcalc [10])
);

DFFPOSX1 _11078_ (
    .CLK(clk_bF$buf40),
    .D(_3489_),
    .Q(\genblk1[4].u_ce.Xcalc [11])
);

DFFPOSX1 _11079_ (
    .CLK(clk_bF$buf39),
    .D(_3490_),
    .Q(\genblk1[4].u_ce.Acalc [0])
);

DFFPOSX1 _11080_ (
    .CLK(clk_bF$buf38),
    .D(_3491_),
    .Q(\genblk1[4].u_ce.Acalc [1])
);

DFFPOSX1 _11081_ (
    .CLK(clk_bF$buf37),
    .D(_3492_),
    .Q(\genblk1[4].u_ce.Acalc [2])
);

DFFPOSX1 _11082_ (
    .CLK(clk_bF$buf36),
    .D(_3493_),
    .Q(\genblk1[4].u_ce.Acalc [3])
);

DFFPOSX1 _11083_ (
    .CLK(clk_bF$buf35),
    .D(_3494_),
    .Q(\genblk1[4].u_ce.Acalc [4])
);

DFFPOSX1 _11084_ (
    .CLK(clk_bF$buf34),
    .D(_3495_),
    .Q(\genblk1[4].u_ce.Acalc [5])
);

DFFPOSX1 _11085_ (
    .CLK(clk_bF$buf33),
    .D(_3496_),
    .Q(\genblk1[4].u_ce.Acalc [6])
);

DFFPOSX1 _11086_ (
    .CLK(clk_bF$buf32),
    .D(_3497_),
    .Q(\genblk1[4].u_ce.Acalc [7])
);

DFFPOSX1 _11087_ (
    .CLK(clk_bF$buf31),
    .D(_3498_),
    .Q(\genblk1[4].u_ce.Acalc [8])
);

DFFPOSX1 _11088_ (
    .CLK(clk_bF$buf30),
    .D(_3499_),
    .Q(\genblk1[4].u_ce.Acalc [9])
);

DFFPOSX1 _11089_ (
    .CLK(clk_bF$buf29),
    .D(_3500_),
    .Q(\genblk1[4].u_ce.Acalc [10])
);

DFFPOSX1 _11090_ (
    .CLK(clk_bF$buf28),
    .D(_3501_),
    .Q(\genblk1[4].u_ce.Acalc [11])
);

DFFPOSX1 _11091_ (
    .CLK(clk_bF$buf27),
    .D(_3502_),
    .Q(\genblk1[4].u_ce.Xin12b [10])
);

DFFPOSX1 _11092_ (
    .CLK(clk_bF$buf26),
    .D(_3503_),
    .Q(\genblk1[4].u_ce.Xin12b [11])
);

DFFPOSX1 _11093_ (
    .CLK(clk_bF$buf25),
    .D(_3504_),
    .Q(\genblk1[4].u_ce.Xin12b [8])
);

DFFPOSX1 _11094_ (
    .CLK(clk_bF$buf24),
    .D(_3505_),
    .Q(\genblk1[4].u_ce.Xin12b [9])
);

DFFPOSX1 _11095_ (
    .CLK(clk_bF$buf23),
    .D(_3506_),
    .Q(\genblk1[4].u_ce.Xin12b [6])
);

DFFPOSX1 _11096_ (
    .CLK(clk_bF$buf22),
    .D(_3507_),
    .Q(\genblk1[4].u_ce.Xin12b [7])
);

DFFPOSX1 _11097_ (
    .CLK(clk_bF$buf21),
    .D(_3508_),
    .Q(\genblk1[4].u_ce.Xin12b [4])
);

DFFPOSX1 _11098_ (
    .CLK(clk_bF$buf20),
    .D(_3509_),
    .Q(\genblk1[4].u_ce.Xin12b [5])
);

DFFPOSX1 _11099_ (
    .CLK(clk_bF$buf19),
    .D(_3510_),
    .Q(\genblk1[4].u_ce.Xin1 [0])
);

DFFPOSX1 _11100_ (
    .CLK(clk_bF$buf18),
    .D(_3511_),
    .Q(\genblk1[4].u_ce.Xin1 [1])
);

DFFPOSX1 _11101_ (
    .CLK(clk_bF$buf17),
    .D(_3512_),
    .Q(\genblk1[4].u_ce.Xin0 [0])
);

DFFPOSX1 _11102_ (
    .CLK(clk_bF$buf16),
    .D(_3513_),
    .Q(\genblk1[4].u_ce.Xin0 [1])
);

DFFPOSX1 _11103_ (
    .CLK(clk_bF$buf15),
    .D(_3514_),
    .Q(\genblk1[4].u_ce.Yin12b [10])
);

DFFPOSX1 _11104_ (
    .CLK(clk_bF$buf14),
    .D(_3515_),
    .Q(\genblk1[4].u_ce.Yin12b [11])
);

DFFPOSX1 _11105_ (
    .CLK(clk_bF$buf13),
    .D(_3516_),
    .Q(\genblk1[4].u_ce.Yin12b [8])
);

DFFPOSX1 _11106_ (
    .CLK(clk_bF$buf12),
    .D(_3517_),
    .Q(\genblk1[4].u_ce.Yin12b [9])
);

DFFPOSX1 _11107_ (
    .CLK(clk_bF$buf11),
    .D(_3518_),
    .Q(\genblk1[4].u_ce.Yin12b [6])
);

DFFPOSX1 _11108_ (
    .CLK(clk_bF$buf10),
    .D(_3519_),
    .Q(\genblk1[4].u_ce.Yin12b [7])
);

DFFPOSX1 _11109_ (
    .CLK(clk_bF$buf9),
    .D(_3520_),
    .Q(\genblk1[4].u_ce.Yin12b [4])
);

DFFPOSX1 _11110_ (
    .CLK(clk_bF$buf8),
    .D(_3521_),
    .Q(\genblk1[4].u_ce.Yin12b [5])
);

DFFPOSX1 _11111_ (
    .CLK(clk_bF$buf7),
    .D(_3522_),
    .Q(\genblk1[4].u_ce.Yin1 [0])
);

DFFPOSX1 _11112_ (
    .CLK(clk_bF$buf6),
    .D(_3523_),
    .Q(\genblk1[4].u_ce.Yin1 [1])
);

DFFPOSX1 _11113_ (
    .CLK(clk_bF$buf5),
    .D(_3524_),
    .Q(\genblk1[4].u_ce.Yin0 [0])
);

DFFPOSX1 _11114_ (
    .CLK(clk_bF$buf4),
    .D(_3525_),
    .Q(\genblk1[4].u_ce.Yin0 [1])
);

DFFPOSX1 _11115_ (
    .CLK(clk_bF$buf3),
    .D(_3526_),
    .Q(\genblk1[4].u_ce.Ain12b [10])
);

DFFPOSX1 _11116_ (
    .CLK(clk_bF$buf2),
    .D(_3527_),
    .Q(\genblk1[4].u_ce.Ain12b [11])
);

DFFPOSX1 _11117_ (
    .CLK(clk_bF$buf1),
    .D(_3528_),
    .Q(\genblk1[4].u_ce.Ain12b [8])
);

DFFPOSX1 _11118_ (
    .CLK(clk_bF$buf0),
    .D(_3529_),
    .Q(\genblk1[4].u_ce.Ain12b [9])
);

DFFPOSX1 _11119_ (
    .CLK(clk_bF$buf75),
    .D(_3530_),
    .Q(\genblk1[4].u_ce.Ain12b [6])
);

DFFPOSX1 _11120_ (
    .CLK(clk_bF$buf74),
    .D(_3531_),
    .Q(\genblk1[4].u_ce.Ain12b [7])
);

DFFPOSX1 _11121_ (
    .CLK(clk_bF$buf73),
    .D(_3532_),
    .Q(\genblk1[4].u_ce.Ain12b [4])
);

DFFPOSX1 _11122_ (
    .CLK(clk_bF$buf72),
    .D(_3533_),
    .Q(\genblk1[4].u_ce.Ain12b [5])
);

DFFPOSX1 _11123_ (
    .CLK(clk_bF$buf71),
    .D(_3534_),
    .Q(\genblk1[4].u_ce.Ain1 [0])
);

DFFPOSX1 _11124_ (
    .CLK(clk_bF$buf70),
    .D(_3535_),
    .Q(\genblk1[4].u_ce.Ain1 [1])
);

DFFPOSX1 _11125_ (
    .CLK(clk_bF$buf69),
    .D(\genblk1[3].u_ce.ISout ),
    .Q(\genblk1[4].u_ce.ISpipe [0])
);

DFFPOSX1 _11126_ (
    .CLK(clk_bF$buf68),
    .D(\genblk1[4].u_ce.ISpipe [0]),
    .Q(\genblk1[4].u_ce.ISpipe [1])
);

DFFPOSX1 _11127_ (
    .CLK(clk_bF$buf67),
    .D(\genblk1[4].u_ce.ISpipe [1]),
    .Q(\genblk1[4].u_ce.ISpipe [2])
);

DFFPOSX1 _11128_ (
    .CLK(clk_bF$buf66),
    .D(\genblk1[4].u_ce.ISpipe [2]),
    .Q(\genblk1[4].u_ce.ISpipe [3])
);

DFFPOSX1 _11129_ (
    .CLK(clk_bF$buf65),
    .D(\genblk1[4].u_ce.ISpipe [3]),
    .Q(\genblk1[4].u_ce.ISpipe [4])
);

DFFPOSX1 _11130_ (
    .CLK(clk_bF$buf64),
    .D(\genblk1[4].u_ce.ISpipe [4]),
    .Q(\genblk1[4].u_ce.ISpipe [5])
);

DFFPOSX1 _11131_ (
    .CLK(clk_bF$buf63),
    .D(\genblk1[4].u_ce.ISpipe [5]),
    .Q(\genblk1[4].u_ce.ISout )
);

DFFPOSX1 _11132_ (
    .CLK(clk_bF$buf62),
    .D(\genblk1[3].u_ce.Vld_bF$buf1 ),
    .Q(\genblk1[4].u_ce.LoadCtl [0])
);

DFFPOSX1 _11133_ (
    .CLK(clk_bF$buf61),
    .D(\genblk1[4].u_ce.LoadCtl_0_bF$buf3 ),
    .Q(\genblk1[4].u_ce.LoadCtl [1])
);

DFFPOSX1 _11134_ (
    .CLK(clk_bF$buf60),
    .D(\genblk1[4].u_ce.LoadCtl [1]),
    .Q(\genblk1[4].u_ce.LoadCtl [2])
);

DFFPOSX1 _11135_ (
    .CLK(clk_bF$buf59),
    .D(\genblk1[4].u_ce.LoadCtl [2]),
    .Q(\genblk1[4].u_ce.LoadCtl [3])
);

DFFPOSX1 _11136_ (
    .CLK(clk_bF$buf58),
    .D(\genblk1[4].u_ce.LoadCtl [3]),
    .Q(\genblk1[4].u_ce.LoadCtl [4])
);

DFFPOSX1 _11137_ (
    .CLK(clk_bF$buf57),
    .D(\genblk1[4].u_ce.LoadCtl [4]),
    .Q(\genblk1[4].u_ce.LoadCtl [5])
);

DFFPOSX1 _11138_ (
    .CLK(clk_bF$buf56),
    .D(\genblk1[4].u_ce.LoadCtl [5]),
    .Q(\genblk1[4].u_ce.Vld )
);

NOR2X1 _11139_ (
    .A(\genblk1[5].u_ce.LoadCtl [3]),
    .B(\genblk1[5].u_ce.LoadCtl [2]),
    .Y(_4416_)
);

INVX2 _11140_ (
    .A(\genblk1[5].u_ce.LoadCtl [2]),
    .Y(_4417_)
);

INVX1 _11141_ (
    .A(\genblk1[5].u_ce.LoadCtl [3]),
    .Y(_4418_)
);

NOR2X1 _11142_ (
    .A(\genblk1[5].u_ce.LoadCtl [2]),
    .B(_4418_),
    .Y(_4419_)
);

NOR2X1 _11143_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[5].u_ce.LoadCtl [1]),
    .Y(_4420_)
);

INVX4 _11144_ (
    .A(_4420_),
    .Y(_4421_)
);

INVX2 _11145_ (
    .A(\genblk1[5].u_ce.LoadCtl [1]),
    .Y(_4422_)
);

NOR2X1 _11146_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_4422_),
    .Y(_4423_)
);

INVX1 _11147_ (
    .A(\genblk1[5].u_ce.Acalc [11]),
    .Y(_4424_)
);

NAND2X1 _11148_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(\genblk1[5].u_ce.Acalc [9]),
    .Y(_4425_)
);

OAI21X1 _11149_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(_4424_),
    .C(_4425_),
    .Y(_4426_)
);

INVX1 _11150_ (
    .A(\genblk1[5].u_ce.Acalc [7]),
    .Y(_4427_)
);

INVX4 _11151_ (
    .A(_4419_),
    .Y(_4428_)
);

NAND2X1 _11152_ (
    .A(\genblk1[5].u_ce.LoadCtl [2]),
    .B(\genblk1[5].u_ce.Acalc [5]),
    .Y(_4429_)
);

OAI21X1 _11153_ (
    .A(_4427_),
    .B(_4428_),
    .C(_4429_),
    .Y(_4430_)
);

AOI21X1 _11154_ (
    .A(_4416_),
    .B(_4426_),
    .C(_4430_),
    .Y(_4431_)
);

AOI22X1 _11155_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[5].u_ce.Acalc [1]),
    .C(_4423_),
    .D(\genblk1[5].u_ce.Acalc [3]),
    .Y(_4432_)
);

OAI21X1 _11156_ (
    .A(_4421_),
    .B(_4431_),
    .C(_4432_),
    .Y(\a[6] [1])
);

INVX1 _11157_ (
    .A(\genblk1[5].u_ce.Ycalc [10]),
    .Y(_4433_)
);

NAND2X1 _11158_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(\genblk1[5].u_ce.Ycalc [8]),
    .Y(_4434_)
);

OAI21X1 _11159_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(_4433_),
    .C(_4434_),
    .Y(_4435_)
);

INVX1 _11160_ (
    .A(\genblk1[5].u_ce.Ycalc [6]),
    .Y(_4436_)
);

INVX1 _11161_ (
    .A(\genblk1[5].u_ce.Ycalc [4]),
    .Y(_4437_)
);

OAI22X1 _11162_ (
    .A(_4417_),
    .B(_4437_),
    .C(_4436_),
    .D(_4428_),
    .Y(_4438_)
);

AOI21X1 _11163_ (
    .A(_4416_),
    .B(_4435_),
    .C(_4438_),
    .Y(_4439_)
);

AOI22X1 _11164_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[5].u_ce.Ycalc [0]),
    .C(_4423_),
    .D(\genblk1[5].u_ce.Ycalc [2]),
    .Y(_4440_)
);

OAI21X1 _11165_ (
    .A(_4421_),
    .B(_4439_),
    .C(_4440_),
    .Y(\genblk1[5].u_ce.Y_ [0])
);

INVX1 _11166_ (
    .A(\genblk1[5].u_ce.Ycalc [11]),
    .Y(_4441_)
);

NAND2X1 _11167_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(\genblk1[5].u_ce.Ycalc [9]),
    .Y(_4442_)
);

OAI21X1 _11168_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(_4441_),
    .C(_4442_),
    .Y(_4443_)
);

INVX1 _11169_ (
    .A(\genblk1[5].u_ce.Ycalc [7]),
    .Y(_4444_)
);

INVX1 _11170_ (
    .A(\genblk1[5].u_ce.Ycalc [5]),
    .Y(_4445_)
);

OAI22X1 _11171_ (
    .A(_4417_),
    .B(_4445_),
    .C(_4444_),
    .D(_4428_),
    .Y(_4446_)
);

AOI21X1 _11172_ (
    .A(_4416_),
    .B(_4443_),
    .C(_4446_),
    .Y(_4447_)
);

AOI22X1 _11173_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[5].u_ce.Ycalc [1]),
    .C(_4423_),
    .D(\genblk1[5].u_ce.Ycalc [3]),
    .Y(_4448_)
);

OAI21X1 _11174_ (
    .A(_4421_),
    .B(_4447_),
    .C(_4448_),
    .Y(\genblk1[5].u_ce.Y_ [1])
);

INVX1 _11175_ (
    .A(\genblk1[5].u_ce.Xcalc [2]),
    .Y(_4449_)
);

INVX2 _11176_ (
    .A(_4423_),
    .Y(_4450_)
);

INVX1 _11177_ (
    .A(\genblk1[5].u_ce.Xcalc [4]),
    .Y(_4451_)
);

INVX1 _11178_ (
    .A(\genblk1[5].u_ce.Xcalc [6]),
    .Y(_4452_)
);

NOR2X1 _11179_ (
    .A(_4418_),
    .B(_4452_),
    .Y(_4453_)
);

INVX1 _11180_ (
    .A(\genblk1[5].u_ce.Xcalc [8]),
    .Y(_4454_)
);

NAND2X1 _11181_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(_4454_),
    .Y(_4455_)
);

OAI21X1 _11182_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(\genblk1[5].u_ce.Xcalc [10]),
    .C(_4455_),
    .Y(_4456_)
);

NOR2X1 _11183_ (
    .A(\genblk1[5].u_ce.LoadCtl [3]),
    .B(_4456_),
    .Y(_4457_)
);

OAI21X1 _11184_ (
    .A(_4453_),
    .B(_4457_),
    .C(_4417_),
    .Y(_4458_)
);

OAI21X1 _11185_ (
    .A(_4417_),
    .B(_4451_),
    .C(_4458_),
    .Y(_4459_)
);

AOI22X1 _11186_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[5].u_ce.Xcalc [0]),
    .C(_4459_),
    .D(_4420_),
    .Y(_4460_)
);

OAI21X1 _11187_ (
    .A(_4449_),
    .B(_4450_),
    .C(_4460_),
    .Y(\genblk1[5].u_ce.X_ [0])
);

INVX1 _11188_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .Y(_4461_)
);

INVX1 _11189_ (
    .A(\genblk1[5].u_ce.Xcalc [9]),
    .Y(_4462_)
);

NAND2X1 _11190_ (
    .A(\genblk1[5].u_ce.Xcalc [11]),
    .B(_4461_),
    .Y(_4463_)
);

OAI21X1 _11191_ (
    .A(_4461_),
    .B(_4462_),
    .C(_4463_),
    .Y(_4464_)
);

INVX1 _11192_ (
    .A(\genblk1[5].u_ce.Xcalc [7]),
    .Y(_4465_)
);

INVX1 _11193_ (
    .A(\genblk1[5].u_ce.Xcalc [5]),
    .Y(_4466_)
);

OAI22X1 _11194_ (
    .A(_4417_),
    .B(_4466_),
    .C(_4465_),
    .D(_4428_),
    .Y(_4467_)
);

AOI21X1 _11195_ (
    .A(_4416_),
    .B(_4464_),
    .C(_4467_),
    .Y(_4468_)
);

AOI22X1 _11196_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[5].u_ce.Xcalc [1]),
    .C(_4423_),
    .D(\genblk1[5].u_ce.Xcalc [3]),
    .Y(_4469_)
);

OAI21X1 _11197_ (
    .A(_4421_),
    .B(_4468_),
    .C(_4469_),
    .Y(\genblk1[5].u_ce.X_ [1])
);

INVX1 _11198_ (
    .A(\genblk1[5].u_ce.Ain0 [0]),
    .Y(_4470_)
);

NAND2X1 _11199_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\a[5] [0]),
    .Y(_4471_)
);

OAI21X1 _11200_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_4470_),
    .C(_4471_),
    .Y(_4330_)
);

INVX1 _11201_ (
    .A(\genblk1[5].u_ce.Ain0 [1]),
    .Y(_4472_)
);

NAND2X1 _11202_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\a[5] [1]),
    .Y(_4473_)
);

OAI21X1 _11203_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_4472_),
    .C(_4473_),
    .Y(_4331_)
);

INVX8 _11204_ (
    .A(\genblk1[5].u_ce.Vld_bF$buf3 ),
    .Y(_4474_)
);

NAND2X1 _11205_ (
    .A(\genblk1[5].u_ce.Ycalc [2]),
    .B(_4474__bF$buf4),
    .Y(_4475_)
);

INVX2 _11206_ (
    .A(1'h1),
    .Y(_4476_)
);

NOR2X1 _11207_ (
    .A(1'h1),
    .B(1'h0),
    .Y(_4477_)
);

NAND2X1 _11208_ (
    .A(_4476_),
    .B(_4477_),
    .Y(_4478_)
);

INVX2 _11209_ (
    .A(_4478_),
    .Y(_4479_)
);

INVX8 _11210_ (
    .A(1'h0),
    .Y(_4480_)
);

MUX2X1 _11211_ (
    .A(\genblk1[5].u_ce.Xin12b [4]),
    .B(\genblk1[5].u_ce.Xin1 [1]),
    .S(1'h1),
    .Y(_4481_)
);

MUX2X1 _11212_ (
    .A(\genblk1[5].u_ce.Xin1 [0]),
    .B(\genblk1[5].u_ce.Xin0 [1]),
    .S(1'h1),
    .Y(_4482_)
);

MUX2X1 _11213_ (
    .A(_4482_),
    .B(_4481_),
    .S(_4480__bF$buf4),
    .Y(_4483_)
);

MUX2X1 _11214_ (
    .A(\genblk1[5].u_ce.Xin12b [8]),
    .B(\genblk1[5].u_ce.Xin12b [7]),
    .S(1'h1),
    .Y(_4484_)
);

MUX2X1 _11215_ (
    .A(\genblk1[5].u_ce.Xin12b [6]),
    .B(\genblk1[5].u_ce.Xin12b [5]),
    .S(1'h1),
    .Y(_4485_)
);

MUX2X1 _11216_ (
    .A(_4485_),
    .B(_4484_),
    .S(_4480__bF$buf3),
    .Y(_4486_)
);

MUX2X1 _11217_ (
    .A(_4486_),
    .B(_4483_),
    .S(1'h1),
    .Y(_4487_)
);

INVX1 _11218_ (
    .A(_4487_),
    .Y(_4488_)
);

MUX2X1 _11219_ (
    .A(\genblk1[5].u_ce.Xin1 [1]),
    .B(\genblk1[5].u_ce.Xin1 [0]),
    .S(1'h1),
    .Y(_4489_)
);

MUX2X1 _11220_ (
    .A(\genblk1[5].u_ce.Xin0 [1]),
    .B(\genblk1[5].u_ce.Xin0 [0]),
    .S(1'h1),
    .Y(_4490_)
);

MUX2X1 _11221_ (
    .A(_4490_),
    .B(_4489_),
    .S(_4480__bF$buf2),
    .Y(_4491_)
);

MUX2X1 _11222_ (
    .A(\genblk1[5].u_ce.Xin12b [7]),
    .B(\genblk1[5].u_ce.Xin12b [6]),
    .S(1'h1),
    .Y(_4492_)
);

MUX2X1 _11223_ (
    .A(\genblk1[5].u_ce.Xin12b [5]),
    .B(\genblk1[5].u_ce.Xin12b [4]),
    .S(1'h1),
    .Y(_4493_)
);

MUX2X1 _11224_ (
    .A(_4493_),
    .B(_4492_),
    .S(_4480__bF$buf1),
    .Y(_4494_)
);

MUX2X1 _11225_ (
    .A(_4494_),
    .B(_4491_),
    .S(1'h1),
    .Y(_4495_)
);

OAI21X1 _11226_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf4 ),
    .B(_4495_),
    .C(_4488_),
    .Y(_4496_)
);

NOR2X1 _11227_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4495_),
    .Y(_4497_)
);

NAND2X1 _11228_ (
    .A(_4487_),
    .B(_4497_),
    .Y(_4498_)
);

NAND3X1 _11229_ (
    .A(\genblk1[5].u_ce.Yin0 [1]),
    .B(_4496_),
    .C(_4498_),
    .Y(_4499_)
);

NOR2X1 _11230_ (
    .A(\genblk1[5].u_ce.Yin0 [0]),
    .B(_4495_),
    .Y(_4500_)
);

AOI21X1 _11231_ (
    .A(_4498_),
    .B(_4496_),
    .C(\genblk1[5].u_ce.Yin0 [1]),
    .Y(_4501_)
);

OAI21X1 _11232_ (
    .A(_4500_),
    .B(_4501_),
    .C(_4499_),
    .Y(_4502_)
);

INVX1 _11233_ (
    .A(\genblk1[5].u_ce.Yin1 [0]),
    .Y(_4503_)
);

MUX2X1 _11234_ (
    .A(\genblk1[5].u_ce.Xin12b [9]),
    .B(\genblk1[5].u_ce.Xin12b [8]),
    .S(1'h1),
    .Y(_4504_)
);

MUX2X1 _11235_ (
    .A(_4504_),
    .B(_4492_),
    .S(1'h0),
    .Y(_4505_)
);

AND2X2 _11236_ (
    .A(_4505_),
    .B(1'h1),
    .Y(_4506_)
);

INVX4 _11237_ (
    .A(1'h1),
    .Y(_4507_)
);

NAND2X1 _11238_ (
    .A(_4507__bF$buf3),
    .B(_4480__bF$buf0),
    .Y(_4508_)
);

NAND2X1 _11239_ (
    .A(1'h0),
    .B(_4507__bF$buf2),
    .Y(_4509_)
);

OAI22X1 _11240_ (
    .A(_4508_),
    .B(_4489_),
    .C(_4493_),
    .D(_4509_),
    .Y(_4510_)
);

INVX1 _11241_ (
    .A(\genblk1[5].u_ce.Xin1 [1]),
    .Y(_4511_)
);

NAND2X1 _11242_ (
    .A(_4476_),
    .B(_4511_),
    .Y(_4512_)
);

INVX1 _11243_ (
    .A(\genblk1[5].u_ce.Xin12b [4]),
    .Y(_4513_)
);

NAND2X1 _11244_ (
    .A(1'h1),
    .B(_4513_),
    .Y(_4514_)
);

NAND3X1 _11245_ (
    .A(1'h0),
    .B(_4514_),
    .C(_4512_),
    .Y(_4515_)
);

INVX1 _11246_ (
    .A(\genblk1[5].u_ce.Xin0 [1]),
    .Y(_4516_)
);

NAND2X1 _11247_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Xin1 [0]),
    .Y(_4517_)
);

OAI21X1 _11248_ (
    .A(1'h1),
    .B(_4516_),
    .C(_4517_),
    .Y(_4518_)
);

NAND2X1 _11249_ (
    .A(_4480__bF$buf4),
    .B(_4518_),
    .Y(_4519_)
);

NAND3X1 _11250_ (
    .A(_4507__bF$buf1),
    .B(_4515_),
    .C(_4519_),
    .Y(_4520_)
);

INVX1 _11251_ (
    .A(\genblk1[5].u_ce.Xin12b [5]),
    .Y(_4521_)
);

NAND2X1 _11252_ (
    .A(_4476_),
    .B(_4521_),
    .Y(_4522_)
);

INVX1 _11253_ (
    .A(\genblk1[5].u_ce.Xin12b [6]),
    .Y(_4523_)
);

NAND2X1 _11254_ (
    .A(1'h1),
    .B(_4523_),
    .Y(_4524_)
);

NAND3X1 _11255_ (
    .A(_4480__bF$buf3),
    .B(_4524_),
    .C(_4522_),
    .Y(_4525_)
);

INVX1 _11256_ (
    .A(\genblk1[5].u_ce.Xin12b [7]),
    .Y(_4526_)
);

NAND2X1 _11257_ (
    .A(_4476_),
    .B(_4526_),
    .Y(_4527_)
);

INVX1 _11258_ (
    .A(\genblk1[5].u_ce.Xin12b [8]),
    .Y(_4528_)
);

NAND2X1 _11259_ (
    .A(1'h1),
    .B(_4528_),
    .Y(_4529_)
);

NAND3X1 _11260_ (
    .A(1'h0),
    .B(_4529_),
    .C(_4527_),
    .Y(_4530_)
);

NAND3X1 _11261_ (
    .A(1'h1),
    .B(_4525_),
    .C(_4530_),
    .Y(_4531_)
);

INVX1 _11262_ (
    .A(\genblk1[5].u_ce.Xin1 [0]),
    .Y(_4532_)
);

NAND2X1 _11263_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Xin1 [1]),
    .Y(_4533_)
);

OAI21X1 _11264_ (
    .A(1'h1),
    .B(_4532_),
    .C(_4533_),
    .Y(_4534_)
);

NAND2X1 _11265_ (
    .A(1'h0),
    .B(_4534_),
    .Y(_4535_)
);

INVX1 _11266_ (
    .A(\genblk1[5].u_ce.Xin0 [0]),
    .Y(_4536_)
);

NAND2X1 _11267_ (
    .A(\genblk1[5].u_ce.Xin0 [1]),
    .B(1'h1),
    .Y(_4537_)
);

OAI21X1 _11268_ (
    .A(1'h1),
    .B(_4536_),
    .C(_4537_),
    .Y(_4538_)
);

NAND2X1 _11269_ (
    .A(_4480__bF$buf2),
    .B(_4538_),
    .Y(_4539_)
);

NAND3X1 _11270_ (
    .A(_4507__bF$buf0),
    .B(_4535_),
    .C(_4539_),
    .Y(_4540_)
);

NAND2X1 _11271_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Xin12b [5]),
    .Y(_4541_)
);

OAI21X1 _11272_ (
    .A(1'h1),
    .B(_4513_),
    .C(_4541_),
    .Y(_4542_)
);

NAND2X1 _11273_ (
    .A(_4480__bF$buf1),
    .B(_4542_),
    .Y(_4543_)
);

NAND2X1 _11274_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Xin12b [7]),
    .Y(_4544_)
);

OAI21X1 _11275_ (
    .A(1'h1),
    .B(_4523_),
    .C(_4544_),
    .Y(_4545_)
);

NAND2X1 _11276_ (
    .A(1'h0),
    .B(_4545_),
    .Y(_4546_)
);

NAND3X1 _11277_ (
    .A(1'h1),
    .B(_4543_),
    .C(_4546_),
    .Y(_4547_)
);

AOI22X1 _11278_ (
    .A(_4520_),
    .B(_4531_),
    .C(_4540_),
    .D(_4547_),
    .Y(_4548_)
);

NOR2X1 _11279_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4548_),
    .Y(_4549_)
);

OAI21X1 _11280_ (
    .A(_4506_),
    .B(_4510_),
    .C(_4549_),
    .Y(_4550_)
);

AOI21X1 _11281_ (
    .A(1'h1),
    .B(_4505_),
    .C(_4510_),
    .Y(_4551_)
);

OAI21X1 _11282_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .B(_4548_),
    .C(_4551_),
    .Y(_4552_)
);

NAND3X1 _11283_ (
    .A(_4503_),
    .B(_4552_),
    .C(_4550_),
    .Y(_4553_)
);

NAND2X1 _11284_ (
    .A(_4551_),
    .B(_4549_),
    .Y(_4554_)
);

OAI22X1 _11285_ (
    .A(_4506_),
    .B(_4510_),
    .C(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .D(_4548_),
    .Y(_4555_)
);

NAND3X1 _11286_ (
    .A(\genblk1[5].u_ce.Yin1 [0]),
    .B(_4555_),
    .C(_4554_),
    .Y(_4556_)
);

NAND3X1 _11287_ (
    .A(_4553_),
    .B(_4556_),
    .C(_4502_),
    .Y(_4557_)
);

INVX1 _11288_ (
    .A(\genblk1[5].u_ce.Yin0 [1]),
    .Y(_4558_)
);

NAND2X1 _11289_ (
    .A(_4488_),
    .B(_4497_),
    .Y(_4559_)
);

OAI21X1 _11290_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf4 ),
    .B(_4495_),
    .C(_4487_),
    .Y(_4560_)
);

AOI21X1 _11291_ (
    .A(_4559_),
    .B(_4560_),
    .C(_4558_),
    .Y(_4561_)
);

INVX1 _11292_ (
    .A(_4500_),
    .Y(_4562_)
);

NAND3X1 _11293_ (
    .A(_4558_),
    .B(_4560_),
    .C(_4559_),
    .Y(_4563_)
);

AOI21X1 _11294_ (
    .A(_4562_),
    .B(_4563_),
    .C(_4561_),
    .Y(_4564_)
);

AOI21X1 _11295_ (
    .A(_4554_),
    .B(_4555_),
    .C(\genblk1[5].u_ce.Yin1 [0]),
    .Y(_4565_)
);

AOI21X1 _11296_ (
    .A(_4550_),
    .B(_4552_),
    .C(_4503_),
    .Y(_4566_)
);

OAI21X1 _11297_ (
    .A(_4565_),
    .B(_4566_),
    .C(_4564_),
    .Y(_4567_)
);

AOI21X1 _11298_ (
    .A(_4557_),
    .B(_4567_),
    .C(_4479_),
    .Y(_4568_)
);

INVX8 _11299_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_4569_)
);

NAND3X1 _11300_ (
    .A(_4507__bF$buf3),
    .B(_4476_),
    .C(_4569__bF$buf5),
    .Y(_4570_)
);

OAI21X1 _11301_ (
    .A(1'h0),
    .B(_4570_),
    .C(\genblk1[5].u_ce.Vld_bF$buf2 ),
    .Y(_4571_)
);

OAI21X1 _11302_ (
    .A(_4571_),
    .B(_4568_),
    .C(_4475_),
    .Y(_4332_)
);

INVX1 _11303_ (
    .A(\genblk1[5].u_ce.Ycalc [3]),
    .Y(_4572_)
);

INVX1 _11304_ (
    .A(\genblk1[5].u_ce.Xin12b [9]),
    .Y(_4573_)
);

NAND2X1 _11305_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Xin12b [10]),
    .Y(_4574_)
);

OAI21X1 _11306_ (
    .A(1'h1),
    .B(_4573_),
    .C(_4574_),
    .Y(_4575_)
);

NAND2X1 _11307_ (
    .A(1'h0),
    .B(_4575_),
    .Y(_4576_)
);

OAI21X1 _11308_ (
    .A(1'h0),
    .B(_4484_),
    .C(_4576_),
    .Y(_4577_)
);

OAI22X1 _11309_ (
    .A(_4508_),
    .B(_4481_),
    .C(_4485_),
    .D(_4509_),
    .Y(_4578_)
);

AOI21X1 _11310_ (
    .A(_4577_),
    .B(1'h1),
    .C(_4578_),
    .Y(_4579_)
);

NAND3X1 _11311_ (
    .A(_4551_),
    .B(_4487_),
    .C(_4495_),
    .Y(_4580_)
);

INVX1 _11312_ (
    .A(_4580_),
    .Y(_4581_)
);

NOR2X1 _11313_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4581_),
    .Y(_4582_)
);

NAND2X1 _11314_ (
    .A(_4579_),
    .B(_4582_),
    .Y(_4583_)
);

INVX1 _11315_ (
    .A(_4579_),
    .Y(_4584_)
);

OAI21X1 _11316_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .B(_4581_),
    .C(_4584_),
    .Y(_4585_)
);

AOI21X1 _11317_ (
    .A(_4583_),
    .B(_4585_),
    .C(\genblk1[5].u_ce.Yin1 [1]),
    .Y(_4586_)
);

AOI21X1 _11318_ (
    .A(_4502_),
    .B(_4553_),
    .C(_4566_),
    .Y(_4587_)
);

NAND3X1 _11319_ (
    .A(\genblk1[5].u_ce.Yin1 [1]),
    .B(_4585_),
    .C(_4583_),
    .Y(_4588_)
);

NAND2X1 _11320_ (
    .A(_4588_),
    .B(_4587_),
    .Y(_4589_)
);

OAI21X1 _11321_ (
    .A(_4565_),
    .B(_4564_),
    .C(_4556_),
    .Y(_4590_)
);

INVX1 _11322_ (
    .A(\genblk1[5].u_ce.Yin1 [1]),
    .Y(_4591_)
);

NAND2X1 _11323_ (
    .A(_4584_),
    .B(_4582_),
    .Y(_4592_)
);

OAI21X1 _11324_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .B(_4581_),
    .C(_4579_),
    .Y(_4593_)
);

AOI21X1 _11325_ (
    .A(_4592_),
    .B(_4593_),
    .C(_4591_),
    .Y(_4594_)
);

OAI21X1 _11326_ (
    .A(_4586_),
    .B(_4594_),
    .C(_4590_),
    .Y(_4595_)
);

OAI21X1 _11327_ (
    .A(_4586_),
    .B(_4589_),
    .C(_4595_),
    .Y(_4596_)
);

OAI21X1 _11328_ (
    .A(_4569__bF$buf4),
    .B(_4478_),
    .C(\genblk1[5].u_ce.Vld_bF$buf1 ),
    .Y(_4597_)
);

INVX1 _11329_ (
    .A(_4597_),
    .Y(_4598_)
);

OAI21X1 _11330_ (
    .A(_4479_),
    .B(_4596_),
    .C(_4598_),
    .Y(_4599_)
);

OAI21X1 _11331_ (
    .A(_4572_),
    .B(\genblk1[5].u_ce.Vld_bF$buf0 ),
    .C(_4599_),
    .Y(_4333_)
);

INVX1 _11332_ (
    .A(_4571_),
    .Y(_4600_)
);

INVX1 _11333_ (
    .A(\genblk1[5].u_ce.Yin12b [4]),
    .Y(_4601_)
);

NAND3X1 _11334_ (
    .A(_4551_),
    .B(_4579_),
    .C(_4548_),
    .Y(_4602_)
);

INVX1 _11335_ (
    .A(\genblk1[5].u_ce.Xin12b [10]),
    .Y(_4603_)
);

NAND2X1 _11336_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Xin12b [11]),
    .Y(_4604_)
);

OAI21X1 _11337_ (
    .A(1'h1),
    .B(_4603_),
    .C(_4604_),
    .Y(_4605_)
);

NAND2X1 _11338_ (
    .A(_4480__bF$buf0),
    .B(_4504_),
    .Y(_4606_)
);

OAI21X1 _11339_ (
    .A(_4480__bF$buf4),
    .B(_4605_),
    .C(_4606_),
    .Y(_4607_)
);

NAND2X1 _11340_ (
    .A(_4507__bF$buf2),
    .B(_4494_),
    .Y(_4608_)
);

OAI21X1 _11341_ (
    .A(_4507__bF$buf1),
    .B(_4607_),
    .C(_4608_),
    .Y(_4609_)
);

INVX1 _11342_ (
    .A(_4609_),
    .Y(_4610_)
);

NAND3X1 _11343_ (
    .A(_4569__bF$buf3),
    .B(_4610_),
    .C(_4602_),
    .Y(_4611_)
);

INVX1 _11344_ (
    .A(_4611_),
    .Y(_4612_)
);

AOI21X1 _11345_ (
    .A(_4602_),
    .B(_4569__bF$buf2),
    .C(_4610_),
    .Y(_4613_)
);

OAI21X1 _11346_ (
    .A(_4613_),
    .B(_4612_),
    .C(_4601_),
    .Y(_4614_)
);

OAI21X1 _11347_ (
    .A(_4580_),
    .B(_4584_),
    .C(_4569__bF$buf1),
    .Y(_4615_)
);

NAND2X1 _11348_ (
    .A(_4609_),
    .B(_4615_),
    .Y(_4616_)
);

NAND3X1 _11349_ (
    .A(\genblk1[5].u_ce.Yin12b [4]),
    .B(_4611_),
    .C(_4616_),
    .Y(_4617_)
);

NAND2X1 _11350_ (
    .A(_4617_),
    .B(_4614_),
    .Y(_4618_)
);

INVX1 _11351_ (
    .A(_4586_),
    .Y(_4619_)
);

OAI21X1 _11352_ (
    .A(_4594_),
    .B(_4590_),
    .C(_4619_),
    .Y(_4620_)
);

AOI21X1 _11353_ (
    .A(_4620_),
    .B(_4618_),
    .C(_4479_),
    .Y(_4621_)
);

OAI21X1 _11354_ (
    .A(_4618_),
    .B(_4620_),
    .C(_4621_),
    .Y(_4622_)
);

AOI22X1 _11355_ (
    .A(_4437_),
    .B(_4474__bF$buf3),
    .C(_4622_),
    .D(_4600_),
    .Y(_4334_)
);

INVX1 _11356_ (
    .A(_4617_),
    .Y(_4623_)
);

AOI21X1 _11357_ (
    .A(_4587_),
    .B(_4588_),
    .C(_4586_),
    .Y(_4624_)
);

AOI21X1 _11358_ (
    .A(_4624_),
    .B(_4614_),
    .C(_4623_),
    .Y(_4625_)
);

INVX1 _11359_ (
    .A(\genblk1[5].u_ce.Yin12b [5]),
    .Y(_4626_)
);

NAND3X1 _11360_ (
    .A(_4579_),
    .B(_4610_),
    .C(_4581_),
    .Y(_4627_)
);

INVX1 _11361_ (
    .A(\genblk1[5].u_ce.Xin12b [11]),
    .Y(_4628_)
);

NOR2X1 _11362_ (
    .A(_4480__bF$buf3),
    .B(_4628_),
    .Y(_4629_)
);

AOI21X1 _11363_ (
    .A(_4480__bF$buf2),
    .B(_4575_),
    .C(_4629_),
    .Y(_4630_)
);

NAND2X1 _11364_ (
    .A(_4507__bF$buf0),
    .B(_4486_),
    .Y(_4631_)
);

OAI21X1 _11365_ (
    .A(_4507__bF$buf3),
    .B(_4630_),
    .C(_4631_),
    .Y(_4632_)
);

NAND3X1 _11366_ (
    .A(_4569__bF$buf0),
    .B(_4632_),
    .C(_4627_),
    .Y(_4633_)
);

INVX1 _11367_ (
    .A(_4632_),
    .Y(_4634_)
);

OAI21X1 _11368_ (
    .A(_4609_),
    .B(_4602_),
    .C(_4569__bF$buf5),
    .Y(_4635_)
);

NAND2X1 _11369_ (
    .A(_4634_),
    .B(_4635_),
    .Y(_4636_)
);

NAND3X1 _11370_ (
    .A(_4626_),
    .B(_4636_),
    .C(_4633_),
    .Y(_4637_)
);

NAND3X1 _11371_ (
    .A(_4569__bF$buf4),
    .B(_4634_),
    .C(_4627_),
    .Y(_4638_)
);

NAND2X1 _11372_ (
    .A(_4632_),
    .B(_4635_),
    .Y(_4639_)
);

NAND3X1 _11373_ (
    .A(\genblk1[5].u_ce.Yin12b [5]),
    .B(_4639_),
    .C(_4638_),
    .Y(_4640_)
);

NAND2X1 _11374_ (
    .A(_4637_),
    .B(_4640_),
    .Y(_4641_)
);

INVX1 _11375_ (
    .A(_4641_),
    .Y(_4642_)
);

NOR2X1 _11376_ (
    .A(_4642_),
    .B(_4625_),
    .Y(_4643_)
);

OAI21X1 _11377_ (
    .A(_4618_),
    .B(_4620_),
    .C(_4617_),
    .Y(_4644_)
);

OAI21X1 _11378_ (
    .A(_4641_),
    .B(_4644_),
    .C(_4478_),
    .Y(_4645_)
);

OAI21X1 _11379_ (
    .A(_4645_),
    .B(_4643_),
    .C(_4600_),
    .Y(_4646_)
);

OAI21X1 _11380_ (
    .A(_4445_),
    .B(\genblk1[5].u_ce.Vld_bF$buf3 ),
    .C(_4646_),
    .Y(_4335_)
);

NOR2X1 _11381_ (
    .A(_4618_),
    .B(_4641_),
    .Y(_4647_)
);

OAI21X1 _11382_ (
    .A(_4617_),
    .B(_4641_),
    .C(_4640_),
    .Y(_4648_)
);

AOI21X1 _11383_ (
    .A(_4647_),
    .B(_4624_),
    .C(_4648_),
    .Y(_4649_)
);

INVX1 _11384_ (
    .A(\genblk1[5].u_ce.Yin12b [6]),
    .Y(_4650_)
);

NOR2X1 _11385_ (
    .A(_4609_),
    .B(_4602_),
    .Y(_4651_)
);

NAND2X1 _11386_ (
    .A(_4634_),
    .B(_4651_),
    .Y(_4652_)
);

AOI21X1 _11387_ (
    .A(_4480__bF$buf1),
    .B(_4605_),
    .C(_4629_),
    .Y(_4653_)
);

NAND2X1 _11388_ (
    .A(_4507__bF$buf2),
    .B(_4505_),
    .Y(_4654_)
);

OAI21X1 _11389_ (
    .A(_4507__bF$buf1),
    .B(_4653_),
    .C(_4654_),
    .Y(_4655_)
);

NAND3X1 _11390_ (
    .A(_4569__bF$buf3),
    .B(_4655_),
    .C(_4652_),
    .Y(_4656_)
);

NOR3X1 _11391_ (
    .A(_4609_),
    .B(_4632_),
    .C(_4602_),
    .Y(_4657_)
);

INVX1 _11392_ (
    .A(_4655_),
    .Y(_4658_)
);

OAI21X1 _11393_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf4 ),
    .B(_4657_),
    .C(_4658_),
    .Y(_4659_)
);

NAND3X1 _11394_ (
    .A(_4650_),
    .B(_4659_),
    .C(_4656_),
    .Y(_4660_)
);

NAND3X1 _11395_ (
    .A(_4569__bF$buf2),
    .B(_4658_),
    .C(_4652_),
    .Y(_4661_)
);

OAI21X1 _11396_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4657_),
    .C(_4655_),
    .Y(_4662_)
);

NAND3X1 _11397_ (
    .A(\genblk1[5].u_ce.Yin12b [6]),
    .B(_4662_),
    .C(_4661_),
    .Y(_4663_)
);

AND2X2 _11398_ (
    .A(_4660_),
    .B(_4663_),
    .Y(_4664_)
);

INVX1 _11399_ (
    .A(_4664_),
    .Y(_4665_)
);

AOI21X1 _11400_ (
    .A(_4649_),
    .B(_4665_),
    .C(_4479_),
    .Y(_4666_)
);

OAI21X1 _11401_ (
    .A(_4649_),
    .B(_4665_),
    .C(_4666_),
    .Y(_4667_)
);

AOI22X1 _11402_ (
    .A(_4436_),
    .B(_4474__bF$buf2),
    .C(_4667_),
    .D(_4600_),
    .Y(_4336_)
);

AND2X2 _11403_ (
    .A(_4614_),
    .B(_4617_),
    .Y(_4668_)
);

NAND3X1 _11404_ (
    .A(_4637_),
    .B(_4640_),
    .C(_4668_),
    .Y(_4669_)
);

INVX1 _11405_ (
    .A(_4640_),
    .Y(_4670_)
);

AOI21X1 _11406_ (
    .A(_4623_),
    .B(_4637_),
    .C(_4670_),
    .Y(_4671_)
);

OAI21X1 _11407_ (
    .A(_4620_),
    .B(_4669_),
    .C(_4671_),
    .Y(_4672_)
);

INVX1 _11408_ (
    .A(_4663_),
    .Y(_4673_)
);

AOI21X1 _11409_ (
    .A(_4672_),
    .B(_4660_),
    .C(_4673_),
    .Y(_4674_)
);

INVX1 _11410_ (
    .A(\genblk1[5].u_ce.Yin12b [7]),
    .Y(_4675_)
);

NAND2X1 _11411_ (
    .A(_4658_),
    .B(_4657_),
    .Y(_4676_)
);

NOR2X1 _11412_ (
    .A(_4507__bF$buf0),
    .B(_4628_),
    .Y(_4677_)
);

AOI21X1 _11413_ (
    .A(_4577_),
    .B(_4507__bF$buf3),
    .C(_4677_),
    .Y(_4678_)
);

INVX1 _11414_ (
    .A(_4678_),
    .Y(_4679_)
);

NAND3X1 _11415_ (
    .A(_4569__bF$buf1),
    .B(_4679_),
    .C(_4676_),
    .Y(_4680_)
);

AND2X2 _11416_ (
    .A(_4657_),
    .B(_4658_),
    .Y(_4681_)
);

OAI21X1 _11417_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4681_),
    .C(_4678_),
    .Y(_4682_)
);

NAND3X1 _11418_ (
    .A(_4675_),
    .B(_4680_),
    .C(_4682_),
    .Y(_4683_)
);

NAND3X1 _11419_ (
    .A(_4569__bF$buf0),
    .B(_4678_),
    .C(_4676_),
    .Y(_4684_)
);

OAI21X1 _11420_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .B(_4681_),
    .C(_4679_),
    .Y(_4685_)
);

NAND3X1 _11421_ (
    .A(\genblk1[5].u_ce.Yin12b [7]),
    .B(_4684_),
    .C(_4685_),
    .Y(_4686_)
);

AND2X2 _11422_ (
    .A(_4683_),
    .B(_4686_),
    .Y(_4687_)
);

NOR2X1 _11423_ (
    .A(_4687_),
    .B(_4674_),
    .Y(_4688_)
);

NAND2X1 _11424_ (
    .A(_4476_),
    .B(_4480__bF$buf0),
    .Y(_4689_)
);

NAND2X1 _11425_ (
    .A(_4687_),
    .B(_4674_),
    .Y(_4690_)
);

OAI21X1 _11426_ (
    .A(1'h1),
    .B(_4689_),
    .C(_4690_),
    .Y(_4691_)
);

OAI21X1 _11427_ (
    .A(_4688_),
    .B(_4691_),
    .C(_4598_),
    .Y(_4692_)
);

OAI21X1 _11428_ (
    .A(_4444_),
    .B(\genblk1[5].u_ce.Vld_bF$buf2 ),
    .C(_4692_),
    .Y(_4337_)
);

INVX1 _11429_ (
    .A(\genblk1[5].u_ce.Ycalc [8]),
    .Y(_4693_)
);

AOI21X1 _11430_ (
    .A(_4682_),
    .B(_4680_),
    .C(_4675_),
    .Y(_4694_)
);

OAI21X1 _11431_ (
    .A(_4673_),
    .B(_4694_),
    .C(_4683_),
    .Y(_4695_)
);

NAND3X1 _11432_ (
    .A(_4664_),
    .B(_4687_),
    .C(_4672_),
    .Y(_4696_)
);

INVX1 _11433_ (
    .A(\genblk1[5].u_ce.Yin12b [8]),
    .Y(_4697_)
);

NAND3X1 _11434_ (
    .A(_4658_),
    .B(_4678_),
    .C(_4657_),
    .Y(_4698_)
);

INVX1 _11435_ (
    .A(_4677_),
    .Y(_4699_)
);

OAI21X1 _11436_ (
    .A(1'h1),
    .B(_4607_),
    .C(_4699_),
    .Y(_4700_)
);

NAND3X1 _11437_ (
    .A(_4569__bF$buf5),
    .B(_4700_),
    .C(_4698_),
    .Y(_4701_)
);

INVX1 _11438_ (
    .A(_4700_),
    .Y(_4702_)
);

NAND2X1 _11439_ (
    .A(_4569__bF$buf4),
    .B(_4698_),
    .Y(_4703_)
);

NAND2X1 _11440_ (
    .A(_4702_),
    .B(_4703_),
    .Y(_4704_)
);

NAND3X1 _11441_ (
    .A(_4697_),
    .B(_4701_),
    .C(_4704_),
    .Y(_4705_)
);

NAND3X1 _11442_ (
    .A(_4569__bF$buf3),
    .B(_4702_),
    .C(_4698_),
    .Y(_4706_)
);

NAND2X1 _11443_ (
    .A(_4700_),
    .B(_4703_),
    .Y(_4707_)
);

NAND3X1 _11444_ (
    .A(\genblk1[5].u_ce.Yin12b [8]),
    .B(_4706_),
    .C(_4707_),
    .Y(_4708_)
);

AND2X2 _11445_ (
    .A(_4705_),
    .B(_4708_),
    .Y(_4709_)
);

INVX1 _11446_ (
    .A(_4709_),
    .Y(_4710_)
);

AOI21X1 _11447_ (
    .A(_4696_),
    .B(_4695_),
    .C(_4710_),
    .Y(_4711_)
);

NAND3X1 _11448_ (
    .A(_4683_),
    .B(_4686_),
    .C(_4664_),
    .Y(_4712_)
);

OAI21X1 _11449_ (
    .A(_4712_),
    .B(_4649_),
    .C(_4695_),
    .Y(_4713_)
);

OAI21X1 _11450_ (
    .A(_4709_),
    .B(_4713_),
    .C(_4478_),
    .Y(_4714_)
);

OR2X2 _11451_ (
    .A(_4714_),
    .B(_4711_),
    .Y(_4715_)
);

AOI22X1 _11452_ (
    .A(_4693_),
    .B(_4474__bF$buf1),
    .C(_4715_),
    .D(_4598_),
    .Y(_4338_)
);

INVX1 _11453_ (
    .A(\genblk1[5].u_ce.Ycalc [9]),
    .Y(_4716_)
);

INVX1 _11454_ (
    .A(_4708_),
    .Y(_4717_)
);

NOR2X1 _11455_ (
    .A(_4717_),
    .B(_4711_),
    .Y(_4718_)
);

INVX1 _11456_ (
    .A(\genblk1[5].u_ce.Yin12b [9]),
    .Y(_4719_)
);

OAI21X1 _11457_ (
    .A(1'h1),
    .B(_4630_),
    .C(_4699_),
    .Y(_4720_)
);

INVX1 _11458_ (
    .A(_4720_),
    .Y(_4721_)
);

OAI21X1 _11459_ (
    .A(_4700_),
    .B(_4698_),
    .C(_4569__bF$buf2),
    .Y(_4722_)
);

NAND2X1 _11460_ (
    .A(_4721_),
    .B(_4722_),
    .Y(_4723_)
);

NAND3X1 _11461_ (
    .A(_4678_),
    .B(_4702_),
    .C(_4681_),
    .Y(_4724_)
);

NAND3X1 _11462_ (
    .A(_4569__bF$buf1),
    .B(_4720_),
    .C(_4724_),
    .Y(_4725_)
);

NAND3X1 _11463_ (
    .A(_4719_),
    .B(_4723_),
    .C(_4725_),
    .Y(_4726_)
);

AND2X2 _11464_ (
    .A(_4722_),
    .B(_4721_),
    .Y(_4727_)
);

NOR2X1 _11465_ (
    .A(_4721_),
    .B(_4722_),
    .Y(_4728_)
);

OAI21X1 _11466_ (
    .A(_4728_),
    .B(_4727_),
    .C(\genblk1[5].u_ce.Yin12b [9]),
    .Y(_4729_)
);

NAND2X1 _11467_ (
    .A(_4726_),
    .B(_4729_),
    .Y(_4730_)
);

AOI21X1 _11468_ (
    .A(_4718_),
    .B(_4730_),
    .C(_4479_),
    .Y(_4731_)
);

OAI21X1 _11469_ (
    .A(_4718_),
    .B(_4730_),
    .C(_4731_),
    .Y(_4732_)
);

AOI22X1 _11470_ (
    .A(_4716_),
    .B(_4474__bF$buf0),
    .C(_4732_),
    .D(_4598_),
    .Y(_4339_)
);

OAI21X1 _11471_ (
    .A(_4708_),
    .B(_4730_),
    .C(_4729_),
    .Y(_4733_)
);

NAND3X1 _11472_ (
    .A(_4726_),
    .B(_4729_),
    .C(_4709_),
    .Y(_4734_)
);

AOI21X1 _11473_ (
    .A(_4695_),
    .B(_4696_),
    .C(_4734_),
    .Y(_4735_)
);

INVX1 _11474_ (
    .A(\genblk1[5].u_ce.Yin12b [10]),
    .Y(_4736_)
);

OAI21X1 _11475_ (
    .A(1'h1),
    .B(_4653_),
    .C(_4699_),
    .Y(_4737_)
);

INVX1 _11476_ (
    .A(_4737_),
    .Y(_4738_)
);

OAI21X1 _11477_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .B(_4721_),
    .C(_4722_),
    .Y(_4739_)
);

NAND2X1 _11478_ (
    .A(_4738_),
    .B(_4739_),
    .Y(_4740_)
);

OAI21X1 _11479_ (
    .A(_4720_),
    .B(_4724_),
    .C(_4569__bF$buf0),
    .Y(_4741_)
);

NAND2X1 _11480_ (
    .A(_4737_),
    .B(_4741_),
    .Y(_4742_)
);

NAND2X1 _11481_ (
    .A(_4740_),
    .B(_4742_),
    .Y(_4743_)
);

NAND2X1 _11482_ (
    .A(_4736_),
    .B(_4743_),
    .Y(_4744_)
);

NAND3X1 _11483_ (
    .A(\genblk1[5].u_ce.Yin12b [10]),
    .B(_4740_),
    .C(_4742_),
    .Y(_4745_)
);

AND2X2 _11484_ (
    .A(_4744_),
    .B(_4745_),
    .Y(_4746_)
);

OAI21X1 _11485_ (
    .A(_4733_),
    .B(_4735_),
    .C(_4746_),
    .Y(_4747_)
);

INVX1 _11486_ (
    .A(_4729_),
    .Y(_4748_)
);

AOI21X1 _11487_ (
    .A(_4717_),
    .B(_4726_),
    .C(_4748_),
    .Y(_4749_)
);

AND2X2 _11488_ (
    .A(_4729_),
    .B(_4726_),
    .Y(_4750_)
);

NAND3X1 _11489_ (
    .A(_4709_),
    .B(_4750_),
    .C(_4713_),
    .Y(_4751_)
);

NAND2X1 _11490_ (
    .A(_4745_),
    .B(_4744_),
    .Y(_4752_)
);

NAND3X1 _11491_ (
    .A(_4749_),
    .B(_4752_),
    .C(_4751_),
    .Y(_4753_)
);

NAND3X1 _11492_ (
    .A(_4478_),
    .B(_4753_),
    .C(_4747_),
    .Y(_4754_)
);

AOI22X1 _11493_ (
    .A(_4433_),
    .B(_4474__bF$buf4),
    .C(_4754_),
    .D(_4600_),
    .Y(_4340_)
);

INVX1 _11494_ (
    .A(_4745_),
    .Y(_4755_)
);

AOI21X1 _11495_ (
    .A(_4751_),
    .B(_4749_),
    .C(_4752_),
    .Y(_4756_)
);

OAI21X1 _11496_ (
    .A(_4737_),
    .B(_4739_),
    .C(_4569__bF$buf5),
    .Y(_4757_)
);

INVX1 _11497_ (
    .A(_4757_),
    .Y(_4758_)
);

NAND2X1 _11498_ (
    .A(\genblk1[5].u_ce.Yin12b [11]),
    .B(_4628_),
    .Y(_4759_)
);

INVX1 _11499_ (
    .A(\genblk1[5].u_ce.Yin12b [11]),
    .Y(_4760_)
);

NAND2X1 _11500_ (
    .A(\genblk1[5].u_ce.Xin12b [11]),
    .B(_4760_),
    .Y(_4761_)
);

NAND2X1 _11501_ (
    .A(_4759_),
    .B(_4761_),
    .Y(_4762_)
);

OR2X2 _11502_ (
    .A(_4758_),
    .B(_4762_),
    .Y(_4763_)
);

NAND2X1 _11503_ (
    .A(_4762_),
    .B(_4758_),
    .Y(_4764_)
);

NAND2X1 _11504_ (
    .A(_4764_),
    .B(_4763_),
    .Y(_4765_)
);

OAI21X1 _11505_ (
    .A(_4755_),
    .B(_4756_),
    .C(_4765_),
    .Y(_4766_)
);

INVX1 _11506_ (
    .A(_4765_),
    .Y(_4767_)
);

NAND3X1 _11507_ (
    .A(_4745_),
    .B(_4767_),
    .C(_4747_),
    .Y(_4768_)
);

NAND3X1 _11508_ (
    .A(_4478_),
    .B(_4768_),
    .C(_4766_),
    .Y(_4769_)
);

AOI22X1 _11509_ (
    .A(_4441_),
    .B(_4474__bF$buf3),
    .C(_4769_),
    .D(_4598_),
    .Y(_4341_)
);

INVX1 _11510_ (
    .A(\genblk1[5].u_ce.Ycalc [0]),
    .Y(_4770_)
);

OAI21X1 _11511_ (
    .A(1'h1),
    .B(_4689_),
    .C(\genblk1[5].u_ce.Vld_bF$buf1 ),
    .Y(_4771_)
);

INVX2 _11512_ (
    .A(_4771_),
    .Y(_4772_)
);

INVX1 _11513_ (
    .A(\genblk1[5].u_ce.Yin0 [0]),
    .Y(_4773_)
);

AOI21X1 _11514_ (
    .A(_4540_),
    .B(_4547_),
    .C(_4773_),
    .Y(_4774_)
);

OAI21X1 _11515_ (
    .A(_4774_),
    .B(_4500_),
    .C(_4772_),
    .Y(_4775_)
);

OAI21X1 _11516_ (
    .A(_4770_),
    .B(\genblk1[5].u_ce.Vld_bF$buf0 ),
    .C(_4775_),
    .Y(_4342_)
);

NAND2X1 _11517_ (
    .A(\genblk1[5].u_ce.Ycalc [1]),
    .B(_4474__bF$buf2),
    .Y(_4776_)
);

NAND3X1 _11518_ (
    .A(_4562_),
    .B(_4499_),
    .C(_4563_),
    .Y(_4777_)
);

OAI21X1 _11519_ (
    .A(_4561_),
    .B(_4501_),
    .C(_4500_),
    .Y(_4778_)
);

AOI21X1 _11520_ (
    .A(_4778_),
    .B(_4777_),
    .C(_4479_),
    .Y(_4779_)
);

OAI21X1 _11521_ (
    .A(_4474__bF$buf1),
    .B(_4779_),
    .C(_4776_),
    .Y(_4343_)
);

NAND2X1 _11522_ (
    .A(\genblk1[5].u_ce.Xcalc [0]),
    .B(_4474__bF$buf0),
    .Y(_4780_)
);

MUX2X1 _11523_ (
    .A(\genblk1[5].u_ce.Yin12b [7]),
    .B(\genblk1[5].u_ce.Yin12b [6]),
    .S(1'h1),
    .Y(_4781_)
);

NAND2X1 _11524_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin12b [5]),
    .Y(_4782_)
);

OAI21X1 _11525_ (
    .A(1'h1),
    .B(_4601_),
    .C(_4782_),
    .Y(_4783_)
);

NAND2X1 _11526_ (
    .A(_4480__bF$buf4),
    .B(_4783_),
    .Y(_4784_)
);

OAI21X1 _11527_ (
    .A(_4480__bF$buf3),
    .B(_4781_),
    .C(_4784_),
    .Y(_4785_)
);

NAND2X1 _11528_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin1 [1]),
    .Y(_4786_)
);

OAI21X1 _11529_ (
    .A(1'h1),
    .B(_4503_),
    .C(_4786_),
    .Y(_4787_)
);

NAND2X1 _11530_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin0 [1]),
    .Y(_4788_)
);

OAI21X1 _11531_ (
    .A(1'h1),
    .B(_4773_),
    .C(_4788_),
    .Y(_4789_)
);

MUX2X1 _11532_ (
    .A(_4789_),
    .B(_4787_),
    .S(_4480__bF$buf2),
    .Y(_4790_)
);

NAND2X1 _11533_ (
    .A(_4507__bF$buf2),
    .B(_4790_),
    .Y(_4791_)
);

OAI21X1 _11534_ (
    .A(_4507__bF$buf1),
    .B(_4785_),
    .C(_4791_),
    .Y(_4792_)
);

INVX1 _11535_ (
    .A(_4792_),
    .Y(_4793_)
);

NOR2X1 _11536_ (
    .A(\genblk1[5].u_ce.Xin0 [0]),
    .B(_4793_),
    .Y(_4794_)
);

OAI21X1 _11537_ (
    .A(_4536_),
    .B(_4792_),
    .C(_4772_),
    .Y(_4795_)
);

OAI21X1 _11538_ (
    .A(_4795_),
    .B(_4794_),
    .C(_4780_),
    .Y(_4344_)
);

NAND2X1 _11539_ (
    .A(\genblk1[5].u_ce.Xcalc [1]),
    .B(_4474__bF$buf4),
    .Y(_4796_)
);

NOR2X1 _11540_ (
    .A(_4536_),
    .B(_4792_),
    .Y(_4797_)
);

NAND2X1 _11541_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin12b [4]),
    .Y(_4798_)
);

OAI21X1 _11542_ (
    .A(1'h1),
    .B(_4591_),
    .C(_4798_),
    .Y(_4799_)
);

NAND2X1 _11543_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin1 [0]),
    .Y(_4800_)
);

OAI21X1 _11544_ (
    .A(1'h1),
    .B(_4558_),
    .C(_4800_),
    .Y(_4801_)
);

MUX2X1 _11545_ (
    .A(_4801_),
    .B(_4799_),
    .S(_4480__bF$buf1),
    .Y(_4802_)
);

NAND2X1 _11546_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin12b [8]),
    .Y(_4803_)
);

OAI21X1 _11547_ (
    .A(1'h1),
    .B(_4675_),
    .C(_4803_),
    .Y(_4804_)
);

NAND2X1 _11548_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin12b [6]),
    .Y(_4805_)
);

OAI21X1 _11549_ (
    .A(1'h1),
    .B(_4626_),
    .C(_4805_),
    .Y(_4806_)
);

MUX2X1 _11550_ (
    .A(_4806_),
    .B(_4804_),
    .S(_4480__bF$buf0),
    .Y(_4807_)
);

MUX2X1 _11551_ (
    .A(_4807_),
    .B(_4802_),
    .S(1'h1),
    .Y(_4808_)
);

NOR2X1 _11552_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf4 ),
    .B(_4792_),
    .Y(_4809_)
);

NAND2X1 _11553_ (
    .A(_4808_),
    .B(_4809_),
    .Y(_4810_)
);

NAND2X1 _11554_ (
    .A(_4507__bF$buf0),
    .B(_4802_),
    .Y(_4811_)
);

NAND2X1 _11555_ (
    .A(1'h1),
    .B(_4807_),
    .Y(_4812_)
);

NAND2X1 _11556_ (
    .A(_4811_),
    .B(_4812_),
    .Y(_4813_)
);

OAI21X1 _11557_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4792_),
    .C(_4813_),
    .Y(_4814_)
);

NAND3X1 _11558_ (
    .A(\genblk1[5].u_ce.Xin0 [1]),
    .B(_4814_),
    .C(_4810_),
    .Y(_4815_)
);

OAI21X1 _11559_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4792_),
    .C(_4808_),
    .Y(_4816_)
);

NAND2X1 _11560_ (
    .A(_4813_),
    .B(_4809_),
    .Y(_4817_)
);

NAND3X1 _11561_ (
    .A(_4516_),
    .B(_4816_),
    .C(_4817_),
    .Y(_4818_)
);

NAND3X1 _11562_ (
    .A(_4797_),
    .B(_4815_),
    .C(_4818_),
    .Y(_4819_)
);

INVX1 _11563_ (
    .A(_4797_),
    .Y(_4820_)
);

AOI21X1 _11564_ (
    .A(_4817_),
    .B(_4816_),
    .C(_4516_),
    .Y(_4821_)
);

AOI21X1 _11565_ (
    .A(_4810_),
    .B(_4814_),
    .C(\genblk1[5].u_ce.Xin0 [1]),
    .Y(_4822_)
);

OAI21X1 _11566_ (
    .A(_4821_),
    .B(_4822_),
    .C(_4820_),
    .Y(_4823_)
);

AOI21X1 _11567_ (
    .A(_4823_),
    .B(_4819_),
    .C(_4479_),
    .Y(_4824_)
);

OAI21X1 _11568_ (
    .A(_4474__bF$buf3),
    .B(_4824_),
    .C(_4796_),
    .Y(_4345_)
);

OAI21X1 _11569_ (
    .A(_4820_),
    .B(_4822_),
    .C(_4815_),
    .Y(_4825_)
);

MUX2X1 _11570_ (
    .A(\genblk1[5].u_ce.Yin12b [9]),
    .B(\genblk1[5].u_ce.Yin12b [8]),
    .S(1'h1),
    .Y(_4826_)
);

MUX2X1 _11571_ (
    .A(_4826_),
    .B(_4781_),
    .S(1'h0),
    .Y(_4827_)
);

NOR2X1 _11572_ (
    .A(1'h1),
    .B(_4480__bF$buf4),
    .Y(_4828_)
);

NAND2X1 _11573_ (
    .A(_4783_),
    .B(_4828_),
    .Y(_4829_)
);

NAND2X1 _11574_ (
    .A(_4477_),
    .B(_4787_),
    .Y(_4830_)
);

NAND2X1 _11575_ (
    .A(_4830_),
    .B(_4829_),
    .Y(_4831_)
);

AOI21X1 _11576_ (
    .A(1'h1),
    .B(_4827_),
    .C(_4831_),
    .Y(_4832_)
);

NAND2X1 _11577_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin12b [7]),
    .Y(_4833_)
);

OAI21X1 _11578_ (
    .A(1'h1),
    .B(_4650_),
    .C(_4833_),
    .Y(_4834_)
);

MUX2X1 _11579_ (
    .A(_4783_),
    .B(_4834_),
    .S(_4480__bF$buf3),
    .Y(_4835_)
);

NAND2X1 _11580_ (
    .A(1'h1),
    .B(_4835_),
    .Y(_4836_)
);

AOI21X1 _11581_ (
    .A(_4791_),
    .B(_4836_),
    .C(_4808_),
    .Y(_4837_)
);

NOR2X1 _11582_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .B(_4837_),
    .Y(_4838_)
);

NAND2X1 _11583_ (
    .A(_4832_),
    .B(_4838_),
    .Y(_4839_)
);

INVX1 _11584_ (
    .A(_4832_),
    .Y(_4840_)
);

OAI21X1 _11585_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .B(_4837_),
    .C(_4840_),
    .Y(_4841_)
);

AOI21X1 _11586_ (
    .A(_4839_),
    .B(_4841_),
    .C(_4532_),
    .Y(_4842_)
);

NAND3X1 _11587_ (
    .A(_4532_),
    .B(_4841_),
    .C(_4839_),
    .Y(_4843_)
);

INVX1 _11588_ (
    .A(_4843_),
    .Y(_4844_)
);

NOR2X1 _11589_ (
    .A(_4842_),
    .B(_4844_),
    .Y(_4845_)
);

NOR2X1 _11590_ (
    .A(_4825_),
    .B(_4845_),
    .Y(_4846_)
);

AOI21X1 _11591_ (
    .A(_4797_),
    .B(_4818_),
    .C(_4821_),
    .Y(_4847_)
);

INVX1 _11592_ (
    .A(_4845_),
    .Y(_4848_)
);

OAI21X1 _11593_ (
    .A(_4847_),
    .B(_4848_),
    .C(_4772_),
    .Y(_4849_)
);

OAI22X1 _11594_ (
    .A(_4449_),
    .B(\genblk1[5].u_ce.Vld_bF$buf3 ),
    .C(_4846_),
    .D(_4849_),
    .Y(_4346_)
);

NAND2X1 _11595_ (
    .A(\genblk1[5].u_ce.Xcalc [3]),
    .B(_4474__bF$buf2),
    .Y(_4850_)
);

AOI21X1 _11596_ (
    .A(_4825_),
    .B(_4843_),
    .C(_4842_),
    .Y(_4851_)
);

NAND2X1 _11597_ (
    .A(1'h1),
    .B(_4736_),
    .Y(_4852_)
);

OAI21X1 _11598_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin12b [9]),
    .C(_4852_),
    .Y(_4853_)
);

NAND2X1 _11599_ (
    .A(_4480__bF$buf2),
    .B(_4804_),
    .Y(_4854_)
);

OAI21X1 _11600_ (
    .A(_4480__bF$buf1),
    .B(_4853_),
    .C(_4854_),
    .Y(_4855_)
);

NAND2X1 _11601_ (
    .A(_4806_),
    .B(_4828_),
    .Y(_4856_)
);

NAND2X1 _11602_ (
    .A(_4477_),
    .B(_4799_),
    .Y(_4857_)
);

NAND2X1 _11603_ (
    .A(_4857_),
    .B(_4856_),
    .Y(_4858_)
);

AOI21X1 _11604_ (
    .A(_4855_),
    .B(1'h1),
    .C(_4858_),
    .Y(_4859_)
);

NAND3X1 _11605_ (
    .A(_4832_),
    .B(_4813_),
    .C(_4792_),
    .Y(_4860_)
);

NAND2X1 _11606_ (
    .A(_4569__bF$buf4),
    .B(_4860_),
    .Y(_4861_)
);

OR2X2 _11607_ (
    .A(_4861_),
    .B(_4859_),
    .Y(_4862_)
);

INVX1 _11608_ (
    .A(_4860_),
    .Y(_4863_)
);

OAI21X1 _11609_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf4 ),
    .B(_4863_),
    .C(_4859_),
    .Y(_4864_)
);

NAND3X1 _11610_ (
    .A(\genblk1[5].u_ce.Xin1 [1]),
    .B(_4864_),
    .C(_4862_),
    .Y(_4865_)
);

INVX1 _11611_ (
    .A(_4859_),
    .Y(_4866_)
);

OR2X2 _11612_ (
    .A(_4861_),
    .B(_4866_),
    .Y(_4867_)
);

OAI21X1 _11613_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .B(_4863_),
    .C(_4866_),
    .Y(_4868_)
);

NAND3X1 _11614_ (
    .A(_4511_),
    .B(_4868_),
    .C(_4867_),
    .Y(_4869_)
);

NAND2X1 _11615_ (
    .A(_4865_),
    .B(_4869_),
    .Y(_4870_)
);

OR2X2 _11616_ (
    .A(_4851_),
    .B(_4870_),
    .Y(_4871_)
);

NAND2X1 _11617_ (
    .A(_4870_),
    .B(_4851_),
    .Y(_4872_)
);

AOI21X1 _11618_ (
    .A(_4871_),
    .B(_4872_),
    .C(_4479_),
    .Y(_4873_)
);

OAI21X1 _11619_ (
    .A(_4474__bF$buf1),
    .B(_4873_),
    .C(_4850_),
    .Y(_4347_)
);

OAI21X1 _11620_ (
    .A(_4870_),
    .B(_4851_),
    .C(_4865_),
    .Y(_4874_)
);

NAND2X1 _11621_ (
    .A(1'h1),
    .B(\genblk1[5].u_ce.Yin12b [11]),
    .Y(_4875_)
);

OAI21X1 _11622_ (
    .A(1'h1),
    .B(_4736_),
    .C(_4875_),
    .Y(_4876_)
);

NAND2X1 _11623_ (
    .A(1'h0),
    .B(_4876_),
    .Y(_4877_)
);

OAI21X1 _11624_ (
    .A(1'h0),
    .B(_4826_),
    .C(_4877_),
    .Y(_4878_)
);

NAND2X1 _11625_ (
    .A(1'h1),
    .B(_4878_),
    .Y(_4879_)
);

OAI21X1 _11626_ (
    .A(1'h1),
    .B(_4835_),
    .C(_4879_),
    .Y(_4880_)
);

INVX1 _11627_ (
    .A(_4880_),
    .Y(_4881_)
);

OAI21X1 _11628_ (
    .A(_4866_),
    .B(_4860_),
    .C(_4569__bF$buf3),
    .Y(_4882_)
);

OR2X2 _11629_ (
    .A(_4882_),
    .B(_4881_),
    .Y(_4883_)
);

NAND2X1 _11630_ (
    .A(_4881_),
    .B(_4882_),
    .Y(_4884_)
);

NAND3X1 _11631_ (
    .A(\genblk1[5].u_ce.Xin12b [4]),
    .B(_4884_),
    .C(_4883_),
    .Y(_4885_)
);

OR2X2 _11632_ (
    .A(_4882_),
    .B(_4880_),
    .Y(_4886_)
);

NAND2X1 _11633_ (
    .A(_4880_),
    .B(_4882_),
    .Y(_4887_)
);

NAND3X1 _11634_ (
    .A(_4513_),
    .B(_4887_),
    .C(_4886_),
    .Y(_4888_)
);

AND2X2 _11635_ (
    .A(_4885_),
    .B(_4888_),
    .Y(_4889_)
);

NAND2X1 _11636_ (
    .A(_4889_),
    .B(_4874_),
    .Y(_4890_)
);

INVX1 _11637_ (
    .A(_4842_),
    .Y(_4891_)
);

OAI21X1 _11638_ (
    .A(_4844_),
    .B(_4847_),
    .C(_4891_),
    .Y(_4892_)
);

INVX1 _11639_ (
    .A(_4865_),
    .Y(_4893_)
);

AOI21X1 _11640_ (
    .A(_4892_),
    .B(_4869_),
    .C(_4893_),
    .Y(_4894_)
);

NAND2X1 _11641_ (
    .A(_4888_),
    .B(_4885_),
    .Y(_4895_)
);

NAND2X1 _11642_ (
    .A(_4895_),
    .B(_4894_),
    .Y(_4896_)
);

NAND2X1 _11643_ (
    .A(_4890_),
    .B(_4896_),
    .Y(_4897_)
);

AOI22X1 _11644_ (
    .A(_4451_),
    .B(_4474__bF$buf0),
    .C(_4897_),
    .D(_4772_),
    .Y(_4348_)
);

NAND3X1 _11645_ (
    .A(_4859_),
    .B(_4881_),
    .C(_4863_),
    .Y(_4898_)
);

NOR2X1 _11646_ (
    .A(1'h0),
    .B(_4853_),
    .Y(_4899_)
);

NOR2X1 _11647_ (
    .A(_4480__bF$buf0),
    .B(_4760_),
    .Y(_4900_)
);

OAI21X1 _11648_ (
    .A(_4900_),
    .B(_4899_),
    .C(1'h1),
    .Y(_4901_)
);

OAI21X1 _11649_ (
    .A(1'h1),
    .B(_4807_),
    .C(_4901_),
    .Y(_4902_)
);

NAND3X1 _11650_ (
    .A(_4569__bF$buf2),
    .B(_4902_),
    .C(_4898_),
    .Y(_4903_)
);

INVX1 _11651_ (
    .A(_4902_),
    .Y(_4904_)
);

NAND3X1 _11652_ (
    .A(_4832_),
    .B(_4859_),
    .C(_4837_),
    .Y(_4905_)
);

OAI21X1 _11653_ (
    .A(_4880_),
    .B(_4905_),
    .C(_4569__bF$buf1),
    .Y(_4906_)
);

NAND2X1 _11654_ (
    .A(_4904_),
    .B(_4906_),
    .Y(_4907_)
);

NAND3X1 _11655_ (
    .A(\genblk1[5].u_ce.Xin12b [5]),
    .B(_4907_),
    .C(_4903_),
    .Y(_4908_)
);

NAND3X1 _11656_ (
    .A(_4569__bF$buf0),
    .B(_4904_),
    .C(_4898_),
    .Y(_4909_)
);

NAND2X1 _11657_ (
    .A(_4902_),
    .B(_4906_),
    .Y(_4910_)
);

NAND3X1 _11658_ (
    .A(_4521_),
    .B(_4910_),
    .C(_4909_),
    .Y(_4911_)
);

NAND2X1 _11659_ (
    .A(_4908_),
    .B(_4911_),
    .Y(_4912_)
);

AOI21X1 _11660_ (
    .A(_4890_),
    .B(_4885_),
    .C(_4912_),
    .Y(_4913_)
);

OAI21X1 _11661_ (
    .A(_4895_),
    .B(_4894_),
    .C(_4885_),
    .Y(_4914_)
);

AND2X2 _11662_ (
    .A(_4908_),
    .B(_4911_),
    .Y(_4915_)
);

OAI21X1 _11663_ (
    .A(_4915_),
    .B(_4914_),
    .C(_4772_),
    .Y(_4916_)
);

OAI22X1 _11664_ (
    .A(_4466_),
    .B(\genblk1[5].u_ce.Vld_bF$buf2 ),
    .C(_4913_),
    .D(_4916_),
    .Y(_4349_)
);

NOR2X1 _11665_ (
    .A(_4880_),
    .B(_4905_),
    .Y(_4917_)
);

NAND2X1 _11666_ (
    .A(_4904_),
    .B(_4917_),
    .Y(_4918_)
);

AOI21X1 _11667_ (
    .A(_4480__bF$buf4),
    .B(_4876_),
    .C(_4900_),
    .Y(_4919_)
);

NAND2X1 _11668_ (
    .A(_4507__bF$buf3),
    .B(_4827_),
    .Y(_4920_)
);

OAI21X1 _11669_ (
    .A(_4507__bF$buf2),
    .B(_4919_),
    .C(_4920_),
    .Y(_4921_)
);

NAND3X1 _11670_ (
    .A(_4569__bF$buf5),
    .B(_4921_),
    .C(_4918_),
    .Y(_4922_)
);

NOR3X1 _11671_ (
    .A(_4880_),
    .B(_4902_),
    .C(_4905_),
    .Y(_4923_)
);

INVX1 _11672_ (
    .A(_4921_),
    .Y(_4924_)
);

OAI21X1 _11673_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_4923_),
    .C(_4924_),
    .Y(_4925_)
);

NAND3X1 _11674_ (
    .A(\genblk1[5].u_ce.Xin12b [6]),
    .B(_4925_),
    .C(_4922_),
    .Y(_4926_)
);

NAND3X1 _11675_ (
    .A(_4569__bF$buf4),
    .B(_4924_),
    .C(_4918_),
    .Y(_4927_)
);

OAI21X1 _11676_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .B(_4923_),
    .C(_4921_),
    .Y(_4928_)
);

NAND3X1 _11677_ (
    .A(_4523_),
    .B(_4928_),
    .C(_4927_),
    .Y(_4929_)
);

AND2X2 _11678_ (
    .A(_4926_),
    .B(_4929_),
    .Y(_4930_)
);

NAND2X1 _11679_ (
    .A(_4889_),
    .B(_4915_),
    .Y(_4931_)
);

INVX1 _11680_ (
    .A(_4885_),
    .Y(_4932_)
);

INVX1 _11681_ (
    .A(_4908_),
    .Y(_4933_)
);

AOI21X1 _11682_ (
    .A(_4932_),
    .B(_4911_),
    .C(_4933_),
    .Y(_4934_)
);

OAI21X1 _11683_ (
    .A(_4894_),
    .B(_4931_),
    .C(_4934_),
    .Y(_4935_)
);

AND2X2 _11684_ (
    .A(_4935_),
    .B(_4930_),
    .Y(_4936_)
);

NOR2X1 _11685_ (
    .A(_4930_),
    .B(_4935_),
    .Y(_4937_)
);

OAI21X1 _11686_ (
    .A(_4937_),
    .B(_4936_),
    .C(_4478_),
    .Y(_4938_)
);

NAND2X1 _11687_ (
    .A(\genblk1[5].u_ce.Vld_bF$buf1 ),
    .B(_4938_),
    .Y(_4939_)
);

OAI21X1 _11688_ (
    .A(_4452_),
    .B(\genblk1[5].u_ce.Vld_bF$buf0 ),
    .C(_4939_),
    .Y(_4350_)
);

INVX1 _11689_ (
    .A(_4926_),
    .Y(_4940_)
);

NOR2X1 _11690_ (
    .A(_4940_),
    .B(_4936_),
    .Y(_4941_)
);

NAND2X1 _11691_ (
    .A(_4924_),
    .B(_4923_),
    .Y(_4942_)
);

NOR2X1 _11692_ (
    .A(_4507__bF$buf1),
    .B(_4760_),
    .Y(_4943_)
);

AOI21X1 _11693_ (
    .A(_4855_),
    .B(_4507__bF$buf0),
    .C(_4943_),
    .Y(_4944_)
);

NAND3X1 _11694_ (
    .A(_4569__bF$buf3),
    .B(_4944_),
    .C(_4942_),
    .Y(_4945_)
);

INVX1 _11695_ (
    .A(_4945_),
    .Y(_4946_)
);

AOI21X1 _11696_ (
    .A(_4942_),
    .B(_4569__bF$buf2),
    .C(_4944_),
    .Y(_4947_)
);

OAI21X1 _11697_ (
    .A(_4947_),
    .B(_4946_),
    .C(\genblk1[5].u_ce.Xin12b [7]),
    .Y(_4948_)
);

INVX1 _11698_ (
    .A(_4947_),
    .Y(_4949_)
);

NAND3X1 _11699_ (
    .A(_4526_),
    .B(_4945_),
    .C(_4949_),
    .Y(_4950_)
);

AND2X2 _11700_ (
    .A(_4950_),
    .B(_4948_),
    .Y(_4951_)
);

OR2X2 _11701_ (
    .A(_4941_),
    .B(_4951_),
    .Y(_4952_)
);

AOI21X1 _11702_ (
    .A(_4941_),
    .B(_4951_),
    .C(_4771_),
    .Y(_4953_)
);

AOI22X1 _11703_ (
    .A(_4465_),
    .B(_4474__bF$buf4),
    .C(_4952_),
    .D(_4953_),
    .Y(_4351_)
);

NOR2X1 _11704_ (
    .A(_4895_),
    .B(_4912_),
    .Y(_4954_)
);

OAI21X1 _11705_ (
    .A(_4885_),
    .B(_4912_),
    .C(_4908_),
    .Y(_4955_)
);

AOI21X1 _11706_ (
    .A(_4954_),
    .B(_4874_),
    .C(_4955_),
    .Y(_4956_)
);

AOI21X1 _11707_ (
    .A(_4949_),
    .B(_4945_),
    .C(_4526_),
    .Y(_4957_)
);

AOI21X1 _11708_ (
    .A(_4940_),
    .B(_4950_),
    .C(_4957_),
    .Y(_4958_)
);

NAND3X1 _11709_ (
    .A(_4930_),
    .B(_4948_),
    .C(_4950_),
    .Y(_4959_)
);

OAI21X1 _11710_ (
    .A(_4959_),
    .B(_4956_),
    .C(_4958_),
    .Y(_4960_)
);

NAND3X1 _11711_ (
    .A(_4924_),
    .B(_4944_),
    .C(_4923_),
    .Y(_4961_)
);

INVX1 _11712_ (
    .A(_4878_),
    .Y(_4962_)
);

INVX1 _11713_ (
    .A(_4943_),
    .Y(_4963_)
);

OAI21X1 _11714_ (
    .A(1'h1),
    .B(_4962_),
    .C(_4963_),
    .Y(_4964_)
);

INVX1 _11715_ (
    .A(_4964_),
    .Y(_4965_)
);

NAND3X1 _11716_ (
    .A(_4569__bF$buf1),
    .B(_4965_),
    .C(_4961_),
    .Y(_4966_)
);

INVX1 _11717_ (
    .A(_4966_),
    .Y(_4967_)
);

AOI21X1 _11718_ (
    .A(_4961_),
    .B(_4569__bF$buf0),
    .C(_4965_),
    .Y(_4968_)
);

OAI21X1 _11719_ (
    .A(_4968_),
    .B(_4967_),
    .C(\genblk1[5].u_ce.Xin12b [8]),
    .Y(_4969_)
);

INVX1 _11720_ (
    .A(_4968_),
    .Y(_4970_)
);

NAND3X1 _11721_ (
    .A(_4528_),
    .B(_4966_),
    .C(_4970_),
    .Y(_4971_)
);

AND2X2 _11722_ (
    .A(_4971_),
    .B(_4969_),
    .Y(_4972_)
);

OR2X2 _11723_ (
    .A(_4960_),
    .B(_4972_),
    .Y(_4973_)
);

INVX1 _11724_ (
    .A(_4973_),
    .Y(_4974_)
);

NAND2X1 _11725_ (
    .A(_4972_),
    .B(_4960_),
    .Y(_4975_)
);

NAND2X1 _11726_ (
    .A(_4772_),
    .B(_4975_),
    .Y(_4976_)
);

OAI22X1 _11727_ (
    .A(_4454_),
    .B(\genblk1[5].u_ce.Vld_bF$buf3 ),
    .C(_4976_),
    .D(_4974_),
    .Y(_4352_)
);

NOR3X1 _11728_ (
    .A(_4902_),
    .B(_4921_),
    .C(_4898_),
    .Y(_4977_)
);

NAND3X1 _11729_ (
    .A(_4944_),
    .B(_4965_),
    .C(_4977_),
    .Y(_4978_)
);

OR2X2 _11730_ (
    .A(_4899_),
    .B(_4900_),
    .Y(_4979_)
);

AOI21X1 _11731_ (
    .A(_4979_),
    .B(_4507__bF$buf3),
    .C(_4943_),
    .Y(_4980_)
);

INVX1 _11732_ (
    .A(_4980_),
    .Y(_4981_)
);

NAND3X1 _11733_ (
    .A(_4569__bF$buf5),
    .B(_4981_),
    .C(_4978_),
    .Y(_4982_)
);

OAI21X1 _11734_ (
    .A(_4964_),
    .B(_4961_),
    .C(_4569__bF$buf4),
    .Y(_4983_)
);

NAND2X1 _11735_ (
    .A(_4980_),
    .B(_4983_),
    .Y(_4984_)
);

NAND3X1 _11736_ (
    .A(\genblk1[5].u_ce.Xin12b [9]),
    .B(_4984_),
    .C(_4982_),
    .Y(_4985_)
);

NAND3X1 _11737_ (
    .A(_4569__bF$buf3),
    .B(_4980_),
    .C(_4978_),
    .Y(_4986_)
);

NAND2X1 _11738_ (
    .A(_4981_),
    .B(_4983_),
    .Y(_4987_)
);

NAND3X1 _11739_ (
    .A(_4573_),
    .B(_4987_),
    .C(_4986_),
    .Y(_4988_)
);

NAND2X1 _11740_ (
    .A(_4985_),
    .B(_4988_),
    .Y(_4989_)
);

AOI21X1 _11741_ (
    .A(_4975_),
    .B(_4969_),
    .C(_4989_),
    .Y(_4990_)
);

NAND3X1 _11742_ (
    .A(_4969_),
    .B(_4989_),
    .C(_4975_),
    .Y(_4991_)
);

NAND2X1 _11743_ (
    .A(_4772_),
    .B(_4991_),
    .Y(_4992_)
);

OAI22X1 _11744_ (
    .A(_4462_),
    .B(\genblk1[5].u_ce.Vld_bF$buf2 ),
    .C(_4990_),
    .D(_4992_),
    .Y(_4353_)
);

NAND2X1 _11745_ (
    .A(\genblk1[5].u_ce.Xcalc [10]),
    .B(_4474__bF$buf3),
    .Y(_4993_)
);

OAI21X1 _11746_ (
    .A(1'h1),
    .B(_4919_),
    .C(_4963_),
    .Y(_4994_)
);

OAI21X1 _11747_ (
    .A(_4981_),
    .B(_4978_),
    .C(_4569__bF$buf2),
    .Y(_4995_)
);

NOR2X1 _11748_ (
    .A(_4994_),
    .B(_4995_),
    .Y(_4996_)
);

NAND2X1 _11749_ (
    .A(_4994_),
    .B(_4995_),
    .Y(_4997_)
);

INVX1 _11750_ (
    .A(_4997_),
    .Y(_4998_)
);

OAI21X1 _11751_ (
    .A(_4996_),
    .B(_4998_),
    .C(\genblk1[5].u_ce.Xin12b [10]),
    .Y(_4999_)
);

INVX1 _11752_ (
    .A(_4996_),
    .Y(_5000_)
);

NAND3X1 _11753_ (
    .A(_4603_),
    .B(_4997_),
    .C(_5000_),
    .Y(_5001_)
);

AND2X2 _11754_ (
    .A(_5001_),
    .B(_4999_),
    .Y(_5002_)
);

OAI21X1 _11755_ (
    .A(_4969_),
    .B(_4989_),
    .C(_4985_),
    .Y(_5003_)
);

NAND3X1 _11756_ (
    .A(_4930_),
    .B(_4935_),
    .C(_4951_),
    .Y(_5004_)
);

NAND3X1 _11757_ (
    .A(_4985_),
    .B(_4988_),
    .C(_4972_),
    .Y(_5005_)
);

AOI21X1 _11758_ (
    .A(_5004_),
    .B(_4958_),
    .C(_5005_),
    .Y(_5006_)
);

OAI21X1 _11759_ (
    .A(_5003_),
    .B(_5006_),
    .C(_5002_),
    .Y(_5007_)
);

NAND2X1 _11760_ (
    .A(_4999_),
    .B(_5001_),
    .Y(_5008_)
);

NAND2X1 _11761_ (
    .A(_4969_),
    .B(_4971_),
    .Y(_5009_)
);

NOR2X1 _11762_ (
    .A(_5009_),
    .B(_4989_),
    .Y(_5010_)
);

AOI21X1 _11763_ (
    .A(_4960_),
    .B(_5010_),
    .C(_5003_),
    .Y(_5011_)
);

NAND2X1 _11764_ (
    .A(_5008_),
    .B(_5011_),
    .Y(_5012_)
);

AOI21X1 _11765_ (
    .A(_5007_),
    .B(_5012_),
    .C(_4479_),
    .Y(_5013_)
);

OAI21X1 _11766_ (
    .A(_4474__bF$buf2),
    .B(_5013_),
    .C(_4993_),
    .Y(_4354_)
);

NAND2X1 _11767_ (
    .A(\genblk1[5].u_ce.Xcalc [11]),
    .B(_4474__bF$buf1),
    .Y(_5014_)
);

OR2X2 _11768_ (
    .A(_4978_),
    .B(_4981_),
    .Y(_5015_)
);

OAI21X1 _11769_ (
    .A(_4994_),
    .B(_5015_),
    .C(_4569__bF$buf1),
    .Y(_5016_)
);

OR2X2 _11770_ (
    .A(_5016_),
    .B(_4762_),
    .Y(_5017_)
);

NAND2X1 _11771_ (
    .A(_4762_),
    .B(_5016_),
    .Y(_5018_)
);

AOI22X1 _11772_ (
    .A(_5017_),
    .B(_5018_),
    .C(_5007_),
    .D(_4999_),
    .Y(_5019_)
);

OAI21X1 _11773_ (
    .A(_5008_),
    .B(_5011_),
    .C(_4999_),
    .Y(_5020_)
);

NAND2X1 _11774_ (
    .A(_5018_),
    .B(_5017_),
    .Y(_5021_)
);

OAI21X1 _11775_ (
    .A(_5021_),
    .B(_5020_),
    .C(_4772_),
    .Y(_5022_)
);

OAI21X1 _11776_ (
    .A(_5019_),
    .B(_5022_),
    .C(_5014_),
    .Y(_4355_)
);

NAND2X1 _11777_ (
    .A(1'h1),
    .B(1'h0),
    .Y(_5023_)
);

OAI21X1 _11778_ (
    .A(_4507__bF$buf2),
    .B(_4689_),
    .C(_5023_),
    .Y(_5024_)
);

NOR2X1 _11779_ (
    .A(_4470_),
    .B(_5024_),
    .Y(_5025_)
);

NAND2X1 _11780_ (
    .A(\genblk1[5].u_ce.Acalc [1]),
    .B(_4474__bF$buf0),
    .Y(_5026_)
);

OAI21X1 _11781_ (
    .A(1'h0),
    .B(_4476_),
    .C(1'h1),
    .Y(_5027_)
);

OAI21X1 _11782_ (
    .A(1'h1),
    .B(_4476_),
    .C(_5027_),
    .Y(_5028_)
);

OAI21X1 _11783_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5024_),
    .C(_5028_),
    .Y(_5029_)
);

OAI21X1 _11784_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf4 ),
    .B(_5028_),
    .C(_5029_),
    .Y(_5030_)
);

OR2X2 _11785_ (
    .A(_5030_),
    .B(\genblk1[5].u_ce.Ain0 [1]),
    .Y(_5031_)
);

NAND2X1 _11786_ (
    .A(\genblk1[5].u_ce.Ain0 [1]),
    .B(_5030_),
    .Y(_5032_)
);

NAND2X1 _11787_ (
    .A(_5032_),
    .B(_5031_),
    .Y(_5033_)
);

NOR2X1 _11788_ (
    .A(_5025_),
    .B(_5033_),
    .Y(_5034_)
);

NAND2X1 _11789_ (
    .A(_5025_),
    .B(_5033_),
    .Y(_5035_)
);

NAND2X1 _11790_ (
    .A(\genblk1[5].u_ce.Vld_bF$buf1 ),
    .B(_5035_),
    .Y(_5036_)
);

OAI21X1 _11791_ (
    .A(_5034_),
    .B(_5036_),
    .C(_5026_),
    .Y(_4356_)
);

OAI21X1 _11792_ (
    .A(_4472_),
    .B(_5030_),
    .C(_5035_),
    .Y(_5037_)
);

OAI21X1 _11793_ (
    .A(_4476_),
    .B(_4480__bF$buf3),
    .C(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_5038_)
);

NAND3X1 _11794_ (
    .A(1'h1),
    .B(_4689_),
    .C(_5038_),
    .Y(_5039_)
);

OAI21X1 _11795_ (
    .A(1'h1),
    .B(_5038_),
    .C(_5039_),
    .Y(_5040_)
);

NAND2X1 _11796_ (
    .A(\genblk1[5].u_ce.Ain1 [0]),
    .B(_5040_),
    .Y(_5041_)
);

OR2X2 _11797_ (
    .A(_5040_),
    .B(\genblk1[5].u_ce.Ain1 [0]),
    .Y(_5042_)
);

NAND2X1 _11798_ (
    .A(_5041_),
    .B(_5042_),
    .Y(_5043_)
);

INVX1 _11799_ (
    .A(_5043_),
    .Y(_5044_)
);

NAND2X1 _11800_ (
    .A(_5044_),
    .B(_5037_),
    .Y(_5045_)
);

NAND2X1 _11801_ (
    .A(_5041_),
    .B(_5045_),
    .Y(_5046_)
);

INVX1 _11802_ (
    .A(_5046_),
    .Y(_5047_)
);

INVX1 _11803_ (
    .A(\genblk1[5].u_ce.Ain1 [1]),
    .Y(_5048_)
);

OAI21X1 _11804_ (
    .A(1'h1),
    .B(_4480__bF$buf2),
    .C(1'h1),
    .Y(_5049_)
);

NAND2X1 _11805_ (
    .A(_4569__bF$buf0),
    .B(_5049_),
    .Y(_5050_)
);

OAI21X1 _11806_ (
    .A(1'h1),
    .B(1'h0),
    .C(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .Y(_5051_)
);

OAI21X1 _11807_ (
    .A(_4476_),
    .B(_5051_),
    .C(_5050_),
    .Y(_5052_)
);

NOR2X1 _11808_ (
    .A(_5048_),
    .B(_5052_),
    .Y(_5053_)
);

NAND2X1 _11809_ (
    .A(_5048_),
    .B(_5052_),
    .Y(_5054_)
);

INVX1 _11810_ (
    .A(_5054_),
    .Y(_5055_)
);

OAI21X1 _11811_ (
    .A(_5053_),
    .B(_5055_),
    .C(_5047_),
    .Y(_5056_)
);

INVX1 _11812_ (
    .A(_5053_),
    .Y(_5057_)
);

NAND3X1 _11813_ (
    .A(_5057_),
    .B(_5054_),
    .C(_5046_),
    .Y(_5058_)
);

NAND2X1 _11814_ (
    .A(_5058_),
    .B(_5056_),
    .Y(_5059_)
);

NAND2X1 _11815_ (
    .A(\genblk1[5].u_ce.Acalc [3]),
    .B(_4474__bF$buf4),
    .Y(_5060_)
);

OAI21X1 _11816_ (
    .A(_4474__bF$buf3),
    .B(_5059_),
    .C(_5060_),
    .Y(_4357_)
);

NOR2X1 _11817_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf1 ),
    .B(_5028_),
    .Y(_5061_)
);

NAND3X1 _11818_ (
    .A(1'h1),
    .B(_4507__bF$buf1),
    .C(_4480__bF$buf1),
    .Y(_5062_)
);

AOI21X1 _11819_ (
    .A(_5027_),
    .B(_5062_),
    .C(_4569__bF$buf5),
    .Y(_5063_)
);

NOR2X1 _11820_ (
    .A(_5063_),
    .B(_5061_),
    .Y(_5064_)
);

NAND2X1 _11821_ (
    .A(\genblk1[5].u_ce.Ain12b [4]),
    .B(_5064_),
    .Y(_5065_)
);

INVX1 _11822_ (
    .A(\genblk1[5].u_ce.Ain12b [4]),
    .Y(_5066_)
);

OAI21X1 _11823_ (
    .A(_5063_),
    .B(_5061_),
    .C(_5066_),
    .Y(_5067_)
);

NAND2X1 _11824_ (
    .A(_5067_),
    .B(_5065_),
    .Y(_5068_)
);

AOI21X1 _11825_ (
    .A(_5046_),
    .B(_5054_),
    .C(_5053_),
    .Y(_5069_)
);

NAND2X1 _11826_ (
    .A(\genblk1[5].u_ce.Acalc [5]),
    .B(_4474__bF$buf2),
    .Y(_5070_)
);

OAI21X1 _11827_ (
    .A(_5068_),
    .B(_5069_),
    .C(_5065_),
    .Y(_5071_)
);

OAI21X1 _11828_ (
    .A(1'h1),
    .B(1'h0),
    .C(_4508_),
    .Y(_5072_)
);

NAND2X1 _11829_ (
    .A(_4569__bF$buf4),
    .B(_5072_),
    .Y(_5073_)
);

INVX1 _11830_ (
    .A(_5073_),
    .Y(_5074_)
);

NOR2X1 _11831_ (
    .A(_4569__bF$buf3),
    .B(_5072_),
    .Y(_5075_)
);

NOR2X1 _11832_ (
    .A(_5075_),
    .B(_5074_),
    .Y(_5076_)
);

NAND2X1 _11833_ (
    .A(\genblk1[5].u_ce.Ain12b [5]),
    .B(_5076_),
    .Y(_5077_)
);

INVX1 _11834_ (
    .A(\genblk1[5].u_ce.Ain12b [5]),
    .Y(_5078_)
);

OAI21X1 _11835_ (
    .A(_5075_),
    .B(_5074_),
    .C(_5078_),
    .Y(_5079_)
);

NAND2X1 _11836_ (
    .A(_5079_),
    .B(_5077_),
    .Y(_5080_)
);

INVX1 _11837_ (
    .A(_5080_),
    .Y(_5081_)
);

NOR2X1 _11838_ (
    .A(_5081_),
    .B(_5071_),
    .Y(_5082_)
);

NAND2X1 _11839_ (
    .A(_5081_),
    .B(_5071_),
    .Y(_5083_)
);

NAND2X1 _11840_ (
    .A(\genblk1[5].u_ce.Vld_bF$buf0 ),
    .B(_5083_),
    .Y(_5084_)
);

OAI21X1 _11841_ (
    .A(_5082_),
    .B(_5084_),
    .C(_5070_),
    .Y(_4358_)
);

INVX1 _11842_ (
    .A(_5069_),
    .Y(_5085_)
);

NOR2X1 _11843_ (
    .A(_5068_),
    .B(_5080_),
    .Y(_5086_)
);

OAI21X1 _11844_ (
    .A(_5065_),
    .B(_5080_),
    .C(_5077_),
    .Y(_5087_)
);

AOI21X1 _11845_ (
    .A(_5085_),
    .B(_5086_),
    .C(_5087_),
    .Y(_5088_)
);

OAI21X1 _11846_ (
    .A(1'h1),
    .B(_5023_),
    .C(_4478_),
    .Y(_5089_)
);

NOR2X1 _11847_ (
    .A(_4569__bF$buf2),
    .B(_5089_),
    .Y(_5090_)
);

NAND2X1 _11848_ (
    .A(_4569__bF$buf1),
    .B(_5089_),
    .Y(_5091_)
);

INVX1 _11849_ (
    .A(_5091_),
    .Y(_5092_)
);

NOR2X1 _11850_ (
    .A(_5090_),
    .B(_5092_),
    .Y(_5093_)
);

NAND2X1 _11851_ (
    .A(\genblk1[5].u_ce.Ain12b [6]),
    .B(_5093_),
    .Y(_5094_)
);

OR2X2 _11852_ (
    .A(_5093_),
    .B(\genblk1[5].u_ce.Ain12b [6]),
    .Y(_5095_)
);

AND2X2 _11853_ (
    .A(_5095_),
    .B(_5094_),
    .Y(_5096_)
);

INVX1 _11854_ (
    .A(_5096_),
    .Y(_5097_)
);

OAI21X1 _11855_ (
    .A(_5097_),
    .B(_5088_),
    .C(_5094_),
    .Y(_5098_)
);

OAI21X1 _11856_ (
    .A(1'h1),
    .B(1'h1),
    .C(\genblk1[5].u_ce.Ain12b_11_bF$buf0 ),
    .Y(_5099_)
);

NAND2X1 _11857_ (
    .A(_5099_),
    .B(_4570_),
    .Y(_5100_)
);

INVX1 _11858_ (
    .A(_5100_),
    .Y(_5101_)
);

NAND2X1 _11859_ (
    .A(\genblk1[5].u_ce.Ain12b [7]),
    .B(_5101_),
    .Y(_5102_)
);

INVX1 _11860_ (
    .A(_5102_),
    .Y(_5103_)
);

NOR2X1 _11861_ (
    .A(\genblk1[5].u_ce.Ain12b [7]),
    .B(_5101_),
    .Y(_5104_)
);

NOR2X1 _11862_ (
    .A(_5104_),
    .B(_5103_),
    .Y(_5105_)
);

INVX1 _11863_ (
    .A(_5105_),
    .Y(_5106_)
);

OR2X2 _11864_ (
    .A(_5098_),
    .B(_5106_),
    .Y(_5107_)
);

AOI21X1 _11865_ (
    .A(_5098_),
    .B(_5106_),
    .C(_4474__bF$buf1),
    .Y(_5108_)
);

AOI22X1 _11866_ (
    .A(_4427_),
    .B(_4474__bF$buf0),
    .C(_5107_),
    .D(_5108_),
    .Y(_4359_)
);

OAI21X1 _11867_ (
    .A(_5104_),
    .B(_5094_),
    .C(_5102_),
    .Y(_5109_)
);

NAND2X1 _11868_ (
    .A(_5105_),
    .B(_5096_),
    .Y(_5110_)
);

INVX1 _11869_ (
    .A(_5110_),
    .Y(_5111_)
);

AOI21X1 _11870_ (
    .A(_5111_),
    .B(_5087_),
    .C(_5109_),
    .Y(_5112_)
);

NAND2X1 _11871_ (
    .A(_5086_),
    .B(_5111_),
    .Y(_5113_)
);

OAI21X1 _11872_ (
    .A(_5113_),
    .B(_5069_),
    .C(_5112_),
    .Y(_5114_)
);

INVX1 _11873_ (
    .A(\genblk1[5].u_ce.Ain12b [8]),
    .Y(_5115_)
);

NAND2X1 _11874_ (
    .A(_4569__bF$buf0),
    .B(_4477_),
    .Y(_5116_)
);

NAND2X1 _11875_ (
    .A(_5051_),
    .B(_5116_),
    .Y(_5117_)
);

OR2X2 _11876_ (
    .A(_5117_),
    .B(_5115_),
    .Y(_5118_)
);

NAND2X1 _11877_ (
    .A(_5115_),
    .B(_5117_),
    .Y(_5119_)
);

AND2X2 _11878_ (
    .A(_5118_),
    .B(_5119_),
    .Y(_5120_)
);

NAND2X1 _11879_ (
    .A(_5120_),
    .B(_5114_),
    .Y(_5121_)
);

NAND2X1 _11880_ (
    .A(\genblk1[5].u_ce.Acalc [9]),
    .B(_4474__bF$buf4),
    .Y(_5122_)
);

OAI21X1 _11881_ (
    .A(_5115_),
    .B(_5117_),
    .C(_5121_),
    .Y(_5123_)
);

INVX1 _11882_ (
    .A(\genblk1[5].u_ce.Ain12b [9]),
    .Y(_5124_)
);

NAND2X1 _11883_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf4 ),
    .B(_5124_),
    .Y(_5125_)
);

NOR2X1 _11884_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf3 ),
    .B(_5124_),
    .Y(_5126_)
);

INVX1 _11885_ (
    .A(_5126_),
    .Y(_5127_)
);

NAND2X1 _11886_ (
    .A(_5125_),
    .B(_5127_),
    .Y(_5128_)
);

INVX1 _11887_ (
    .A(_5128_),
    .Y(_5129_)
);

NOR2X1 _11888_ (
    .A(_5129_),
    .B(_5123_),
    .Y(_5130_)
);

NAND2X1 _11889_ (
    .A(_5129_),
    .B(_5123_),
    .Y(_5131_)
);

NAND2X1 _11890_ (
    .A(\genblk1[5].u_ce.Vld_bF$buf3 ),
    .B(_5131_),
    .Y(_5132_)
);

OAI21X1 _11891_ (
    .A(_5130_),
    .B(_5132_),
    .C(_5122_),
    .Y(_4360_)
);

AOI21X1 _11892_ (
    .A(_5123_),
    .B(_5125_),
    .C(_5126_),
    .Y(_5133_)
);

INVX1 _11893_ (
    .A(\genblk1[5].u_ce.Ain12b [10]),
    .Y(_5134_)
);

NAND2X1 _11894_ (
    .A(\genblk1[5].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5134_),
    .Y(_5135_)
);

NAND2X1 _11895_ (
    .A(\genblk1[5].u_ce.Ain12b [10]),
    .B(_4569__bF$buf5),
    .Y(_5136_)
);

NAND2X1 _11896_ (
    .A(_5135_),
    .B(_5136_),
    .Y(_5137_)
);

NAND2X1 _11897_ (
    .A(\genblk1[5].u_ce.Acalc [11]),
    .B(_4474__bF$buf3),
    .Y(_5138_)
);

OAI21X1 _11898_ (
    .A(_5137_),
    .B(_5133_),
    .C(_5136_),
    .Y(_5139_)
);

OAI21X1 _11899_ (
    .A(_4474__bF$buf2),
    .B(_5139_),
    .C(_5138_),
    .Y(_4361_)
);

INVX1 _11900_ (
    .A(_4416_),
    .Y(_5140_)
);

NAND3X1 _11901_ (
    .A(_4461_),
    .B(\genblk1[5].u_ce.LoadCtl [5]),
    .C(_4420_),
    .Y(_5141_)
);

NOR2X1 _11902_ (
    .A(_5140_),
    .B(_5141_),
    .Y(_5142_)
);

NAND2X1 _11903_ (
    .A(\genblk1[4].u_ce.X_ [0]),
    .B(_5142_),
    .Y(_5143_)
);

OAI21X1 _11904_ (
    .A(_4603_),
    .B(_5142_),
    .C(_5143_),
    .Y(_4362_)
);

NAND2X1 _11905_ (
    .A(\genblk1[4].u_ce.X_ [1]),
    .B(_5142_),
    .Y(_5144_)
);

OAI21X1 _11906_ (
    .A(_4628_),
    .B(_5142_),
    .C(_5144_),
    .Y(_4363_)
);

INVX1 _11907_ (
    .A(\genblk1[4].u_ce.X_ [0]),
    .Y(_5145_)
);

NAND3X1 _11908_ (
    .A(\genblk1[5].u_ce.LoadCtl [4]),
    .B(_4416_),
    .C(_4420_),
    .Y(_5146_)
);

NAND2X1 _11909_ (
    .A(\genblk1[5].u_ce.Xin12b [8]),
    .B(_5146_),
    .Y(_5147_)
);

OAI21X1 _11910_ (
    .A(_5145_),
    .B(_5146_),
    .C(_5147_),
    .Y(_4364_)
);

INVX1 _11911_ (
    .A(\genblk1[4].u_ce.X_ [1]),
    .Y(_5148_)
);

NAND2X1 _11912_ (
    .A(\genblk1[5].u_ce.Xin12b [9]),
    .B(_5146_),
    .Y(_5149_)
);

OAI21X1 _11913_ (
    .A(_5148_),
    .B(_5146_),
    .C(_5149_),
    .Y(_4365_)
);

NAND2X1 _11914_ (
    .A(_4420_),
    .B(_4419_),
    .Y(_5150_)
);

OAI21X1 _11915_ (
    .A(_4421_),
    .B(_4428_),
    .C(\genblk1[5].u_ce.Xin12b [6]),
    .Y(_5151_)
);

OAI21X1 _11916_ (
    .A(_5145_),
    .B(_5150_),
    .C(_5151_),
    .Y(_4366_)
);

OAI21X1 _11917_ (
    .A(_4421_),
    .B(_4428_),
    .C(\genblk1[5].u_ce.Xin12b [7]),
    .Y(_5152_)
);

OAI21X1 _11918_ (
    .A(_5148_),
    .B(_5150_),
    .C(_5152_),
    .Y(_4367_)
);

NOR2X1 _11919_ (
    .A(_4417_),
    .B(_4421_),
    .Y(_5153_)
);

NAND2X1 _11920_ (
    .A(\genblk1[4].u_ce.X_ [0]),
    .B(_5153_),
    .Y(_5154_)
);

OAI21X1 _11921_ (
    .A(_4513_),
    .B(_5153_),
    .C(_5154_),
    .Y(_4368_)
);

NAND2X1 _11922_ (
    .A(\genblk1[4].u_ce.X_ [1]),
    .B(_5153_),
    .Y(_5155_)
);

OAI21X1 _11923_ (
    .A(_4521_),
    .B(_5153_),
    .C(_5155_),
    .Y(_4369_)
);

OAI21X1 _11924_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_4422_),
    .C(\genblk1[5].u_ce.Xin1 [0]),
    .Y(_5156_)
);

OAI21X1 _11925_ (
    .A(_5145_),
    .B(_4450_),
    .C(_5156_),
    .Y(_4370_)
);

OAI21X1 _11926_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_4422_),
    .C(\genblk1[5].u_ce.Xin1 [1]),
    .Y(_5157_)
);

OAI21X1 _11927_ (
    .A(_5148_),
    .B(_4450_),
    .C(_5157_),
    .Y(_4371_)
);

NAND2X1 _11928_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[4].u_ce.X_ [0]),
    .Y(_5158_)
);

OAI21X1 _11929_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_4536_),
    .C(_5158_),
    .Y(_4372_)
);

NAND2X1 _11930_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[4].u_ce.X_ [1]),
    .Y(_5159_)
);

OAI21X1 _11931_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_4516_),
    .C(_5159_),
    .Y(_4373_)
);

NAND2X1 _11932_ (
    .A(\genblk1[4].u_ce.Y_ [0]),
    .B(_5142_),
    .Y(_5160_)
);

OAI21X1 _11933_ (
    .A(_4736_),
    .B(_5142_),
    .C(_5160_),
    .Y(_4374_)
);

NAND2X1 _11934_ (
    .A(\genblk1[4].u_ce.Y_ [1]),
    .B(_5142_),
    .Y(_5161_)
);

OAI21X1 _11935_ (
    .A(_4760_),
    .B(_5142_),
    .C(_5161_),
    .Y(_4375_)
);

INVX1 _11936_ (
    .A(\genblk1[4].u_ce.Y_ [0]),
    .Y(_5162_)
);

NAND2X1 _11937_ (
    .A(\genblk1[5].u_ce.Yin12b [8]),
    .B(_5146_),
    .Y(_5163_)
);

OAI21X1 _11938_ (
    .A(_5162_),
    .B(_5146_),
    .C(_5163_),
    .Y(_4376_)
);

INVX1 _11939_ (
    .A(\genblk1[4].u_ce.Y_ [1]),
    .Y(_5164_)
);

NAND2X1 _11940_ (
    .A(\genblk1[5].u_ce.Yin12b [9]),
    .B(_5146_),
    .Y(_5165_)
);

OAI21X1 _11941_ (
    .A(_5164_),
    .B(_5146_),
    .C(_5165_),
    .Y(_4377_)
);

OAI21X1 _11942_ (
    .A(_4421_),
    .B(_4428_),
    .C(\genblk1[5].u_ce.Yin12b [6]),
    .Y(_4396_)
);

OAI21X1 _11943_ (
    .A(_5162_),
    .B(_5150_),
    .C(_4396_),
    .Y(_4378_)
);

OAI21X1 _11944_ (
    .A(_4421_),
    .B(_4428_),
    .C(\genblk1[5].u_ce.Yin12b [7]),
    .Y(_4397_)
);

OAI21X1 _11945_ (
    .A(_5164_),
    .B(_5150_),
    .C(_4397_),
    .Y(_4379_)
);

NAND2X1 _11946_ (
    .A(\genblk1[4].u_ce.Y_ [0]),
    .B(_5153_),
    .Y(_4398_)
);

OAI21X1 _11947_ (
    .A(_4601_),
    .B(_5153_),
    .C(_4398_),
    .Y(_4380_)
);

NAND2X1 _11948_ (
    .A(\genblk1[4].u_ce.Y_ [1]),
    .B(_5153_),
    .Y(_4399_)
);

OAI21X1 _11949_ (
    .A(_4626_),
    .B(_5153_),
    .C(_4399_),
    .Y(_4381_)
);

OAI21X1 _11950_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_4422_),
    .C(\genblk1[5].u_ce.Yin1 [0]),
    .Y(_4400_)
);

OAI21X1 _11951_ (
    .A(_5162_),
    .B(_4450_),
    .C(_4400_),
    .Y(_4382_)
);

OAI21X1 _11952_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_4422_),
    .C(\genblk1[5].u_ce.Yin1 [1]),
    .Y(_4401_)
);

OAI21X1 _11953_ (
    .A(_5164_),
    .B(_4450_),
    .C(_4401_),
    .Y(_4383_)
);

NAND2X1 _11954_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[4].u_ce.Y_ [0]),
    .Y(_4402_)
);

OAI21X1 _11955_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_4773_),
    .C(_4402_),
    .Y(_4384_)
);

NAND2X1 _11956_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[4].u_ce.Y_ [1]),
    .Y(_4403_)
);

OAI21X1 _11957_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_4558_),
    .C(_4403_),
    .Y(_4385_)
);

NAND2X1 _11958_ (
    .A(\a[5] [0]),
    .B(_5142_),
    .Y(_4404_)
);

OAI21X1 _11959_ (
    .A(_5134_),
    .B(_5142_),
    .C(_4404_),
    .Y(_4386_)
);

NAND2X1 _11960_ (
    .A(\a[5] [1]),
    .B(_5142_),
    .Y(_4405_)
);

OAI21X1 _11961_ (
    .A(_4569__bF$buf4),
    .B(_5142_),
    .C(_4405_),
    .Y(_4387_)
);

INVX1 _11962_ (
    .A(\a[5] [0]),
    .Y(_4406_)
);

NAND2X1 _11963_ (
    .A(\genblk1[5].u_ce.Ain12b [8]),
    .B(_5146_),
    .Y(_4407_)
);

OAI21X1 _11964_ (
    .A(_4406_),
    .B(_5146_),
    .C(_4407_),
    .Y(_4388_)
);

INVX1 _11965_ (
    .A(\a[5] [1]),
    .Y(_4408_)
);

NAND2X1 _11966_ (
    .A(\genblk1[5].u_ce.Ain12b [9]),
    .B(_5146_),
    .Y(_4409_)
);

OAI21X1 _11967_ (
    .A(_4408_),
    .B(_5146_),
    .C(_4409_),
    .Y(_4389_)
);

OAI21X1 _11968_ (
    .A(_4421_),
    .B(_4428_),
    .C(\genblk1[5].u_ce.Ain12b [6]),
    .Y(_4410_)
);

OAI21X1 _11969_ (
    .A(_4406_),
    .B(_5150_),
    .C(_4410_),
    .Y(_4390_)
);

OAI21X1 _11970_ (
    .A(_4421_),
    .B(_4428_),
    .C(\genblk1[5].u_ce.Ain12b [7]),
    .Y(_4411_)
);

OAI21X1 _11971_ (
    .A(_4408_),
    .B(_5150_),
    .C(_4411_),
    .Y(_4391_)
);

NAND2X1 _11972_ (
    .A(\a[5] [0]),
    .B(_5153_),
    .Y(_4412_)
);

OAI21X1 _11973_ (
    .A(_5066_),
    .B(_5153_),
    .C(_4412_),
    .Y(_4392_)
);

NAND2X1 _11974_ (
    .A(\a[5] [1]),
    .B(_5153_),
    .Y(_4413_)
);

OAI21X1 _11975_ (
    .A(_5078_),
    .B(_5153_),
    .C(_4413_),
    .Y(_4393_)
);

OAI21X1 _11976_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_4422_),
    .C(\genblk1[5].u_ce.Ain1 [0]),
    .Y(_4414_)
);

OAI21X1 _11977_ (
    .A(_4406_),
    .B(_4450_),
    .C(_4414_),
    .Y(_4394_)
);

OAI21X1 _11978_ (
    .A(\genblk1[5].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_4422_),
    .C(\genblk1[5].u_ce.Ain1 [1]),
    .Y(_4415_)
);

OAI21X1 _11979_ (
    .A(_4408_),
    .B(_4450_),
    .C(_4415_),
    .Y(_4395_)
);

DFFPOSX1 _11980_ (
    .CLK(clk_bF$buf55),
    .D(_4330_),
    .Q(\genblk1[5].u_ce.Ain0 [0])
);

DFFPOSX1 _11981_ (
    .CLK(clk_bF$buf54),
    .D(_4331_),
    .Q(\genblk1[5].u_ce.Ain0 [1])
);

DFFPOSX1 _11982_ (
    .CLK(clk_bF$buf53),
    .D(_4332_),
    .Q(\genblk1[5].u_ce.Ycalc [2])
);

DFFPOSX1 _11983_ (
    .CLK(clk_bF$buf52),
    .D(_4333_),
    .Q(\genblk1[5].u_ce.Ycalc [3])
);

DFFPOSX1 _11984_ (
    .CLK(clk_bF$buf51),
    .D(_4334_),
    .Q(\genblk1[5].u_ce.Ycalc [4])
);

DFFPOSX1 _11985_ (
    .CLK(clk_bF$buf50),
    .D(_4335_),
    .Q(\genblk1[5].u_ce.Ycalc [5])
);

DFFPOSX1 _11986_ (
    .CLK(clk_bF$buf49),
    .D(_4336_),
    .Q(\genblk1[5].u_ce.Ycalc [6])
);

DFFPOSX1 _11987_ (
    .CLK(clk_bF$buf48),
    .D(_4337_),
    .Q(\genblk1[5].u_ce.Ycalc [7])
);

DFFPOSX1 _11988_ (
    .CLK(clk_bF$buf47),
    .D(_4338_),
    .Q(\genblk1[5].u_ce.Ycalc [8])
);

DFFPOSX1 _11989_ (
    .CLK(clk_bF$buf46),
    .D(_4339_),
    .Q(\genblk1[5].u_ce.Ycalc [9])
);

DFFPOSX1 _11990_ (
    .CLK(clk_bF$buf45),
    .D(_4340_),
    .Q(\genblk1[5].u_ce.Ycalc [10])
);

DFFPOSX1 _11991_ (
    .CLK(clk_bF$buf44),
    .D(_4341_),
    .Q(\genblk1[5].u_ce.Ycalc [11])
);

DFFPOSX1 _11992_ (
    .CLK(clk_bF$buf43),
    .D(_4342_),
    .Q(\genblk1[5].u_ce.Ycalc [0])
);

DFFPOSX1 _11993_ (
    .CLK(clk_bF$buf42),
    .D(_4343_),
    .Q(\genblk1[5].u_ce.Ycalc [1])
);

DFFPOSX1 _11994_ (
    .CLK(clk_bF$buf41),
    .D(_4344_),
    .Q(\genblk1[5].u_ce.Xcalc [0])
);

DFFPOSX1 _11995_ (
    .CLK(clk_bF$buf40),
    .D(_4345_),
    .Q(\genblk1[5].u_ce.Xcalc [1])
);

DFFPOSX1 _11996_ (
    .CLK(clk_bF$buf39),
    .D(_4346_),
    .Q(\genblk1[5].u_ce.Xcalc [2])
);

DFFPOSX1 _11997_ (
    .CLK(clk_bF$buf38),
    .D(_4347_),
    .Q(\genblk1[5].u_ce.Xcalc [3])
);

DFFPOSX1 _11998_ (
    .CLK(clk_bF$buf37),
    .D(_4348_),
    .Q(\genblk1[5].u_ce.Xcalc [4])
);

DFFPOSX1 _11999_ (
    .CLK(clk_bF$buf36),
    .D(_4349_),
    .Q(\genblk1[5].u_ce.Xcalc [5])
);

DFFPOSX1 _12000_ (
    .CLK(clk_bF$buf35),
    .D(_4350_),
    .Q(\genblk1[5].u_ce.Xcalc [6])
);

DFFPOSX1 _12001_ (
    .CLK(clk_bF$buf34),
    .D(_4351_),
    .Q(\genblk1[5].u_ce.Xcalc [7])
);

DFFPOSX1 _12002_ (
    .CLK(clk_bF$buf33),
    .D(_4352_),
    .Q(\genblk1[5].u_ce.Xcalc [8])
);

DFFPOSX1 _12003_ (
    .CLK(clk_bF$buf32),
    .D(_4353_),
    .Q(\genblk1[5].u_ce.Xcalc [9])
);

DFFPOSX1 _12004_ (
    .CLK(clk_bF$buf31),
    .D(_4354_),
    .Q(\genblk1[5].u_ce.Xcalc [10])
);

DFFPOSX1 _12005_ (
    .CLK(clk_bF$buf30),
    .D(_4355_),
    .Q(\genblk1[5].u_ce.Xcalc [11])
);

DFFPOSX1 _12006_ (
    .CLK(clk_bF$buf29),
    .D(_4356_),
    .Q(\genblk1[5].u_ce.Acalc [1])
);

DFFPOSX1 _12007_ (
    .CLK(clk_bF$buf28),
    .D(_4357_),
    .Q(\genblk1[5].u_ce.Acalc [3])
);

DFFPOSX1 _12008_ (
    .CLK(clk_bF$buf27),
    .D(_4358_),
    .Q(\genblk1[5].u_ce.Acalc [5])
);

DFFPOSX1 _12009_ (
    .CLK(clk_bF$buf26),
    .D(_4359_),
    .Q(\genblk1[5].u_ce.Acalc [7])
);

DFFPOSX1 _12010_ (
    .CLK(clk_bF$buf25),
    .D(_4360_),
    .Q(\genblk1[5].u_ce.Acalc [9])
);

DFFPOSX1 _12011_ (
    .CLK(clk_bF$buf24),
    .D(_4361_),
    .Q(\genblk1[5].u_ce.Acalc [11])
);

DFFPOSX1 _12012_ (
    .CLK(clk_bF$buf23),
    .D(_4362_),
    .Q(\genblk1[5].u_ce.Xin12b [10])
);

DFFPOSX1 _12013_ (
    .CLK(clk_bF$buf22),
    .D(_4363_),
    .Q(\genblk1[5].u_ce.Xin12b [11])
);

DFFPOSX1 _12014_ (
    .CLK(clk_bF$buf21),
    .D(_4364_),
    .Q(\genblk1[5].u_ce.Xin12b [8])
);

DFFPOSX1 _12015_ (
    .CLK(clk_bF$buf20),
    .D(_4365_),
    .Q(\genblk1[5].u_ce.Xin12b [9])
);

DFFPOSX1 _12016_ (
    .CLK(clk_bF$buf19),
    .D(_4366_),
    .Q(\genblk1[5].u_ce.Xin12b [6])
);

DFFPOSX1 _12017_ (
    .CLK(clk_bF$buf18),
    .D(_4367_),
    .Q(\genblk1[5].u_ce.Xin12b [7])
);

DFFPOSX1 _12018_ (
    .CLK(clk_bF$buf17),
    .D(_4368_),
    .Q(\genblk1[5].u_ce.Xin12b [4])
);

DFFPOSX1 _12019_ (
    .CLK(clk_bF$buf16),
    .D(_4369_),
    .Q(\genblk1[5].u_ce.Xin12b [5])
);

DFFPOSX1 _12020_ (
    .CLK(clk_bF$buf15),
    .D(_4370_),
    .Q(\genblk1[5].u_ce.Xin1 [0])
);

DFFPOSX1 _12021_ (
    .CLK(clk_bF$buf14),
    .D(_4371_),
    .Q(\genblk1[5].u_ce.Xin1 [1])
);

DFFPOSX1 _12022_ (
    .CLK(clk_bF$buf13),
    .D(_4372_),
    .Q(\genblk1[5].u_ce.Xin0 [0])
);

DFFPOSX1 _12023_ (
    .CLK(clk_bF$buf12),
    .D(_4373_),
    .Q(\genblk1[5].u_ce.Xin0 [1])
);

DFFPOSX1 _12024_ (
    .CLK(clk_bF$buf11),
    .D(_4374_),
    .Q(\genblk1[5].u_ce.Yin12b [10])
);

DFFPOSX1 _12025_ (
    .CLK(clk_bF$buf10),
    .D(_4375_),
    .Q(\genblk1[5].u_ce.Yin12b [11])
);

DFFPOSX1 _12026_ (
    .CLK(clk_bF$buf9),
    .D(_4376_),
    .Q(\genblk1[5].u_ce.Yin12b [8])
);

DFFPOSX1 _12027_ (
    .CLK(clk_bF$buf8),
    .D(_4377_),
    .Q(\genblk1[5].u_ce.Yin12b [9])
);

DFFPOSX1 _12028_ (
    .CLK(clk_bF$buf7),
    .D(_4378_),
    .Q(\genblk1[5].u_ce.Yin12b [6])
);

DFFPOSX1 _12029_ (
    .CLK(clk_bF$buf6),
    .D(_4379_),
    .Q(\genblk1[5].u_ce.Yin12b [7])
);

DFFPOSX1 _12030_ (
    .CLK(clk_bF$buf5),
    .D(_4380_),
    .Q(\genblk1[5].u_ce.Yin12b [4])
);

DFFPOSX1 _12031_ (
    .CLK(clk_bF$buf4),
    .D(_4381_),
    .Q(\genblk1[5].u_ce.Yin12b [5])
);

DFFPOSX1 _12032_ (
    .CLK(clk_bF$buf3),
    .D(_4382_),
    .Q(\genblk1[5].u_ce.Yin1 [0])
);

DFFPOSX1 _12033_ (
    .CLK(clk_bF$buf2),
    .D(_4383_),
    .Q(\genblk1[5].u_ce.Yin1 [1])
);

DFFPOSX1 _12034_ (
    .CLK(clk_bF$buf1),
    .D(_4384_),
    .Q(\genblk1[5].u_ce.Yin0 [0])
);

DFFPOSX1 _12035_ (
    .CLK(clk_bF$buf0),
    .D(_4385_),
    .Q(\genblk1[5].u_ce.Yin0 [1])
);

DFFPOSX1 _12036_ (
    .CLK(clk_bF$buf75),
    .D(_4386_),
    .Q(\genblk1[5].u_ce.Ain12b [10])
);

DFFPOSX1 _12037_ (
    .CLK(clk_bF$buf74),
    .D(_4387_),
    .Q(\genblk1[5].u_ce.Ain12b [11])
);

DFFPOSX1 _12038_ (
    .CLK(clk_bF$buf73),
    .D(_4388_),
    .Q(\genblk1[5].u_ce.Ain12b [8])
);

DFFPOSX1 _12039_ (
    .CLK(clk_bF$buf72),
    .D(_4389_),
    .Q(\genblk1[5].u_ce.Ain12b [9])
);

DFFPOSX1 _12040_ (
    .CLK(clk_bF$buf71),
    .D(_4390_),
    .Q(\genblk1[5].u_ce.Ain12b [6])
);

DFFPOSX1 _12041_ (
    .CLK(clk_bF$buf70),
    .D(_4391_),
    .Q(\genblk1[5].u_ce.Ain12b [7])
);

DFFPOSX1 _12042_ (
    .CLK(clk_bF$buf69),
    .D(_4392_),
    .Q(\genblk1[5].u_ce.Ain12b [4])
);

DFFPOSX1 _12043_ (
    .CLK(clk_bF$buf68),
    .D(_4393_),
    .Q(\genblk1[5].u_ce.Ain12b [5])
);

DFFPOSX1 _12044_ (
    .CLK(clk_bF$buf67),
    .D(_4394_),
    .Q(\genblk1[5].u_ce.Ain1 [0])
);

DFFPOSX1 _12045_ (
    .CLK(clk_bF$buf66),
    .D(_4395_),
    .Q(\genblk1[5].u_ce.Ain1 [1])
);

DFFPOSX1 _12046_ (
    .CLK(clk_bF$buf65),
    .D(\genblk1[4].u_ce.ISout ),
    .Q(\genblk1[5].u_ce.ISpipe [0])
);

DFFPOSX1 _12047_ (
    .CLK(clk_bF$buf64),
    .D(\genblk1[5].u_ce.ISpipe [0]),
    .Q(\genblk1[5].u_ce.ISpipe [1])
);

DFFPOSX1 _12048_ (
    .CLK(clk_bF$buf63),
    .D(\genblk1[5].u_ce.ISpipe [1]),
    .Q(\genblk1[5].u_ce.ISpipe [2])
);

DFFPOSX1 _12049_ (
    .CLK(clk_bF$buf62),
    .D(\genblk1[5].u_ce.ISpipe [2]),
    .Q(\genblk1[5].u_ce.ISpipe [3])
);

DFFPOSX1 _12050_ (
    .CLK(clk_bF$buf61),
    .D(\genblk1[5].u_ce.ISpipe [3]),
    .Q(\genblk1[5].u_ce.ISpipe [4])
);

DFFPOSX1 _12051_ (
    .CLK(clk_bF$buf60),
    .D(\genblk1[5].u_ce.ISpipe [4]),
    .Q(\genblk1[5].u_ce.ISpipe [5])
);

DFFPOSX1 _12052_ (
    .CLK(clk_bF$buf59),
    .D(\genblk1[5].u_ce.ISpipe [5]),
    .Q(\genblk1[5].u_ce.ISout )
);

DFFPOSX1 _12053_ (
    .CLK(clk_bF$buf58),
    .D(\genblk1[4].u_ce.Vld_bF$buf0 ),
    .Q(\genblk1[5].u_ce.LoadCtl [0])
);

DFFPOSX1 _12054_ (
    .CLK(clk_bF$buf57),
    .D(\genblk1[5].u_ce.LoadCtl_0_bF$buf4 ),
    .Q(\genblk1[5].u_ce.LoadCtl [1])
);

DFFPOSX1 _12055_ (
    .CLK(clk_bF$buf56),
    .D(\genblk1[5].u_ce.LoadCtl [1]),
    .Q(\genblk1[5].u_ce.LoadCtl [2])
);

DFFPOSX1 _12056_ (
    .CLK(clk_bF$buf55),
    .D(\genblk1[5].u_ce.LoadCtl [2]),
    .Q(\genblk1[5].u_ce.LoadCtl [3])
);

DFFPOSX1 _12057_ (
    .CLK(clk_bF$buf54),
    .D(\genblk1[5].u_ce.LoadCtl [3]),
    .Q(\genblk1[5].u_ce.LoadCtl [4])
);

DFFPOSX1 _12058_ (
    .CLK(clk_bF$buf53),
    .D(\genblk1[5].u_ce.LoadCtl [4]),
    .Q(\genblk1[5].u_ce.LoadCtl [5])
);

DFFPOSX1 _12059_ (
    .CLK(clk_bF$buf52),
    .D(\genblk1[5].u_ce.LoadCtl [5]),
    .Q(\genblk1[5].u_ce.Vld )
);

NOR2X1 _12060_ (
    .A(\genblk1[6].u_ce.LoadCtl [3]),
    .B(\genblk1[6].u_ce.LoadCtl [2]),
    .Y(_5224_)
);

INVX2 _12061_ (
    .A(\genblk1[6].u_ce.LoadCtl [2]),
    .Y(_5225_)
);

INVX1 _12062_ (
    .A(\genblk1[6].u_ce.LoadCtl [3]),
    .Y(_5226_)
);

NOR2X1 _12063_ (
    .A(\genblk1[6].u_ce.LoadCtl [2]),
    .B(_5226_),
    .Y(_5227_)
);

NOR2X1 _12064_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[6].u_ce.LoadCtl [1]),
    .Y(_5228_)
);

INVX2 _12065_ (
    .A(_5228_),
    .Y(_5229_)
);

INVX2 _12066_ (
    .A(\genblk1[6].u_ce.LoadCtl [1]),
    .Y(_5230_)
);

NOR2X1 _12067_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_5230_),
    .Y(_5231_)
);

INVX2 _12068_ (
    .A(_5227_),
    .Y(_5232_)
);

INVX1 _12069_ (
    .A(\genblk1[6].u_ce.Ycalc [10]),
    .Y(_5233_)
);

NAND2X1 _12070_ (
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(\genblk1[6].u_ce.Ycalc [8]),
    .Y(_5234_)
);

OAI21X1 _12071_ (
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(_5233_),
    .C(_5234_),
    .Y(_5235_)
);

INVX1 _12072_ (
    .A(\genblk1[6].u_ce.Ycalc [6]),
    .Y(_5236_)
);

INVX1 _12073_ (
    .A(\genblk1[6].u_ce.Ycalc [4]),
    .Y(_5237_)
);

OAI22X1 _12074_ (
    .A(_5225_),
    .B(_5237_),
    .C(_5236_),
    .D(_5232_),
    .Y(_5238_)
);

AOI21X1 _12075_ (
    .A(_5224_),
    .B(_5235_),
    .C(_5238_),
    .Y(_5239_)
);

AOI22X1 _12076_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[6].u_ce.Ycalc [0]),
    .C(_5231_),
    .D(\genblk1[6].u_ce.Ycalc [2]),
    .Y(_5240_)
);

OAI21X1 _12077_ (
    .A(_5229_),
    .B(_5239_),
    .C(_5240_),
    .Y(\genblk1[6].u_ce.Y_ [0])
);

INVX1 _12078_ (
    .A(\genblk1[6].u_ce.Ycalc [11]),
    .Y(_5241_)
);

NAND2X1 _12079_ (
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(\genblk1[6].u_ce.Ycalc [9]),
    .Y(_5242_)
);

OAI21X1 _12080_ (
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(_5241_),
    .C(_5242_),
    .Y(_5243_)
);

INVX1 _12081_ (
    .A(\genblk1[6].u_ce.Ycalc [7]),
    .Y(_5244_)
);

INVX1 _12082_ (
    .A(\genblk1[6].u_ce.Ycalc [5]),
    .Y(_5245_)
);

OAI22X1 _12083_ (
    .A(_5225_),
    .B(_5245_),
    .C(_5244_),
    .D(_5232_),
    .Y(_5246_)
);

AOI21X1 _12084_ (
    .A(_5224_),
    .B(_5243_),
    .C(_5246_),
    .Y(_5247_)
);

AOI22X1 _12085_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[6].u_ce.Ycalc [1]),
    .C(_5231_),
    .D(\genblk1[6].u_ce.Ycalc [3]),
    .Y(_5248_)
);

OAI21X1 _12086_ (
    .A(_5229_),
    .B(_5247_),
    .C(_5248_),
    .Y(\genblk1[6].u_ce.Y_ [1])
);

INVX1 _12087_ (
    .A(\genblk1[6].u_ce.Xcalc [2]),
    .Y(_5249_)
);

INVX2 _12088_ (
    .A(_5231_),
    .Y(_5250_)
);

INVX1 _12089_ (
    .A(\genblk1[6].u_ce.Xcalc [4]),
    .Y(_5251_)
);

INVX1 _12090_ (
    .A(\genblk1[6].u_ce.Xcalc [6]),
    .Y(_5252_)
);

NOR2X1 _12091_ (
    .A(_5226_),
    .B(_5252_),
    .Y(_5253_)
);

INVX1 _12092_ (
    .A(\genblk1[6].u_ce.Xcalc [8]),
    .Y(_5254_)
);

NAND2X1 _12093_ (
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(_5254_),
    .Y(_5255_)
);

OAI21X1 _12094_ (
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(\genblk1[6].u_ce.Xcalc [10]),
    .C(_5255_),
    .Y(_5256_)
);

NOR2X1 _12095_ (
    .A(\genblk1[6].u_ce.LoadCtl [3]),
    .B(_5256_),
    .Y(_5257_)
);

OAI21X1 _12096_ (
    .A(_5253_),
    .B(_5257_),
    .C(_5225_),
    .Y(_5258_)
);

OAI21X1 _12097_ (
    .A(_5225_),
    .B(_5251_),
    .C(_5258_),
    .Y(_5259_)
);

AOI22X1 _12098_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[6].u_ce.Xcalc [0]),
    .C(_5259_),
    .D(_5228_),
    .Y(_5260_)
);

OAI21X1 _12099_ (
    .A(_5249_),
    .B(_5250_),
    .C(_5260_),
    .Y(\genblk1[6].u_ce.X_ [0])
);

INVX1 _12100_ (
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .Y(_5261_)
);

INVX1 _12101_ (
    .A(\genblk1[6].u_ce.Xcalc [9]),
    .Y(_5262_)
);

NAND2X1 _12102_ (
    .A(\genblk1[6].u_ce.Xcalc [11]),
    .B(_5261_),
    .Y(_5263_)
);

OAI21X1 _12103_ (
    .A(_5261_),
    .B(_5262_),
    .C(_5263_),
    .Y(_5264_)
);

INVX1 _12104_ (
    .A(\genblk1[6].u_ce.Xcalc [7]),
    .Y(_5265_)
);

INVX1 _12105_ (
    .A(\genblk1[6].u_ce.Xcalc [5]),
    .Y(_5266_)
);

OAI22X1 _12106_ (
    .A(_5225_),
    .B(_5266_),
    .C(_5265_),
    .D(_5232_),
    .Y(_5267_)
);

AOI21X1 _12107_ (
    .A(_5224_),
    .B(_5264_),
    .C(_5267_),
    .Y(_5268_)
);

AOI22X1 _12108_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[6].u_ce.Xcalc [1]),
    .C(_5231_),
    .D(\genblk1[6].u_ce.Xcalc [3]),
    .Y(_5269_)
);

OAI21X1 _12109_ (
    .A(_5229_),
    .B(_5268_),
    .C(_5269_),
    .Y(\genblk1[6].u_ce.X_ [1])
);

INVX4 _12110_ (
    .A(\genblk1[6].u_ce.Vld ),
    .Y(_5270_)
);

NAND2X1 _12111_ (
    .A(\genblk1[6].u_ce.Ycalc [2]),
    .B(_5270__bF$buf3),
    .Y(_5271_)
);

INVX1 _12112_ (
    .A(1'h0),
    .Y(_5272_)
);

NOR2X1 _12113_ (
    .A(1'h1),
    .B(1'h1),
    .Y(_5273_)
);

NAND2X1 _12114_ (
    .A(_5272_),
    .B(_5273_),
    .Y(_5274_)
);

INVX2 _12115_ (
    .A(_5274_),
    .Y(_5275_)
);

INVX8 _12116_ (
    .A(1'h1),
    .Y(_5276_)
);

MUX2X1 _12117_ (
    .A(\genblk1[6].u_ce.Xin12b [4]),
    .B(\genblk1[6].u_ce.Xin1 [1]),
    .S(1'h0),
    .Y(_5277_)
);

MUX2X1 _12118_ (
    .A(\genblk1[6].u_ce.Xin1 [0]),
    .B(\genblk1[6].u_ce.Xin0 [1]),
    .S(1'h0),
    .Y(_5278_)
);

MUX2X1 _12119_ (
    .A(_5278_),
    .B(_5277_),
    .S(_5276__bF$buf4),
    .Y(_5279_)
);

MUX2X1 _12120_ (
    .A(\genblk1[6].u_ce.Xin12b [8]),
    .B(\genblk1[6].u_ce.Xin12b [7]),
    .S(1'h0),
    .Y(_5280_)
);

MUX2X1 _12121_ (
    .A(\genblk1[6].u_ce.Xin12b [6]),
    .B(\genblk1[6].u_ce.Xin12b [5]),
    .S(1'h0),
    .Y(_5281_)
);

MUX2X1 _12122_ (
    .A(_5281_),
    .B(_5280_),
    .S(_5276__bF$buf3),
    .Y(_5282_)
);

MUX2X1 _12123_ (
    .A(_5282_),
    .B(_5279_),
    .S(1'h1),
    .Y(_5283_)
);

INVX1 _12124_ (
    .A(_5283_),
    .Y(_5284_)
);

MUX2X1 _12125_ (
    .A(\genblk1[6].u_ce.Xin1 [1]),
    .B(\genblk1[6].u_ce.Xin1 [0]),
    .S(1'h0),
    .Y(_5285_)
);

MUX2X1 _12126_ (
    .A(\genblk1[6].u_ce.Xin0 [1]),
    .B(\genblk1[6].u_ce.Xin0 [0]),
    .S(1'h0),
    .Y(_5286_)
);

MUX2X1 _12127_ (
    .A(_5286_),
    .B(_5285_),
    .S(_5276__bF$buf2),
    .Y(_5287_)
);

MUX2X1 _12128_ (
    .A(\genblk1[6].u_ce.Xin12b [7]),
    .B(\genblk1[6].u_ce.Xin12b [6]),
    .S(1'h0),
    .Y(_5288_)
);

MUX2X1 _12129_ (
    .A(\genblk1[6].u_ce.Xin12b [5]),
    .B(\genblk1[6].u_ce.Xin12b [4]),
    .S(1'h0),
    .Y(_5289_)
);

MUX2X1 _12130_ (
    .A(_5289_),
    .B(_5288_),
    .S(_5276__bF$buf1),
    .Y(_5290_)
);

MUX2X1 _12131_ (
    .A(_5290_),
    .B(_5287_),
    .S(1'h1),
    .Y(_5291_)
);

OAI21X1 _12132_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .B(_5291_),
    .C(_5284_),
    .Y(_5292_)
);

NOR2X1 _12133_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5291_),
    .Y(_5293_)
);

NAND2X1 _12134_ (
    .A(_5283_),
    .B(_5293_),
    .Y(_5294_)
);

NAND3X1 _12135_ (
    .A(\genblk1[6].u_ce.Yin0 [1]),
    .B(_5292_),
    .C(_5294_),
    .Y(_5295_)
);

NOR2X1 _12136_ (
    .A(\genblk1[6].u_ce.Yin0 [0]),
    .B(_5291_),
    .Y(_5296_)
);

AOI21X1 _12137_ (
    .A(_5294_),
    .B(_5292_),
    .C(\genblk1[6].u_ce.Yin0 [1]),
    .Y(_5297_)
);

OAI21X1 _12138_ (
    .A(_5296_),
    .B(_5297_),
    .C(_5295_),
    .Y(_5298_)
);

INVX1 _12139_ (
    .A(\genblk1[6].u_ce.Yin1 [0]),
    .Y(_5299_)
);

MUX2X1 _12140_ (
    .A(\genblk1[6].u_ce.Xin12b [9]),
    .B(\genblk1[6].u_ce.Xin12b [8]),
    .S(1'h0),
    .Y(_5300_)
);

MUX2X1 _12141_ (
    .A(_5300_),
    .B(_5288_),
    .S(1'h1),
    .Y(_5301_)
);

AND2X2 _12142_ (
    .A(_5301_),
    .B(1'h1),
    .Y(_5302_)
);

INVX4 _12143_ (
    .A(1'h1),
    .Y(_5303_)
);

NAND2X1 _12144_ (
    .A(_5303__bF$buf3),
    .B(_5276__bF$buf0),
    .Y(_5304_)
);

NAND2X1 _12145_ (
    .A(1'h1),
    .B(_5303__bF$buf2),
    .Y(_5305_)
);

OAI22X1 _12146_ (
    .A(_5304_),
    .B(_5285_),
    .C(_5289_),
    .D(_5305_),
    .Y(_5306_)
);

INVX1 _12147_ (
    .A(\genblk1[6].u_ce.Xin1 [1]),
    .Y(_5307_)
);

NAND2X1 _12148_ (
    .A(_5272_),
    .B(_5307_),
    .Y(_5308_)
);

INVX1 _12149_ (
    .A(\genblk1[6].u_ce.Xin12b [4]),
    .Y(_5309_)
);

NAND2X1 _12150_ (
    .A(1'h0),
    .B(_5309_),
    .Y(_5310_)
);

NAND3X1 _12151_ (
    .A(1'h1),
    .B(_5310_),
    .C(_5308_),
    .Y(_5311_)
);

INVX1 _12152_ (
    .A(\genblk1[6].u_ce.Xin0 [1]),
    .Y(_5312_)
);

NAND2X1 _12153_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Xin1 [0]),
    .Y(_5313_)
);

OAI21X1 _12154_ (
    .A(1'h0),
    .B(_5312_),
    .C(_5313_),
    .Y(_5314_)
);

NAND2X1 _12155_ (
    .A(_5276__bF$buf4),
    .B(_5314_),
    .Y(_5315_)
);

NAND3X1 _12156_ (
    .A(_5303__bF$buf1),
    .B(_5311_),
    .C(_5315_),
    .Y(_5316_)
);

INVX1 _12157_ (
    .A(\genblk1[6].u_ce.Xin12b [5]),
    .Y(_5317_)
);

NAND2X1 _12158_ (
    .A(_5272_),
    .B(_5317_),
    .Y(_5318_)
);

INVX1 _12159_ (
    .A(\genblk1[6].u_ce.Xin12b [6]),
    .Y(_5319_)
);

NAND2X1 _12160_ (
    .A(1'h0),
    .B(_5319_),
    .Y(_5320_)
);

NAND3X1 _12161_ (
    .A(_5276__bF$buf3),
    .B(_5320_),
    .C(_5318_),
    .Y(_5321_)
);

INVX1 _12162_ (
    .A(\genblk1[6].u_ce.Xin12b [7]),
    .Y(_5322_)
);

NAND2X1 _12163_ (
    .A(_5272_),
    .B(_5322_),
    .Y(_5323_)
);

INVX1 _12164_ (
    .A(\genblk1[6].u_ce.Xin12b [8]),
    .Y(_5324_)
);

NAND2X1 _12165_ (
    .A(1'h0),
    .B(_5324_),
    .Y(_5325_)
);

NAND3X1 _12166_ (
    .A(1'h1),
    .B(_5325_),
    .C(_5323_),
    .Y(_5326_)
);

NAND3X1 _12167_ (
    .A(1'h1),
    .B(_5321_),
    .C(_5326_),
    .Y(_5327_)
);

INVX1 _12168_ (
    .A(\genblk1[6].u_ce.Xin1 [0]),
    .Y(_5328_)
);

NAND2X1 _12169_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Xin1 [1]),
    .Y(_5329_)
);

OAI21X1 _12170_ (
    .A(1'h0),
    .B(_5328_),
    .C(_5329_),
    .Y(_5330_)
);

NAND2X1 _12171_ (
    .A(1'h1),
    .B(_5330_),
    .Y(_5331_)
);

INVX1 _12172_ (
    .A(\genblk1[6].u_ce.Xin0 [0]),
    .Y(_5332_)
);

NAND2X1 _12173_ (
    .A(\genblk1[6].u_ce.Xin0 [1]),
    .B(1'h0),
    .Y(_5333_)
);

OAI21X1 _12174_ (
    .A(1'h0),
    .B(_5332_),
    .C(_5333_),
    .Y(_5334_)
);

NAND2X1 _12175_ (
    .A(_5276__bF$buf2),
    .B(_5334_),
    .Y(_5335_)
);

NAND3X1 _12176_ (
    .A(_5303__bF$buf0),
    .B(_5331_),
    .C(_5335_),
    .Y(_5336_)
);

NAND2X1 _12177_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Xin12b [5]),
    .Y(_5337_)
);

OAI21X1 _12178_ (
    .A(1'h0),
    .B(_5309_),
    .C(_5337_),
    .Y(_5338_)
);

NAND2X1 _12179_ (
    .A(_5276__bF$buf1),
    .B(_5338_),
    .Y(_5339_)
);

NAND2X1 _12180_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Xin12b [7]),
    .Y(_5340_)
);

OAI21X1 _12181_ (
    .A(1'h0),
    .B(_5319_),
    .C(_5340_),
    .Y(_5341_)
);

NAND2X1 _12182_ (
    .A(1'h1),
    .B(_5341_),
    .Y(_5342_)
);

NAND3X1 _12183_ (
    .A(1'h1),
    .B(_5339_),
    .C(_5342_),
    .Y(_5343_)
);

AOI22X1 _12184_ (
    .A(_5316_),
    .B(_5327_),
    .C(_5336_),
    .D(_5343_),
    .Y(_5344_)
);

NOR2X1 _12185_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .B(_5344_),
    .Y(_5345_)
);

OAI21X1 _12186_ (
    .A(_5302_),
    .B(_5306_),
    .C(_5345_),
    .Y(_5346_)
);

AOI21X1 _12187_ (
    .A(1'h1),
    .B(_5301_),
    .C(_5306_),
    .Y(_5347_)
);

OAI21X1 _12188_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5344_),
    .C(_5347_),
    .Y(_5348_)
);

NAND3X1 _12189_ (
    .A(_5299_),
    .B(_5348_),
    .C(_5346_),
    .Y(_5349_)
);

NAND2X1 _12190_ (
    .A(_5347_),
    .B(_5345_),
    .Y(_5350_)
);

OAI22X1 _12191_ (
    .A(_5302_),
    .B(_5306_),
    .C(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .D(_5344_),
    .Y(_5351_)
);

NAND3X1 _12192_ (
    .A(\genblk1[6].u_ce.Yin1 [0]),
    .B(_5351_),
    .C(_5350_),
    .Y(_5352_)
);

NAND3X1 _12193_ (
    .A(_5349_),
    .B(_5352_),
    .C(_5298_),
    .Y(_5353_)
);

INVX1 _12194_ (
    .A(\genblk1[6].u_ce.Yin0 [1]),
    .Y(_5354_)
);

NAND2X1 _12195_ (
    .A(_5284_),
    .B(_5293_),
    .Y(_5355_)
);

OAI21X1 _12196_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5291_),
    .C(_5283_),
    .Y(_5356_)
);

AOI21X1 _12197_ (
    .A(_5355_),
    .B(_5356_),
    .C(_5354_),
    .Y(_5357_)
);

INVX1 _12198_ (
    .A(_5296_),
    .Y(_5358_)
);

NAND3X1 _12199_ (
    .A(_5354_),
    .B(_5356_),
    .C(_5355_),
    .Y(_5359_)
);

AOI21X1 _12200_ (
    .A(_5358_),
    .B(_5359_),
    .C(_5357_),
    .Y(_5360_)
);

AOI21X1 _12201_ (
    .A(_5350_),
    .B(_5351_),
    .C(\genblk1[6].u_ce.Yin1 [0]),
    .Y(_5361_)
);

AOI21X1 _12202_ (
    .A(_5346_),
    .B(_5348_),
    .C(_5299_),
    .Y(_5362_)
);

OAI21X1 _12203_ (
    .A(_5361_),
    .B(_5362_),
    .C(_5360_),
    .Y(_5363_)
);

AOI21X1 _12204_ (
    .A(_5353_),
    .B(_5363_),
    .C(_5275_),
    .Y(_5364_)
);

INVX8 _12205_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_5365_)
);

NAND3X1 _12206_ (
    .A(_5303__bF$buf3),
    .B(_5272_),
    .C(_5365__bF$buf5),
    .Y(_5366_)
);

OAI21X1 _12207_ (
    .A(1'h1),
    .B(_5366_),
    .C(\genblk1[6].u_ce.Vld ),
    .Y(_5367_)
);

OAI21X1 _12208_ (
    .A(_5367_),
    .B(_5364_),
    .C(_5271_),
    .Y(_5166_)
);

INVX1 _12209_ (
    .A(\genblk1[6].u_ce.Ycalc [3]),
    .Y(_5368_)
);

INVX1 _12210_ (
    .A(\genblk1[6].u_ce.Xin12b [9]),
    .Y(_5369_)
);

NAND2X1 _12211_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Xin12b [10]),
    .Y(_5370_)
);

OAI21X1 _12212_ (
    .A(1'h0),
    .B(_5369_),
    .C(_5370_),
    .Y(_5371_)
);

NAND2X1 _12213_ (
    .A(1'h1),
    .B(_5371_),
    .Y(_5372_)
);

OAI21X1 _12214_ (
    .A(1'h1),
    .B(_5280_),
    .C(_5372_),
    .Y(_5373_)
);

OAI22X1 _12215_ (
    .A(_5304_),
    .B(_5277_),
    .C(_5281_),
    .D(_5305_),
    .Y(_5374_)
);

AOI21X1 _12216_ (
    .A(_5373_),
    .B(1'h1),
    .C(_5374_),
    .Y(_5375_)
);

NAND3X1 _12217_ (
    .A(_5347_),
    .B(_5283_),
    .C(_5291_),
    .Y(_5376_)
);

INVX1 _12218_ (
    .A(_5376_),
    .Y(_5377_)
);

NOR2X1 _12219_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5377_),
    .Y(_5378_)
);

NAND2X1 _12220_ (
    .A(_5375_),
    .B(_5378_),
    .Y(_5379_)
);

INVX1 _12221_ (
    .A(_5375_),
    .Y(_5380_)
);

OAI21X1 _12222_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .B(_5377_),
    .C(_5380_),
    .Y(_5381_)
);

AOI21X1 _12223_ (
    .A(_5379_),
    .B(_5381_),
    .C(\genblk1[6].u_ce.Yin1 [1]),
    .Y(_5382_)
);

AOI21X1 _12224_ (
    .A(_5298_),
    .B(_5349_),
    .C(_5362_),
    .Y(_5383_)
);

NAND3X1 _12225_ (
    .A(\genblk1[6].u_ce.Yin1 [1]),
    .B(_5381_),
    .C(_5379_),
    .Y(_5384_)
);

NAND2X1 _12226_ (
    .A(_5384_),
    .B(_5383_),
    .Y(_5385_)
);

OAI21X1 _12227_ (
    .A(_5361_),
    .B(_5360_),
    .C(_5352_),
    .Y(_5386_)
);

INVX1 _12228_ (
    .A(\genblk1[6].u_ce.Yin1 [1]),
    .Y(_5387_)
);

NAND2X1 _12229_ (
    .A(_5380_),
    .B(_5378_),
    .Y(_5388_)
);

OAI21X1 _12230_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5377_),
    .C(_5375_),
    .Y(_5389_)
);

AOI21X1 _12231_ (
    .A(_5388_),
    .B(_5389_),
    .C(_5387_),
    .Y(_5390_)
);

OAI21X1 _12232_ (
    .A(_5382_),
    .B(_5390_),
    .C(_5386_),
    .Y(_5391_)
);

OAI21X1 _12233_ (
    .A(_5382_),
    .B(_5385_),
    .C(_5391_),
    .Y(_5392_)
);

OAI21X1 _12234_ (
    .A(_5365__bF$buf4),
    .B(_5274_),
    .C(\genblk1[6].u_ce.Vld ),
    .Y(_5393_)
);

INVX1 _12235_ (
    .A(_5393_),
    .Y(_5394_)
);

OAI21X1 _12236_ (
    .A(_5275_),
    .B(_5392_),
    .C(_5394_),
    .Y(_5395_)
);

OAI21X1 _12237_ (
    .A(_5368_),
    .B(\genblk1[6].u_ce.Vld ),
    .C(_5395_),
    .Y(_5167_)
);

INVX1 _12238_ (
    .A(_5367_),
    .Y(_5396_)
);

INVX1 _12239_ (
    .A(\genblk1[6].u_ce.Yin12b [4]),
    .Y(_5397_)
);

NAND3X1 _12240_ (
    .A(_5347_),
    .B(_5375_),
    .C(_5344_),
    .Y(_5398_)
);

INVX1 _12241_ (
    .A(\genblk1[6].u_ce.Xin12b [10]),
    .Y(_5399_)
);

NAND2X1 _12242_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Xin12b [11]),
    .Y(_5400_)
);

OAI21X1 _12243_ (
    .A(1'h0),
    .B(_5399_),
    .C(_5400_),
    .Y(_5401_)
);

NAND2X1 _12244_ (
    .A(_5276__bF$buf0),
    .B(_5300_),
    .Y(_5402_)
);

OAI21X1 _12245_ (
    .A(_5276__bF$buf4),
    .B(_5401_),
    .C(_5402_),
    .Y(_5403_)
);

NAND2X1 _12246_ (
    .A(_5303__bF$buf2),
    .B(_5290_),
    .Y(_5404_)
);

OAI21X1 _12247_ (
    .A(_5303__bF$buf1),
    .B(_5403_),
    .C(_5404_),
    .Y(_5405_)
);

INVX1 _12248_ (
    .A(_5405_),
    .Y(_5406_)
);

NAND3X1 _12249_ (
    .A(_5365__bF$buf3),
    .B(_5406_),
    .C(_5398_),
    .Y(_5407_)
);

INVX1 _12250_ (
    .A(_5407_),
    .Y(_5408_)
);

AOI21X1 _12251_ (
    .A(_5398_),
    .B(_5365__bF$buf2),
    .C(_5406_),
    .Y(_5409_)
);

OAI21X1 _12252_ (
    .A(_5409_),
    .B(_5408_),
    .C(_5397_),
    .Y(_5410_)
);

OAI21X1 _12253_ (
    .A(_5376_),
    .B(_5380_),
    .C(_5365__bF$buf1),
    .Y(_5411_)
);

NAND2X1 _12254_ (
    .A(_5405_),
    .B(_5411_),
    .Y(_5412_)
);

NAND3X1 _12255_ (
    .A(\genblk1[6].u_ce.Yin12b [4]),
    .B(_5407_),
    .C(_5412_),
    .Y(_5413_)
);

NAND2X1 _12256_ (
    .A(_5413_),
    .B(_5410_),
    .Y(_5414_)
);

INVX1 _12257_ (
    .A(_5382_),
    .Y(_5415_)
);

OAI21X1 _12258_ (
    .A(_5390_),
    .B(_5386_),
    .C(_5415_),
    .Y(_5416_)
);

AOI21X1 _12259_ (
    .A(_5416_),
    .B(_5414_),
    .C(_5275_),
    .Y(_5417_)
);

OAI21X1 _12260_ (
    .A(_5414_),
    .B(_5416_),
    .C(_5417_),
    .Y(_5418_)
);

AOI22X1 _12261_ (
    .A(_5237_),
    .B(_5270__bF$buf2),
    .C(_5418_),
    .D(_5396_),
    .Y(_5168_)
);

INVX1 _12262_ (
    .A(_5413_),
    .Y(_5419_)
);

AOI21X1 _12263_ (
    .A(_5383_),
    .B(_5384_),
    .C(_5382_),
    .Y(_5420_)
);

AOI21X1 _12264_ (
    .A(_5420_),
    .B(_5410_),
    .C(_5419_),
    .Y(_5421_)
);

INVX1 _12265_ (
    .A(\genblk1[6].u_ce.Yin12b [5]),
    .Y(_5422_)
);

NAND3X1 _12266_ (
    .A(_5375_),
    .B(_5406_),
    .C(_5377_),
    .Y(_5423_)
);

INVX1 _12267_ (
    .A(\genblk1[6].u_ce.Xin12b [11]),
    .Y(_5424_)
);

NOR2X1 _12268_ (
    .A(_5276__bF$buf3),
    .B(_5424_),
    .Y(_5425_)
);

AOI21X1 _12269_ (
    .A(_5276__bF$buf2),
    .B(_5371_),
    .C(_5425_),
    .Y(_5426_)
);

NAND2X1 _12270_ (
    .A(_5303__bF$buf0),
    .B(_5282_),
    .Y(_5427_)
);

OAI21X1 _12271_ (
    .A(_5303__bF$buf3),
    .B(_5426_),
    .C(_5427_),
    .Y(_5428_)
);

NAND3X1 _12272_ (
    .A(_5365__bF$buf0),
    .B(_5428_),
    .C(_5423_),
    .Y(_5429_)
);

INVX1 _12273_ (
    .A(_5428_),
    .Y(_5430_)
);

OAI21X1 _12274_ (
    .A(_5405_),
    .B(_5398_),
    .C(_5365__bF$buf5),
    .Y(_5431_)
);

NAND2X1 _12275_ (
    .A(_5430_),
    .B(_5431_),
    .Y(_5432_)
);

NAND3X1 _12276_ (
    .A(_5422_),
    .B(_5432_),
    .C(_5429_),
    .Y(_5433_)
);

NAND3X1 _12277_ (
    .A(_5365__bF$buf4),
    .B(_5430_),
    .C(_5423_),
    .Y(_5434_)
);

NAND2X1 _12278_ (
    .A(_5428_),
    .B(_5431_),
    .Y(_5435_)
);

NAND3X1 _12279_ (
    .A(\genblk1[6].u_ce.Yin12b [5]),
    .B(_5435_),
    .C(_5434_),
    .Y(_5436_)
);

NAND2X1 _12280_ (
    .A(_5433_),
    .B(_5436_),
    .Y(_5437_)
);

INVX1 _12281_ (
    .A(_5437_),
    .Y(_5438_)
);

NOR2X1 _12282_ (
    .A(_5438_),
    .B(_5421_),
    .Y(_5439_)
);

OAI21X1 _12283_ (
    .A(_5414_),
    .B(_5416_),
    .C(_5413_),
    .Y(_5440_)
);

OAI21X1 _12284_ (
    .A(_5437_),
    .B(_5440_),
    .C(_5274_),
    .Y(_5441_)
);

OAI21X1 _12285_ (
    .A(_5441_),
    .B(_5439_),
    .C(_5396_),
    .Y(_5442_)
);

OAI21X1 _12286_ (
    .A(_5245_),
    .B(\genblk1[6].u_ce.Vld ),
    .C(_5442_),
    .Y(_5169_)
);

NOR2X1 _12287_ (
    .A(_5414_),
    .B(_5437_),
    .Y(_5443_)
);

OAI21X1 _12288_ (
    .A(_5413_),
    .B(_5437_),
    .C(_5436_),
    .Y(_5444_)
);

AOI21X1 _12289_ (
    .A(_5443_),
    .B(_5420_),
    .C(_5444_),
    .Y(_5445_)
);

INVX1 _12290_ (
    .A(\genblk1[6].u_ce.Yin12b [6]),
    .Y(_5446_)
);

NOR2X1 _12291_ (
    .A(_5405_),
    .B(_5398_),
    .Y(_5447_)
);

NAND2X1 _12292_ (
    .A(_5430_),
    .B(_5447_),
    .Y(_5448_)
);

AOI21X1 _12293_ (
    .A(_5276__bF$buf1),
    .B(_5401_),
    .C(_5425_),
    .Y(_5449_)
);

NAND2X1 _12294_ (
    .A(_5303__bF$buf2),
    .B(_5301_),
    .Y(_5450_)
);

OAI21X1 _12295_ (
    .A(_5303__bF$buf1),
    .B(_5449_),
    .C(_5450_),
    .Y(_5451_)
);

NAND3X1 _12296_ (
    .A(_5365__bF$buf3),
    .B(_5451_),
    .C(_5448_),
    .Y(_5452_)
);

NOR3X1 _12297_ (
    .A(_5405_),
    .B(_5428_),
    .C(_5398_),
    .Y(_5453_)
);

INVX1 _12298_ (
    .A(_5451_),
    .Y(_5454_)
);

OAI21X1 _12299_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .B(_5453_),
    .C(_5454_),
    .Y(_5455_)
);

NAND3X1 _12300_ (
    .A(_5446_),
    .B(_5455_),
    .C(_5452_),
    .Y(_5456_)
);

NAND3X1 _12301_ (
    .A(_5365__bF$buf2),
    .B(_5454_),
    .C(_5448_),
    .Y(_5457_)
);

OAI21X1 _12302_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5453_),
    .C(_5451_),
    .Y(_5458_)
);

NAND3X1 _12303_ (
    .A(\genblk1[6].u_ce.Yin12b [6]),
    .B(_5458_),
    .C(_5457_),
    .Y(_5459_)
);

AND2X2 _12304_ (
    .A(_5456_),
    .B(_5459_),
    .Y(_5460_)
);

INVX1 _12305_ (
    .A(_5460_),
    .Y(_5461_)
);

AOI21X1 _12306_ (
    .A(_5445_),
    .B(_5461_),
    .C(_5275_),
    .Y(_5462_)
);

OAI21X1 _12307_ (
    .A(_5445_),
    .B(_5461_),
    .C(_5462_),
    .Y(_5463_)
);

AOI22X1 _12308_ (
    .A(_5236_),
    .B(_5270__bF$buf1),
    .C(_5463_),
    .D(_5396_),
    .Y(_5170_)
);

AND2X2 _12309_ (
    .A(_5410_),
    .B(_5413_),
    .Y(_5464_)
);

NAND3X1 _12310_ (
    .A(_5433_),
    .B(_5436_),
    .C(_5464_),
    .Y(_5465_)
);

INVX1 _12311_ (
    .A(_5436_),
    .Y(_5466_)
);

AOI21X1 _12312_ (
    .A(_5419_),
    .B(_5433_),
    .C(_5466_),
    .Y(_5467_)
);

OAI21X1 _12313_ (
    .A(_5416_),
    .B(_5465_),
    .C(_5467_),
    .Y(_5468_)
);

INVX1 _12314_ (
    .A(_5459_),
    .Y(_5469_)
);

AOI21X1 _12315_ (
    .A(_5468_),
    .B(_5456_),
    .C(_5469_),
    .Y(_5470_)
);

INVX1 _12316_ (
    .A(\genblk1[6].u_ce.Yin12b [7]),
    .Y(_5471_)
);

NAND2X1 _12317_ (
    .A(_5454_),
    .B(_5453_),
    .Y(_5472_)
);

NOR2X1 _12318_ (
    .A(_5303__bF$buf0),
    .B(_5424_),
    .Y(_5473_)
);

AOI21X1 _12319_ (
    .A(_5373_),
    .B(_5303__bF$buf3),
    .C(_5473_),
    .Y(_5474_)
);

INVX1 _12320_ (
    .A(_5474_),
    .Y(_5475_)
);

NAND3X1 _12321_ (
    .A(_5365__bF$buf1),
    .B(_5475_),
    .C(_5472_),
    .Y(_5476_)
);

AND2X2 _12322_ (
    .A(_5453_),
    .B(_5454_),
    .Y(_5477_)
);

OAI21X1 _12323_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .B(_5477_),
    .C(_5474_),
    .Y(_5478_)
);

NAND3X1 _12324_ (
    .A(_5471_),
    .B(_5476_),
    .C(_5478_),
    .Y(_5479_)
);

NAND3X1 _12325_ (
    .A(_5365__bF$buf0),
    .B(_5474_),
    .C(_5472_),
    .Y(_5480_)
);

OAI21X1 _12326_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5477_),
    .C(_5475_),
    .Y(_5481_)
);

NAND3X1 _12327_ (
    .A(\genblk1[6].u_ce.Yin12b [7]),
    .B(_5480_),
    .C(_5481_),
    .Y(_5482_)
);

AND2X2 _12328_ (
    .A(_5479_),
    .B(_5482_),
    .Y(_5483_)
);

NOR2X1 _12329_ (
    .A(_5483_),
    .B(_5470_),
    .Y(_5484_)
);

NAND2X1 _12330_ (
    .A(_5272_),
    .B(_5276__bF$buf0),
    .Y(_5485_)
);

NAND2X1 _12331_ (
    .A(_5483_),
    .B(_5470_),
    .Y(_5486_)
);

OAI21X1 _12332_ (
    .A(1'h1),
    .B(_5485_),
    .C(_5486_),
    .Y(_5487_)
);

OAI21X1 _12333_ (
    .A(_5484_),
    .B(_5487_),
    .C(_5394_),
    .Y(_5488_)
);

OAI21X1 _12334_ (
    .A(_5244_),
    .B(\genblk1[6].u_ce.Vld ),
    .C(_5488_),
    .Y(_5171_)
);

INVX1 _12335_ (
    .A(\genblk1[6].u_ce.Ycalc [8]),
    .Y(_5489_)
);

AOI21X1 _12336_ (
    .A(_5478_),
    .B(_5476_),
    .C(_5471_),
    .Y(_5490_)
);

OAI21X1 _12337_ (
    .A(_5469_),
    .B(_5490_),
    .C(_5479_),
    .Y(_5491_)
);

NAND3X1 _12338_ (
    .A(_5460_),
    .B(_5483_),
    .C(_5468_),
    .Y(_5492_)
);

INVX1 _12339_ (
    .A(\genblk1[6].u_ce.Yin12b [8]),
    .Y(_5493_)
);

NAND3X1 _12340_ (
    .A(_5454_),
    .B(_5474_),
    .C(_5453_),
    .Y(_5494_)
);

INVX1 _12341_ (
    .A(_5473_),
    .Y(_5495_)
);

OAI21X1 _12342_ (
    .A(1'h1),
    .B(_5403_),
    .C(_5495_),
    .Y(_5496_)
);

NAND3X1 _12343_ (
    .A(_5365__bF$buf5),
    .B(_5496_),
    .C(_5494_),
    .Y(_5497_)
);

INVX1 _12344_ (
    .A(_5496_),
    .Y(_5498_)
);

NAND2X1 _12345_ (
    .A(_5365__bF$buf4),
    .B(_5494_),
    .Y(_5499_)
);

NAND2X1 _12346_ (
    .A(_5498_),
    .B(_5499_),
    .Y(_5500_)
);

NAND3X1 _12347_ (
    .A(_5493_),
    .B(_5497_),
    .C(_5500_),
    .Y(_5501_)
);

NAND3X1 _12348_ (
    .A(_5365__bF$buf3),
    .B(_5498_),
    .C(_5494_),
    .Y(_5502_)
);

NAND2X1 _12349_ (
    .A(_5496_),
    .B(_5499_),
    .Y(_5503_)
);

NAND3X1 _12350_ (
    .A(\genblk1[6].u_ce.Yin12b [8]),
    .B(_5502_),
    .C(_5503_),
    .Y(_5504_)
);

AND2X2 _12351_ (
    .A(_5501_),
    .B(_5504_),
    .Y(_5505_)
);

INVX1 _12352_ (
    .A(_5505_),
    .Y(_5506_)
);

AOI21X1 _12353_ (
    .A(_5492_),
    .B(_5491_),
    .C(_5506_),
    .Y(_5507_)
);

NAND3X1 _12354_ (
    .A(_5479_),
    .B(_5482_),
    .C(_5460_),
    .Y(_5508_)
);

OAI21X1 _12355_ (
    .A(_5508_),
    .B(_5445_),
    .C(_5491_),
    .Y(_5509_)
);

OAI21X1 _12356_ (
    .A(_5505_),
    .B(_5509_),
    .C(_5274_),
    .Y(_5510_)
);

OR2X2 _12357_ (
    .A(_5510_),
    .B(_5507_),
    .Y(_5511_)
);

AOI22X1 _12358_ (
    .A(_5489_),
    .B(_5270__bF$buf0),
    .C(_5511_),
    .D(_5394_),
    .Y(_5172_)
);

INVX1 _12359_ (
    .A(\genblk1[6].u_ce.Ycalc [9]),
    .Y(_5512_)
);

INVX1 _12360_ (
    .A(_5504_),
    .Y(_5513_)
);

NOR2X1 _12361_ (
    .A(_5513_),
    .B(_5507_),
    .Y(_5514_)
);

INVX1 _12362_ (
    .A(\genblk1[6].u_ce.Yin12b [9]),
    .Y(_5515_)
);

OAI21X1 _12363_ (
    .A(1'h1),
    .B(_5426_),
    .C(_5495_),
    .Y(_5516_)
);

INVX1 _12364_ (
    .A(_5516_),
    .Y(_5517_)
);

OAI21X1 _12365_ (
    .A(_5496_),
    .B(_5494_),
    .C(_5365__bF$buf2),
    .Y(_5518_)
);

NAND2X1 _12366_ (
    .A(_5517_),
    .B(_5518_),
    .Y(_5519_)
);

NAND3X1 _12367_ (
    .A(_5474_),
    .B(_5498_),
    .C(_5477_),
    .Y(_5520_)
);

NAND3X1 _12368_ (
    .A(_5365__bF$buf1),
    .B(_5516_),
    .C(_5520_),
    .Y(_5521_)
);

NAND3X1 _12369_ (
    .A(_5515_),
    .B(_5519_),
    .C(_5521_),
    .Y(_5522_)
);

AND2X2 _12370_ (
    .A(_5518_),
    .B(_5517_),
    .Y(_5523_)
);

NOR2X1 _12371_ (
    .A(_5517_),
    .B(_5518_),
    .Y(_5524_)
);

OAI21X1 _12372_ (
    .A(_5524_),
    .B(_5523_),
    .C(\genblk1[6].u_ce.Yin12b [9]),
    .Y(_5525_)
);

NAND2X1 _12373_ (
    .A(_5522_),
    .B(_5525_),
    .Y(_5526_)
);

AOI21X1 _12374_ (
    .A(_5514_),
    .B(_5526_),
    .C(_5275_),
    .Y(_5527_)
);

OAI21X1 _12375_ (
    .A(_5514_),
    .B(_5526_),
    .C(_5527_),
    .Y(_5528_)
);

AOI22X1 _12376_ (
    .A(_5512_),
    .B(_5270__bF$buf3),
    .C(_5528_),
    .D(_5394_),
    .Y(_5173_)
);

OAI21X1 _12377_ (
    .A(_5504_),
    .B(_5526_),
    .C(_5525_),
    .Y(_5529_)
);

NAND3X1 _12378_ (
    .A(_5522_),
    .B(_5525_),
    .C(_5505_),
    .Y(_5530_)
);

AOI21X1 _12379_ (
    .A(_5491_),
    .B(_5492_),
    .C(_5530_),
    .Y(_5531_)
);

INVX1 _12380_ (
    .A(\genblk1[6].u_ce.Yin12b [10]),
    .Y(_5532_)
);

OAI21X1 _12381_ (
    .A(1'h1),
    .B(_5449_),
    .C(_5495_),
    .Y(_5533_)
);

INVX1 _12382_ (
    .A(_5533_),
    .Y(_5534_)
);

OAI21X1 _12383_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .B(_5517_),
    .C(_5518_),
    .Y(_5535_)
);

NAND2X1 _12384_ (
    .A(_5534_),
    .B(_5535_),
    .Y(_5536_)
);

OAI21X1 _12385_ (
    .A(_5516_),
    .B(_5520_),
    .C(_5365__bF$buf0),
    .Y(_5537_)
);

NAND2X1 _12386_ (
    .A(_5533_),
    .B(_5537_),
    .Y(_5538_)
);

NAND2X1 _12387_ (
    .A(_5536_),
    .B(_5538_),
    .Y(_5539_)
);

NAND2X1 _12388_ (
    .A(_5532_),
    .B(_5539_),
    .Y(_5540_)
);

NAND3X1 _12389_ (
    .A(\genblk1[6].u_ce.Yin12b [10]),
    .B(_5536_),
    .C(_5538_),
    .Y(_5541_)
);

AND2X2 _12390_ (
    .A(_5540_),
    .B(_5541_),
    .Y(_5542_)
);

OAI21X1 _12391_ (
    .A(_5529_),
    .B(_5531_),
    .C(_5542_),
    .Y(_5543_)
);

INVX1 _12392_ (
    .A(_5525_),
    .Y(_5544_)
);

AOI21X1 _12393_ (
    .A(_5513_),
    .B(_5522_),
    .C(_5544_),
    .Y(_5545_)
);

AND2X2 _12394_ (
    .A(_5525_),
    .B(_5522_),
    .Y(_5546_)
);

NAND3X1 _12395_ (
    .A(_5505_),
    .B(_5546_),
    .C(_5509_),
    .Y(_5547_)
);

NAND2X1 _12396_ (
    .A(_5541_),
    .B(_5540_),
    .Y(_5548_)
);

NAND3X1 _12397_ (
    .A(_5545_),
    .B(_5548_),
    .C(_5547_),
    .Y(_5549_)
);

NAND3X1 _12398_ (
    .A(_5274_),
    .B(_5549_),
    .C(_5543_),
    .Y(_5550_)
);

AOI22X1 _12399_ (
    .A(_5233_),
    .B(_5270__bF$buf2),
    .C(_5550_),
    .D(_5396_),
    .Y(_5174_)
);

INVX1 _12400_ (
    .A(_5541_),
    .Y(_5551_)
);

AOI21X1 _12401_ (
    .A(_5547_),
    .B(_5545_),
    .C(_5548_),
    .Y(_5552_)
);

OAI21X1 _12402_ (
    .A(_5533_),
    .B(_5535_),
    .C(_5365__bF$buf5),
    .Y(_5553_)
);

INVX1 _12403_ (
    .A(_5553_),
    .Y(_5554_)
);

NAND2X1 _12404_ (
    .A(\genblk1[6].u_ce.Yin12b [11]),
    .B(_5424_),
    .Y(_5555_)
);

INVX1 _12405_ (
    .A(\genblk1[6].u_ce.Yin12b [11]),
    .Y(_5556_)
);

NAND2X1 _12406_ (
    .A(\genblk1[6].u_ce.Xin12b [11]),
    .B(_5556_),
    .Y(_5557_)
);

NAND2X1 _12407_ (
    .A(_5555_),
    .B(_5557_),
    .Y(_5558_)
);

OR2X2 _12408_ (
    .A(_5554_),
    .B(_5558_),
    .Y(_5559_)
);

NAND2X1 _12409_ (
    .A(_5558_),
    .B(_5554_),
    .Y(_5560_)
);

NAND2X1 _12410_ (
    .A(_5560_),
    .B(_5559_),
    .Y(_5561_)
);

OAI21X1 _12411_ (
    .A(_5551_),
    .B(_5552_),
    .C(_5561_),
    .Y(_5562_)
);

INVX1 _12412_ (
    .A(_5561_),
    .Y(_5563_)
);

NAND3X1 _12413_ (
    .A(_5541_),
    .B(_5563_),
    .C(_5543_),
    .Y(_5564_)
);

NAND3X1 _12414_ (
    .A(_5274_),
    .B(_5564_),
    .C(_5562_),
    .Y(_5565_)
);

AOI22X1 _12415_ (
    .A(_5241_),
    .B(_5270__bF$buf1),
    .C(_5565_),
    .D(_5394_),
    .Y(_5175_)
);

INVX1 _12416_ (
    .A(\genblk1[6].u_ce.Ycalc [0]),
    .Y(_5566_)
);

OAI21X1 _12417_ (
    .A(1'h1),
    .B(_5485_),
    .C(\genblk1[6].u_ce.Vld ),
    .Y(_5567_)
);

INVX2 _12418_ (
    .A(_5567_),
    .Y(_5568_)
);

INVX1 _12419_ (
    .A(\genblk1[6].u_ce.Yin0 [0]),
    .Y(_5569_)
);

AOI21X1 _12420_ (
    .A(_5336_),
    .B(_5343_),
    .C(_5569_),
    .Y(_5570_)
);

OAI21X1 _12421_ (
    .A(_5570_),
    .B(_5296_),
    .C(_5568_),
    .Y(_5571_)
);

OAI21X1 _12422_ (
    .A(_5566_),
    .B(\genblk1[6].u_ce.Vld ),
    .C(_5571_),
    .Y(_5176_)
);

NAND2X1 _12423_ (
    .A(\genblk1[6].u_ce.Ycalc [1]),
    .B(_5270__bF$buf0),
    .Y(_5572_)
);

NAND3X1 _12424_ (
    .A(_5358_),
    .B(_5295_),
    .C(_5359_),
    .Y(_5573_)
);

OAI21X1 _12425_ (
    .A(_5357_),
    .B(_5297_),
    .C(_5296_),
    .Y(_5574_)
);

AOI21X1 _12426_ (
    .A(_5574_),
    .B(_5573_),
    .C(_5275_),
    .Y(_5575_)
);

OAI21X1 _12427_ (
    .A(_5270__bF$buf3),
    .B(_5575_),
    .C(_5572_),
    .Y(_5177_)
);

NAND2X1 _12428_ (
    .A(\genblk1[6].u_ce.Xcalc [0]),
    .B(_5270__bF$buf2),
    .Y(_5576_)
);

MUX2X1 _12429_ (
    .A(\genblk1[6].u_ce.Yin12b [7]),
    .B(\genblk1[6].u_ce.Yin12b [6]),
    .S(1'h0),
    .Y(_5577_)
);

NAND2X1 _12430_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin12b [5]),
    .Y(_5578_)
);

OAI21X1 _12431_ (
    .A(1'h0),
    .B(_5397_),
    .C(_5578_),
    .Y(_5579_)
);

NAND2X1 _12432_ (
    .A(_5276__bF$buf4),
    .B(_5579_),
    .Y(_5580_)
);

OAI21X1 _12433_ (
    .A(_5276__bF$buf3),
    .B(_5577_),
    .C(_5580_),
    .Y(_5581_)
);

NAND2X1 _12434_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin1 [1]),
    .Y(_5582_)
);

OAI21X1 _12435_ (
    .A(1'h0),
    .B(_5299_),
    .C(_5582_),
    .Y(_5583_)
);

NAND2X1 _12436_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin0 [1]),
    .Y(_5584_)
);

OAI21X1 _12437_ (
    .A(1'h0),
    .B(_5569_),
    .C(_5584_),
    .Y(_5585_)
);

MUX2X1 _12438_ (
    .A(_5585_),
    .B(_5583_),
    .S(_5276__bF$buf2),
    .Y(_5586_)
);

NAND2X1 _12439_ (
    .A(_5303__bF$buf2),
    .B(_5586_),
    .Y(_5587_)
);

OAI21X1 _12440_ (
    .A(_5303__bF$buf1),
    .B(_5581_),
    .C(_5587_),
    .Y(_5588_)
);

INVX1 _12441_ (
    .A(_5588_),
    .Y(_5589_)
);

NOR2X1 _12442_ (
    .A(\genblk1[6].u_ce.Xin0 [0]),
    .B(_5589_),
    .Y(_5590_)
);

OAI21X1 _12443_ (
    .A(_5332_),
    .B(_5588_),
    .C(_5568_),
    .Y(_5591_)
);

OAI21X1 _12444_ (
    .A(_5591_),
    .B(_5590_),
    .C(_5576_),
    .Y(_5178_)
);

NAND2X1 _12445_ (
    .A(\genblk1[6].u_ce.Xcalc [1]),
    .B(_5270__bF$buf1),
    .Y(_5592_)
);

NOR2X1 _12446_ (
    .A(_5332_),
    .B(_5588_),
    .Y(_5593_)
);

NAND2X1 _12447_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin12b [4]),
    .Y(_5594_)
);

OAI21X1 _12448_ (
    .A(1'h0),
    .B(_5387_),
    .C(_5594_),
    .Y(_5595_)
);

NAND2X1 _12449_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin1 [0]),
    .Y(_5596_)
);

OAI21X1 _12450_ (
    .A(1'h0),
    .B(_5354_),
    .C(_5596_),
    .Y(_5597_)
);

MUX2X1 _12451_ (
    .A(_5597_),
    .B(_5595_),
    .S(_5276__bF$buf1),
    .Y(_5598_)
);

NAND2X1 _12452_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin12b [8]),
    .Y(_5599_)
);

OAI21X1 _12453_ (
    .A(1'h0),
    .B(_5471_),
    .C(_5599_),
    .Y(_5600_)
);

NAND2X1 _12454_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin12b [6]),
    .Y(_5601_)
);

OAI21X1 _12455_ (
    .A(1'h0),
    .B(_5422_),
    .C(_5601_),
    .Y(_5602_)
);

MUX2X1 _12456_ (
    .A(_5602_),
    .B(_5600_),
    .S(_5276__bF$buf0),
    .Y(_5603_)
);

MUX2X1 _12457_ (
    .A(_5603_),
    .B(_5598_),
    .S(1'h1),
    .Y(_5604_)
);

NOR2X1 _12458_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5588_),
    .Y(_5605_)
);

NAND2X1 _12459_ (
    .A(_5604_),
    .B(_5605_),
    .Y(_5606_)
);

NAND2X1 _12460_ (
    .A(_5303__bF$buf0),
    .B(_5598_),
    .Y(_5607_)
);

NAND2X1 _12461_ (
    .A(1'h1),
    .B(_5603_),
    .Y(_5608_)
);

NAND2X1 _12462_ (
    .A(_5607_),
    .B(_5608_),
    .Y(_5609_)
);

OAI21X1 _12463_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .B(_5588_),
    .C(_5609_),
    .Y(_5610_)
);

NAND3X1 _12464_ (
    .A(\genblk1[6].u_ce.Xin0 [1]),
    .B(_5610_),
    .C(_5606_),
    .Y(_5611_)
);

OAI21X1 _12465_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5588_),
    .C(_5604_),
    .Y(_5612_)
);

NAND2X1 _12466_ (
    .A(_5609_),
    .B(_5605_),
    .Y(_5613_)
);

NAND3X1 _12467_ (
    .A(_5312_),
    .B(_5612_),
    .C(_5613_),
    .Y(_5614_)
);

NAND3X1 _12468_ (
    .A(_5593_),
    .B(_5611_),
    .C(_5614_),
    .Y(_5615_)
);

INVX1 _12469_ (
    .A(_5593_),
    .Y(_5616_)
);

AOI21X1 _12470_ (
    .A(_5613_),
    .B(_5612_),
    .C(_5312_),
    .Y(_5617_)
);

AOI21X1 _12471_ (
    .A(_5606_),
    .B(_5610_),
    .C(\genblk1[6].u_ce.Xin0 [1]),
    .Y(_5618_)
);

OAI21X1 _12472_ (
    .A(_5617_),
    .B(_5618_),
    .C(_5616_),
    .Y(_5619_)
);

AOI21X1 _12473_ (
    .A(_5619_),
    .B(_5615_),
    .C(_5275_),
    .Y(_5620_)
);

OAI21X1 _12474_ (
    .A(_5270__bF$buf0),
    .B(_5620_),
    .C(_5592_),
    .Y(_5179_)
);

OAI21X1 _12475_ (
    .A(_5616_),
    .B(_5618_),
    .C(_5611_),
    .Y(_5621_)
);

MUX2X1 _12476_ (
    .A(\genblk1[6].u_ce.Yin12b [9]),
    .B(\genblk1[6].u_ce.Yin12b [8]),
    .S(1'h0),
    .Y(_5622_)
);

MUX2X1 _12477_ (
    .A(_5622_),
    .B(_5577_),
    .S(1'h1),
    .Y(_5623_)
);

NOR2X1 _12478_ (
    .A(1'h1),
    .B(_5276__bF$buf4),
    .Y(_5624_)
);

NAND2X1 _12479_ (
    .A(_5579_),
    .B(_5624_),
    .Y(_5625_)
);

NAND2X1 _12480_ (
    .A(_5273_),
    .B(_5583_),
    .Y(_5626_)
);

NAND2X1 _12481_ (
    .A(_5626_),
    .B(_5625_),
    .Y(_5627_)
);

AOI21X1 _12482_ (
    .A(1'h1),
    .B(_5623_),
    .C(_5627_),
    .Y(_5628_)
);

NAND2X1 _12483_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin12b [7]),
    .Y(_5629_)
);

OAI21X1 _12484_ (
    .A(1'h0),
    .B(_5446_),
    .C(_5629_),
    .Y(_5630_)
);

MUX2X1 _12485_ (
    .A(_5579_),
    .B(_5630_),
    .S(_5276__bF$buf3),
    .Y(_5631_)
);

NAND2X1 _12486_ (
    .A(1'h1),
    .B(_5631_),
    .Y(_5632_)
);

AOI21X1 _12487_ (
    .A(_5587_),
    .B(_5632_),
    .C(_5604_),
    .Y(_5633_)
);

NOR2X1 _12488_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .B(_5633_),
    .Y(_5634_)
);

NAND2X1 _12489_ (
    .A(_5628_),
    .B(_5634_),
    .Y(_5635_)
);

INVX1 _12490_ (
    .A(_5628_),
    .Y(_5636_)
);

OAI21X1 _12491_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5633_),
    .C(_5636_),
    .Y(_5637_)
);

AOI21X1 _12492_ (
    .A(_5635_),
    .B(_5637_),
    .C(_5328_),
    .Y(_5638_)
);

NAND3X1 _12493_ (
    .A(_5328_),
    .B(_5637_),
    .C(_5635_),
    .Y(_5639_)
);

INVX1 _12494_ (
    .A(_5639_),
    .Y(_5640_)
);

NOR2X1 _12495_ (
    .A(_5638_),
    .B(_5640_),
    .Y(_5641_)
);

NOR2X1 _12496_ (
    .A(_5621_),
    .B(_5641_),
    .Y(_5642_)
);

AOI21X1 _12497_ (
    .A(_5593_),
    .B(_5614_),
    .C(_5617_),
    .Y(_5643_)
);

INVX1 _12498_ (
    .A(_5641_),
    .Y(_5644_)
);

OAI21X1 _12499_ (
    .A(_5643_),
    .B(_5644_),
    .C(_5568_),
    .Y(_5645_)
);

OAI22X1 _12500_ (
    .A(_5249_),
    .B(\genblk1[6].u_ce.Vld ),
    .C(_5642_),
    .D(_5645_),
    .Y(_5180_)
);

NAND2X1 _12501_ (
    .A(\genblk1[6].u_ce.Xcalc [3]),
    .B(_5270__bF$buf3),
    .Y(_5646_)
);

AOI21X1 _12502_ (
    .A(_5621_),
    .B(_5639_),
    .C(_5638_),
    .Y(_5647_)
);

NAND2X1 _12503_ (
    .A(1'h0),
    .B(_5532_),
    .Y(_5648_)
);

OAI21X1 _12504_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin12b [9]),
    .C(_5648_),
    .Y(_5649_)
);

NAND2X1 _12505_ (
    .A(_5276__bF$buf2),
    .B(_5600_),
    .Y(_5650_)
);

OAI21X1 _12506_ (
    .A(_5276__bF$buf1),
    .B(_5649_),
    .C(_5650_),
    .Y(_5651_)
);

NAND2X1 _12507_ (
    .A(_5602_),
    .B(_5624_),
    .Y(_5652_)
);

NAND2X1 _12508_ (
    .A(_5273_),
    .B(_5595_),
    .Y(_5653_)
);

NAND2X1 _12509_ (
    .A(_5653_),
    .B(_5652_),
    .Y(_5654_)
);

AOI21X1 _12510_ (
    .A(_5651_),
    .B(1'h1),
    .C(_5654_),
    .Y(_5655_)
);

NAND3X1 _12511_ (
    .A(_5628_),
    .B(_5609_),
    .C(_5588_),
    .Y(_5656_)
);

NAND2X1 _12512_ (
    .A(_5365__bF$buf4),
    .B(_5656_),
    .Y(_5657_)
);

OR2X2 _12513_ (
    .A(_5657_),
    .B(_5655_),
    .Y(_5658_)
);

INVX1 _12514_ (
    .A(_5656_),
    .Y(_5659_)
);

OAI21X1 _12515_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf3 ),
    .B(_5659_),
    .C(_5655_),
    .Y(_5660_)
);

NAND3X1 _12516_ (
    .A(\genblk1[6].u_ce.Xin1 [1]),
    .B(_5660_),
    .C(_5658_),
    .Y(_5661_)
);

INVX1 _12517_ (
    .A(_5655_),
    .Y(_5662_)
);

OR2X2 _12518_ (
    .A(_5657_),
    .B(_5662_),
    .Y(_5663_)
);

OAI21X1 _12519_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf2 ),
    .B(_5659_),
    .C(_5662_),
    .Y(_5664_)
);

NAND3X1 _12520_ (
    .A(_5307_),
    .B(_5664_),
    .C(_5663_),
    .Y(_5665_)
);

NAND2X1 _12521_ (
    .A(_5661_),
    .B(_5665_),
    .Y(_5666_)
);

OR2X2 _12522_ (
    .A(_5647_),
    .B(_5666_),
    .Y(_5667_)
);

NAND2X1 _12523_ (
    .A(_5666_),
    .B(_5647_),
    .Y(_5668_)
);

AOI21X1 _12524_ (
    .A(_5667_),
    .B(_5668_),
    .C(_5275_),
    .Y(_5669_)
);

OAI21X1 _12525_ (
    .A(_5270__bF$buf2),
    .B(_5669_),
    .C(_5646_),
    .Y(_5181_)
);

OAI21X1 _12526_ (
    .A(_5666_),
    .B(_5647_),
    .C(_5661_),
    .Y(_5670_)
);

NAND2X1 _12527_ (
    .A(1'h0),
    .B(\genblk1[6].u_ce.Yin12b [11]),
    .Y(_5671_)
);

OAI21X1 _12528_ (
    .A(1'h0),
    .B(_5532_),
    .C(_5671_),
    .Y(_5672_)
);

NAND2X1 _12529_ (
    .A(1'h1),
    .B(_5672_),
    .Y(_5673_)
);

OAI21X1 _12530_ (
    .A(1'h1),
    .B(_5622_),
    .C(_5673_),
    .Y(_5674_)
);

NAND2X1 _12531_ (
    .A(1'h1),
    .B(_5674_),
    .Y(_5675_)
);

OAI21X1 _12532_ (
    .A(1'h1),
    .B(_5631_),
    .C(_5675_),
    .Y(_5676_)
);

INVX1 _12533_ (
    .A(_5676_),
    .Y(_5677_)
);

OAI21X1 _12534_ (
    .A(_5662_),
    .B(_5656_),
    .C(_5365__bF$buf3),
    .Y(_5678_)
);

OR2X2 _12535_ (
    .A(_5678_),
    .B(_5677_),
    .Y(_5679_)
);

NAND2X1 _12536_ (
    .A(_5677_),
    .B(_5678_),
    .Y(_5680_)
);

NAND3X1 _12537_ (
    .A(\genblk1[6].u_ce.Xin12b [4]),
    .B(_5680_),
    .C(_5679_),
    .Y(_5681_)
);

OR2X2 _12538_ (
    .A(_5678_),
    .B(_5676_),
    .Y(_5682_)
);

NAND2X1 _12539_ (
    .A(_5676_),
    .B(_5678_),
    .Y(_5683_)
);

NAND3X1 _12540_ (
    .A(_5309_),
    .B(_5683_),
    .C(_5682_),
    .Y(_5684_)
);

AND2X2 _12541_ (
    .A(_5681_),
    .B(_5684_),
    .Y(_5685_)
);

NAND2X1 _12542_ (
    .A(_5685_),
    .B(_5670_),
    .Y(_5686_)
);

INVX1 _12543_ (
    .A(_5638_),
    .Y(_5687_)
);

OAI21X1 _12544_ (
    .A(_5640_),
    .B(_5643_),
    .C(_5687_),
    .Y(_5688_)
);

INVX1 _12545_ (
    .A(_5661_),
    .Y(_5689_)
);

AOI21X1 _12546_ (
    .A(_5688_),
    .B(_5665_),
    .C(_5689_),
    .Y(_5690_)
);

NAND2X1 _12547_ (
    .A(_5684_),
    .B(_5681_),
    .Y(_5691_)
);

NAND2X1 _12548_ (
    .A(_5691_),
    .B(_5690_),
    .Y(_5692_)
);

NAND2X1 _12549_ (
    .A(_5686_),
    .B(_5692_),
    .Y(_5693_)
);

AOI22X1 _12550_ (
    .A(_5251_),
    .B(_5270__bF$buf1),
    .C(_5693_),
    .D(_5568_),
    .Y(_5182_)
);

NAND3X1 _12551_ (
    .A(_5655_),
    .B(_5677_),
    .C(_5659_),
    .Y(_5694_)
);

NOR2X1 _12552_ (
    .A(1'h1),
    .B(_5649_),
    .Y(_5695_)
);

NOR2X1 _12553_ (
    .A(_5276__bF$buf0),
    .B(_5556_),
    .Y(_5696_)
);

OAI21X1 _12554_ (
    .A(_5696_),
    .B(_5695_),
    .C(1'h1),
    .Y(_5697_)
);

OAI21X1 _12555_ (
    .A(1'h1),
    .B(_5603_),
    .C(_5697_),
    .Y(_5698_)
);

NAND3X1 _12556_ (
    .A(_5365__bF$buf2),
    .B(_5698_),
    .C(_5694_),
    .Y(_5699_)
);

INVX1 _12557_ (
    .A(_5698_),
    .Y(_5700_)
);

NAND3X1 _12558_ (
    .A(_5628_),
    .B(_5655_),
    .C(_5633_),
    .Y(_5701_)
);

OAI21X1 _12559_ (
    .A(_5676_),
    .B(_5701_),
    .C(_5365__bF$buf1),
    .Y(_5702_)
);

NAND2X1 _12560_ (
    .A(_5700_),
    .B(_5702_),
    .Y(_5703_)
);

NAND3X1 _12561_ (
    .A(\genblk1[6].u_ce.Xin12b [5]),
    .B(_5703_),
    .C(_5699_),
    .Y(_5704_)
);

NAND3X1 _12562_ (
    .A(_5365__bF$buf0),
    .B(_5700_),
    .C(_5694_),
    .Y(_5705_)
);

NAND2X1 _12563_ (
    .A(_5698_),
    .B(_5702_),
    .Y(_5706_)
);

NAND3X1 _12564_ (
    .A(_5317_),
    .B(_5706_),
    .C(_5705_),
    .Y(_5707_)
);

NAND2X1 _12565_ (
    .A(_5704_),
    .B(_5707_),
    .Y(_5708_)
);

AOI21X1 _12566_ (
    .A(_5686_),
    .B(_5681_),
    .C(_5708_),
    .Y(_5709_)
);

OAI21X1 _12567_ (
    .A(_5691_),
    .B(_5690_),
    .C(_5681_),
    .Y(_5710_)
);

AND2X2 _12568_ (
    .A(_5704_),
    .B(_5707_),
    .Y(_5711_)
);

OAI21X1 _12569_ (
    .A(_5711_),
    .B(_5710_),
    .C(_5568_),
    .Y(_5712_)
);

OAI22X1 _12570_ (
    .A(_5266_),
    .B(\genblk1[6].u_ce.Vld ),
    .C(_5709_),
    .D(_5712_),
    .Y(_5183_)
);

NOR2X1 _12571_ (
    .A(_5676_),
    .B(_5701_),
    .Y(_5713_)
);

NAND2X1 _12572_ (
    .A(_5700_),
    .B(_5713_),
    .Y(_5714_)
);

AOI21X1 _12573_ (
    .A(_5276__bF$buf4),
    .B(_5672_),
    .C(_5696_),
    .Y(_5715_)
);

NAND2X1 _12574_ (
    .A(_5303__bF$buf3),
    .B(_5623_),
    .Y(_5716_)
);

OAI21X1 _12575_ (
    .A(_5303__bF$buf2),
    .B(_5715_),
    .C(_5716_),
    .Y(_5717_)
);

NAND3X1 _12576_ (
    .A(_5365__bF$buf5),
    .B(_5717_),
    .C(_5714_),
    .Y(_5718_)
);

NOR3X1 _12577_ (
    .A(_5676_),
    .B(_5698_),
    .C(_5701_),
    .Y(_5719_)
);

INVX1 _12578_ (
    .A(_5717_),
    .Y(_5720_)
);

OAI21X1 _12579_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf1 ),
    .B(_5719_),
    .C(_5720_),
    .Y(_5721_)
);

NAND3X1 _12580_ (
    .A(\genblk1[6].u_ce.Xin12b [6]),
    .B(_5721_),
    .C(_5718_),
    .Y(_5722_)
);

NAND3X1 _12581_ (
    .A(_5365__bF$buf4),
    .B(_5720_),
    .C(_5714_),
    .Y(_5723_)
);

OAI21X1 _12582_ (
    .A(\genblk1[6].u_ce.Ain12b_11_bF$buf0 ),
    .B(_5719_),
    .C(_5717_),
    .Y(_5724_)
);

NAND3X1 _12583_ (
    .A(_5319_),
    .B(_5724_),
    .C(_5723_),
    .Y(_5725_)
);

AND2X2 _12584_ (
    .A(_5722_),
    .B(_5725_),
    .Y(_5726_)
);

NAND2X1 _12585_ (
    .A(_5685_),
    .B(_5711_),
    .Y(_5727_)
);

INVX1 _12586_ (
    .A(_5681_),
    .Y(_5728_)
);

INVX1 _12587_ (
    .A(_5704_),
    .Y(_5729_)
);

AOI21X1 _12588_ (
    .A(_5728_),
    .B(_5707_),
    .C(_5729_),
    .Y(_5730_)
);

OAI21X1 _12589_ (
    .A(_5690_),
    .B(_5727_),
    .C(_5730_),
    .Y(_5731_)
);

AND2X2 _12590_ (
    .A(_5731_),
    .B(_5726_),
    .Y(_5732_)
);

NOR2X1 _12591_ (
    .A(_5726_),
    .B(_5731_),
    .Y(_5733_)
);

OAI21X1 _12592_ (
    .A(_5733_),
    .B(_5732_),
    .C(_5274_),
    .Y(_5734_)
);

NAND2X1 _12593_ (
    .A(\genblk1[6].u_ce.Vld ),
    .B(_5734_),
    .Y(_5735_)
);

OAI21X1 _12594_ (
    .A(_5252_),
    .B(\genblk1[6].u_ce.Vld ),
    .C(_5735_),
    .Y(_5184_)
);

INVX1 _12595_ (
    .A(_5722_),
    .Y(_5736_)
);

NOR2X1 _12596_ (
    .A(_5736_),
    .B(_5732_),
    .Y(_5737_)
);

NAND2X1 _12597_ (
    .A(_5720_),
    .B(_5719_),
    .Y(_5738_)
);

NOR2X1 _12598_ (
    .A(_5303__bF$buf1),
    .B(_5556_),
    .Y(_5739_)
);

AOI21X1 _12599_ (
    .A(_5651_),
    .B(_5303__bF$buf0),
    .C(_5739_),
    .Y(_5740_)
);

NAND3X1 _12600_ (
    .A(_5365__bF$buf3),
    .B(_5740_),
    .C(_5738_),
    .Y(_5741_)
);

INVX1 _12601_ (
    .A(_5741_),
    .Y(_5742_)
);

AOI21X1 _12602_ (
    .A(_5738_),
    .B(_5365__bF$buf2),
    .C(_5740_),
    .Y(_5743_)
);

OAI21X1 _12603_ (
    .A(_5743_),
    .B(_5742_),
    .C(\genblk1[6].u_ce.Xin12b [7]),
    .Y(_5744_)
);

INVX1 _12604_ (
    .A(_5743_),
    .Y(_5745_)
);

NAND3X1 _12605_ (
    .A(_5322_),
    .B(_5741_),
    .C(_5745_),
    .Y(_5746_)
);

AND2X2 _12606_ (
    .A(_5746_),
    .B(_5744_),
    .Y(_5747_)
);

OR2X2 _12607_ (
    .A(_5737_),
    .B(_5747_),
    .Y(_5748_)
);

AOI21X1 _12608_ (
    .A(_5737_),
    .B(_5747_),
    .C(_5567_),
    .Y(_5749_)
);

AOI22X1 _12609_ (
    .A(_5265_),
    .B(_5270__bF$buf0),
    .C(_5748_),
    .D(_5749_),
    .Y(_5185_)
);

NOR2X1 _12610_ (
    .A(_5691_),
    .B(_5708_),
    .Y(_5750_)
);

OAI21X1 _12611_ (
    .A(_5681_),
    .B(_5708_),
    .C(_5704_),
    .Y(_5751_)
);

AOI21X1 _12612_ (
    .A(_5750_),
    .B(_5670_),
    .C(_5751_),
    .Y(_5752_)
);

AOI21X1 _12613_ (
    .A(_5745_),
    .B(_5741_),
    .C(_5322_),
    .Y(_5753_)
);

AOI21X1 _12614_ (
    .A(_5736_),
    .B(_5746_),
    .C(_5753_),
    .Y(_5754_)
);

NAND3X1 _12615_ (
    .A(_5726_),
    .B(_5744_),
    .C(_5746_),
    .Y(_5755_)
);

OAI21X1 _12616_ (
    .A(_5755_),
    .B(_5752_),
    .C(_5754_),
    .Y(_5756_)
);

NAND3X1 _12617_ (
    .A(_5720_),
    .B(_5740_),
    .C(_5719_),
    .Y(_5757_)
);

INVX1 _12618_ (
    .A(_5674_),
    .Y(_5758_)
);

INVX1 _12619_ (
    .A(_5739_),
    .Y(_5759_)
);

OAI21X1 _12620_ (
    .A(1'h1),
    .B(_5758_),
    .C(_5759_),
    .Y(_5760_)
);

INVX1 _12621_ (
    .A(_5760_),
    .Y(_5761_)
);

NAND3X1 _12622_ (
    .A(_5365__bF$buf1),
    .B(_5761_),
    .C(_5757_),
    .Y(_5762_)
);

INVX1 _12623_ (
    .A(_5762_),
    .Y(_5763_)
);

AOI21X1 _12624_ (
    .A(_5757_),
    .B(_5365__bF$buf0),
    .C(_5761_),
    .Y(_5764_)
);

OAI21X1 _12625_ (
    .A(_5764_),
    .B(_5763_),
    .C(\genblk1[6].u_ce.Xin12b [8]),
    .Y(_5765_)
);

INVX1 _12626_ (
    .A(_5764_),
    .Y(_5766_)
);

NAND3X1 _12627_ (
    .A(_5324_),
    .B(_5762_),
    .C(_5766_),
    .Y(_5767_)
);

AND2X2 _12628_ (
    .A(_5767_),
    .B(_5765_),
    .Y(_5768_)
);

OR2X2 _12629_ (
    .A(_5756_),
    .B(_5768_),
    .Y(_5769_)
);

INVX1 _12630_ (
    .A(_5769_),
    .Y(_5770_)
);

NAND2X1 _12631_ (
    .A(_5768_),
    .B(_5756_),
    .Y(_5771_)
);

NAND2X1 _12632_ (
    .A(_5568_),
    .B(_5771_),
    .Y(_5772_)
);

OAI22X1 _12633_ (
    .A(_5254_),
    .B(\genblk1[6].u_ce.Vld ),
    .C(_5772_),
    .D(_5770_),
    .Y(_5186_)
);

NOR3X1 _12634_ (
    .A(_5698_),
    .B(_5717_),
    .C(_5694_),
    .Y(_5773_)
);

NAND3X1 _12635_ (
    .A(_5740_),
    .B(_5761_),
    .C(_5773_),
    .Y(_5774_)
);

OR2X2 _12636_ (
    .A(_5695_),
    .B(_5696_),
    .Y(_5775_)
);

AOI21X1 _12637_ (
    .A(_5775_),
    .B(_5303__bF$buf3),
    .C(_5739_),
    .Y(_5776_)
);

INVX1 _12638_ (
    .A(_5776_),
    .Y(_5777_)
);

NAND3X1 _12639_ (
    .A(_5365__bF$buf5),
    .B(_5777_),
    .C(_5774_),
    .Y(_5778_)
);

OAI21X1 _12640_ (
    .A(_5760_),
    .B(_5757_),
    .C(_5365__bF$buf4),
    .Y(_5779_)
);

NAND2X1 _12641_ (
    .A(_5776_),
    .B(_5779_),
    .Y(_5780_)
);

NAND3X1 _12642_ (
    .A(\genblk1[6].u_ce.Xin12b [9]),
    .B(_5780_),
    .C(_5778_),
    .Y(_5781_)
);

NAND3X1 _12643_ (
    .A(_5365__bF$buf3),
    .B(_5776_),
    .C(_5774_),
    .Y(_5782_)
);

NAND2X1 _12644_ (
    .A(_5777_),
    .B(_5779_),
    .Y(_5783_)
);

NAND3X1 _12645_ (
    .A(_5369_),
    .B(_5783_),
    .C(_5782_),
    .Y(_5784_)
);

NAND2X1 _12646_ (
    .A(_5781_),
    .B(_5784_),
    .Y(_5785_)
);

AOI21X1 _12647_ (
    .A(_5771_),
    .B(_5765_),
    .C(_5785_),
    .Y(_5786_)
);

NAND3X1 _12648_ (
    .A(_5765_),
    .B(_5785_),
    .C(_5771_),
    .Y(_5787_)
);

NAND2X1 _12649_ (
    .A(_5568_),
    .B(_5787_),
    .Y(_5788_)
);

OAI22X1 _12650_ (
    .A(_5262_),
    .B(\genblk1[6].u_ce.Vld ),
    .C(_5786_),
    .D(_5788_),
    .Y(_5187_)
);

NAND2X1 _12651_ (
    .A(\genblk1[6].u_ce.Xcalc [10]),
    .B(_5270__bF$buf3),
    .Y(_5789_)
);

OAI21X1 _12652_ (
    .A(1'h1),
    .B(_5715_),
    .C(_5759_),
    .Y(_5790_)
);

OAI21X1 _12653_ (
    .A(_5777_),
    .B(_5774_),
    .C(_5365__bF$buf2),
    .Y(_5791_)
);

NOR2X1 _12654_ (
    .A(_5790_),
    .B(_5791_),
    .Y(_5792_)
);

NAND2X1 _12655_ (
    .A(_5790_),
    .B(_5791_),
    .Y(_5793_)
);

INVX1 _12656_ (
    .A(_5793_),
    .Y(_5794_)
);

OAI21X1 _12657_ (
    .A(_5792_),
    .B(_5794_),
    .C(\genblk1[6].u_ce.Xin12b [10]),
    .Y(_5795_)
);

INVX1 _12658_ (
    .A(_5792_),
    .Y(_5796_)
);

NAND3X1 _12659_ (
    .A(_5399_),
    .B(_5793_),
    .C(_5796_),
    .Y(_5797_)
);

AND2X2 _12660_ (
    .A(_5797_),
    .B(_5795_),
    .Y(_5798_)
);

OAI21X1 _12661_ (
    .A(_5765_),
    .B(_5785_),
    .C(_5781_),
    .Y(_5799_)
);

NAND3X1 _12662_ (
    .A(_5726_),
    .B(_5731_),
    .C(_5747_),
    .Y(_5800_)
);

NAND3X1 _12663_ (
    .A(_5781_),
    .B(_5784_),
    .C(_5768_),
    .Y(_5801_)
);

AOI21X1 _12664_ (
    .A(_5800_),
    .B(_5754_),
    .C(_5801_),
    .Y(_5802_)
);

OAI21X1 _12665_ (
    .A(_5799_),
    .B(_5802_),
    .C(_5798_),
    .Y(_5803_)
);

NAND2X1 _12666_ (
    .A(_5795_),
    .B(_5797_),
    .Y(_5804_)
);

NAND2X1 _12667_ (
    .A(_5765_),
    .B(_5767_),
    .Y(_5805_)
);

NOR2X1 _12668_ (
    .A(_5805_),
    .B(_5785_),
    .Y(_5806_)
);

AOI21X1 _12669_ (
    .A(_5756_),
    .B(_5806_),
    .C(_5799_),
    .Y(_5807_)
);

NAND2X1 _12670_ (
    .A(_5804_),
    .B(_5807_),
    .Y(_5808_)
);

AOI21X1 _12671_ (
    .A(_5803_),
    .B(_5808_),
    .C(_5275_),
    .Y(_5809_)
);

OAI21X1 _12672_ (
    .A(_5270__bF$buf2),
    .B(_5809_),
    .C(_5789_),
    .Y(_5188_)
);

NAND2X1 _12673_ (
    .A(\genblk1[6].u_ce.Xcalc [11]),
    .B(_5270__bF$buf1),
    .Y(_5810_)
);

OR2X2 _12674_ (
    .A(_5774_),
    .B(_5777_),
    .Y(_5811_)
);

OAI21X1 _12675_ (
    .A(_5790_),
    .B(_5811_),
    .C(_5365__bF$buf1),
    .Y(_5812_)
);

OR2X2 _12676_ (
    .A(_5812_),
    .B(_5558_),
    .Y(_5813_)
);

NAND2X1 _12677_ (
    .A(_5558_),
    .B(_5812_),
    .Y(_5814_)
);

AOI22X1 _12678_ (
    .A(_5813_),
    .B(_5814_),
    .C(_5803_),
    .D(_5795_),
    .Y(_5815_)
);

OAI21X1 _12679_ (
    .A(_5804_),
    .B(_5807_),
    .C(_5795_),
    .Y(_5816_)
);

NAND2X1 _12680_ (
    .A(_5814_),
    .B(_5813_),
    .Y(_5817_)
);

OAI21X1 _12681_ (
    .A(_5817_),
    .B(_5816_),
    .C(_5568_),
    .Y(_5818_)
);

OAI21X1 _12682_ (
    .A(_5815_),
    .B(_5818_),
    .C(_5810_),
    .Y(_5189_)
);

INVX1 _12683_ (
    .A(_5224_),
    .Y(_5819_)
);

NAND3X1 _12684_ (
    .A(_5261_),
    .B(\genblk1[6].u_ce.LoadCtl [5]),
    .C(_5228_),
    .Y(_5820_)
);

NOR2X1 _12685_ (
    .A(_5819_),
    .B(_5820_),
    .Y(_5821_)
);

NAND2X1 _12686_ (
    .A(\genblk1[5].u_ce.X_ [0]),
    .B(_5821_),
    .Y(_5822_)
);

OAI21X1 _12687_ (
    .A(_5399_),
    .B(_5821_),
    .C(_5822_),
    .Y(_5190_)
);

NAND2X1 _12688_ (
    .A(\genblk1[5].u_ce.X_ [1]),
    .B(_5821_),
    .Y(_5823_)
);

OAI21X1 _12689_ (
    .A(_5424_),
    .B(_5821_),
    .C(_5823_),
    .Y(_5191_)
);

INVX1 _12690_ (
    .A(\genblk1[5].u_ce.X_ [0]),
    .Y(_5824_)
);

NAND3X1 _12691_ (
    .A(\genblk1[6].u_ce.LoadCtl [4]),
    .B(_5224_),
    .C(_5228_),
    .Y(_5825_)
);

NAND2X1 _12692_ (
    .A(\genblk1[6].u_ce.Xin12b [8]),
    .B(_5825_),
    .Y(_5826_)
);

OAI21X1 _12693_ (
    .A(_5824_),
    .B(_5825_),
    .C(_5826_),
    .Y(_5192_)
);

INVX1 _12694_ (
    .A(\genblk1[5].u_ce.X_ [1]),
    .Y(_5827_)
);

NAND2X1 _12695_ (
    .A(\genblk1[6].u_ce.Xin12b [9]),
    .B(_5825_),
    .Y(_5828_)
);

OAI21X1 _12696_ (
    .A(_5827_),
    .B(_5825_),
    .C(_5828_),
    .Y(_5193_)
);

NAND2X1 _12697_ (
    .A(_5228_),
    .B(_5227_),
    .Y(_5829_)
);

OAI21X1 _12698_ (
    .A(_5229_),
    .B(_5232_),
    .C(\genblk1[6].u_ce.Xin12b [6]),
    .Y(_5830_)
);

OAI21X1 _12699_ (
    .A(_5824_),
    .B(_5829_),
    .C(_5830_),
    .Y(_5194_)
);

OAI21X1 _12700_ (
    .A(_5229_),
    .B(_5232_),
    .C(\genblk1[6].u_ce.Xin12b [7]),
    .Y(_5831_)
);

OAI21X1 _12701_ (
    .A(_5827_),
    .B(_5829_),
    .C(_5831_),
    .Y(_5195_)
);

NOR2X1 _12702_ (
    .A(_5225_),
    .B(_5229_),
    .Y(_5832_)
);

NAND2X1 _12703_ (
    .A(\genblk1[5].u_ce.X_ [0]),
    .B(_5832_),
    .Y(_5833_)
);

OAI21X1 _12704_ (
    .A(_5309_),
    .B(_5832_),
    .C(_5833_),
    .Y(_5196_)
);

NAND2X1 _12705_ (
    .A(\genblk1[5].u_ce.X_ [1]),
    .B(_5832_),
    .Y(_5834_)
);

OAI21X1 _12706_ (
    .A(_5317_),
    .B(_5832_),
    .C(_5834_),
    .Y(_5197_)
);

OAI21X1 _12707_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_5230_),
    .C(\genblk1[6].u_ce.Xin1 [0]),
    .Y(_5835_)
);

OAI21X1 _12708_ (
    .A(_5824_),
    .B(_5250_),
    .C(_5835_),
    .Y(_5198_)
);

OAI21X1 _12709_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_5230_),
    .C(\genblk1[6].u_ce.Xin1 [1]),
    .Y(_5836_)
);

OAI21X1 _12710_ (
    .A(_5827_),
    .B(_5250_),
    .C(_5836_),
    .Y(_5199_)
);

NAND2X1 _12711_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[5].u_ce.X_ [0]),
    .Y(_5837_)
);

OAI21X1 _12712_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_5332_),
    .C(_5837_),
    .Y(_5200_)
);

NAND2X1 _12713_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[5].u_ce.X_ [1]),
    .Y(_5838_)
);

OAI21X1 _12714_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_5312_),
    .C(_5838_),
    .Y(_5201_)
);

NAND2X1 _12715_ (
    .A(\genblk1[5].u_ce.Y_ [0]),
    .B(_5821_),
    .Y(_5839_)
);

OAI21X1 _12716_ (
    .A(_5532_),
    .B(_5821_),
    .C(_5839_),
    .Y(_5202_)
);

NAND2X1 _12717_ (
    .A(\genblk1[5].u_ce.Y_ [1]),
    .B(_5821_),
    .Y(_5840_)
);

OAI21X1 _12718_ (
    .A(_5556_),
    .B(_5821_),
    .C(_5840_),
    .Y(_5203_)
);

INVX1 _12719_ (
    .A(\genblk1[5].u_ce.Y_ [0]),
    .Y(_5841_)
);

NAND2X1 _12720_ (
    .A(\genblk1[6].u_ce.Yin12b [8]),
    .B(_5825_),
    .Y(_5842_)
);

OAI21X1 _12721_ (
    .A(_5841_),
    .B(_5825_),
    .C(_5842_),
    .Y(_5204_)
);

INVX1 _12722_ (
    .A(\genblk1[5].u_ce.Y_ [1]),
    .Y(_5843_)
);

NAND2X1 _12723_ (
    .A(\genblk1[6].u_ce.Yin12b [9]),
    .B(_5825_),
    .Y(_5844_)
);

OAI21X1 _12724_ (
    .A(_5843_),
    .B(_5825_),
    .C(_5844_),
    .Y(_5205_)
);

OAI21X1 _12725_ (
    .A(_5229_),
    .B(_5232_),
    .C(\genblk1[6].u_ce.Yin12b [6]),
    .Y(_5215_)
);

OAI21X1 _12726_ (
    .A(_5841_),
    .B(_5829_),
    .C(_5215_),
    .Y(_5206_)
);

OAI21X1 _12727_ (
    .A(_5229_),
    .B(_5232_),
    .C(\genblk1[6].u_ce.Yin12b [7]),
    .Y(_5216_)
);

OAI21X1 _12728_ (
    .A(_5843_),
    .B(_5829_),
    .C(_5216_),
    .Y(_5207_)
);

NAND2X1 _12729_ (
    .A(\genblk1[5].u_ce.Y_ [0]),
    .B(_5832_),
    .Y(_5217_)
);

OAI21X1 _12730_ (
    .A(_5397_),
    .B(_5832_),
    .C(_5217_),
    .Y(_5208_)
);

NAND2X1 _12731_ (
    .A(\genblk1[5].u_ce.Y_ [1]),
    .B(_5832_),
    .Y(_5218_)
);

OAI21X1 _12732_ (
    .A(_5422_),
    .B(_5832_),
    .C(_5218_),
    .Y(_5209_)
);

OAI21X1 _12733_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_5230_),
    .C(\genblk1[6].u_ce.Yin1 [0]),
    .Y(_5219_)
);

OAI21X1 _12734_ (
    .A(_5841_),
    .B(_5250_),
    .C(_5219_),
    .Y(_5210_)
);

OAI21X1 _12735_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_5230_),
    .C(\genblk1[6].u_ce.Yin1 [1]),
    .Y(_5220_)
);

OAI21X1 _12736_ (
    .A(_5843_),
    .B(_5250_),
    .C(_5220_),
    .Y(_5211_)
);

NAND2X1 _12737_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[5].u_ce.Y_ [0]),
    .Y(_5221_)
);

OAI21X1 _12738_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_5569_),
    .C(_5221_),
    .Y(_5212_)
);

NAND2X1 _12739_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[5].u_ce.Y_ [1]),
    .Y(_5222_)
);

OAI21X1 _12740_ (
    .A(\genblk1[6].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_5354_),
    .C(_5222_),
    .Y(_5213_)
);

NAND2X1 _12741_ (
    .A(\a[6] [1]),
    .B(_5821_),
    .Y(_5223_)
);

OAI21X1 _12742_ (
    .A(_5365__bF$buf0),
    .B(_5821_),
    .C(_5223_),
    .Y(_5214_)
);

DFFPOSX1 _12743_ (
    .CLK(clk_bF$buf51),
    .D(_5166_),
    .Q(\genblk1[6].u_ce.Ycalc [2])
);

DFFPOSX1 _12744_ (
    .CLK(clk_bF$buf50),
    .D(_5167_),
    .Q(\genblk1[6].u_ce.Ycalc [3])
);

DFFPOSX1 _12745_ (
    .CLK(clk_bF$buf49),
    .D(_5168_),
    .Q(\genblk1[6].u_ce.Ycalc [4])
);

DFFPOSX1 _12746_ (
    .CLK(clk_bF$buf48),
    .D(_5169_),
    .Q(\genblk1[6].u_ce.Ycalc [5])
);

DFFPOSX1 _12747_ (
    .CLK(clk_bF$buf47),
    .D(_5170_),
    .Q(\genblk1[6].u_ce.Ycalc [6])
);

DFFPOSX1 _12748_ (
    .CLK(clk_bF$buf46),
    .D(_5171_),
    .Q(\genblk1[6].u_ce.Ycalc [7])
);

DFFPOSX1 _12749_ (
    .CLK(clk_bF$buf45),
    .D(_5172_),
    .Q(\genblk1[6].u_ce.Ycalc [8])
);

DFFPOSX1 _12750_ (
    .CLK(clk_bF$buf44),
    .D(_5173_),
    .Q(\genblk1[6].u_ce.Ycalc [9])
);

DFFPOSX1 _12751_ (
    .CLK(clk_bF$buf43),
    .D(_5174_),
    .Q(\genblk1[6].u_ce.Ycalc [10])
);

DFFPOSX1 _12752_ (
    .CLK(clk_bF$buf42),
    .D(_5175_),
    .Q(\genblk1[6].u_ce.Ycalc [11])
);

DFFPOSX1 _12753_ (
    .CLK(clk_bF$buf41),
    .D(_5176_),
    .Q(\genblk1[6].u_ce.Ycalc [0])
);

DFFPOSX1 _12754_ (
    .CLK(clk_bF$buf40),
    .D(_5177_),
    .Q(\genblk1[6].u_ce.Ycalc [1])
);

DFFPOSX1 _12755_ (
    .CLK(clk_bF$buf39),
    .D(_5178_),
    .Q(\genblk1[6].u_ce.Xcalc [0])
);

DFFPOSX1 _12756_ (
    .CLK(clk_bF$buf38),
    .D(_5179_),
    .Q(\genblk1[6].u_ce.Xcalc [1])
);

DFFPOSX1 _12757_ (
    .CLK(clk_bF$buf37),
    .D(_5180_),
    .Q(\genblk1[6].u_ce.Xcalc [2])
);

DFFPOSX1 _12758_ (
    .CLK(clk_bF$buf36),
    .D(_5181_),
    .Q(\genblk1[6].u_ce.Xcalc [3])
);

DFFPOSX1 _12759_ (
    .CLK(clk_bF$buf35),
    .D(_5182_),
    .Q(\genblk1[6].u_ce.Xcalc [4])
);

DFFPOSX1 _12760_ (
    .CLK(clk_bF$buf34),
    .D(_5183_),
    .Q(\genblk1[6].u_ce.Xcalc [5])
);

DFFPOSX1 _12761_ (
    .CLK(clk_bF$buf33),
    .D(_5184_),
    .Q(\genblk1[6].u_ce.Xcalc [6])
);

DFFPOSX1 _12762_ (
    .CLK(clk_bF$buf32),
    .D(_5185_),
    .Q(\genblk1[6].u_ce.Xcalc [7])
);

DFFPOSX1 _12763_ (
    .CLK(clk_bF$buf31),
    .D(_5186_),
    .Q(\genblk1[6].u_ce.Xcalc [8])
);

DFFPOSX1 _12764_ (
    .CLK(clk_bF$buf30),
    .D(_5187_),
    .Q(\genblk1[6].u_ce.Xcalc [9])
);

DFFPOSX1 _12765_ (
    .CLK(clk_bF$buf29),
    .D(_5188_),
    .Q(\genblk1[6].u_ce.Xcalc [10])
);

DFFPOSX1 _12766_ (
    .CLK(clk_bF$buf28),
    .D(_5189_),
    .Q(\genblk1[6].u_ce.Xcalc [11])
);

DFFPOSX1 _12767_ (
    .CLK(clk_bF$buf27),
    .D(_5190_),
    .Q(\genblk1[6].u_ce.Xin12b [10])
);

DFFPOSX1 _12768_ (
    .CLK(clk_bF$buf26),
    .D(_5191_),
    .Q(\genblk1[6].u_ce.Xin12b [11])
);

DFFPOSX1 _12769_ (
    .CLK(clk_bF$buf25),
    .D(_5192_),
    .Q(\genblk1[6].u_ce.Xin12b [8])
);

DFFPOSX1 _12770_ (
    .CLK(clk_bF$buf24),
    .D(_5193_),
    .Q(\genblk1[6].u_ce.Xin12b [9])
);

DFFPOSX1 _12771_ (
    .CLK(clk_bF$buf23),
    .D(_5194_),
    .Q(\genblk1[6].u_ce.Xin12b [6])
);

DFFPOSX1 _12772_ (
    .CLK(clk_bF$buf22),
    .D(_5195_),
    .Q(\genblk1[6].u_ce.Xin12b [7])
);

DFFPOSX1 _12773_ (
    .CLK(clk_bF$buf21),
    .D(_5196_),
    .Q(\genblk1[6].u_ce.Xin12b [4])
);

DFFPOSX1 _12774_ (
    .CLK(clk_bF$buf20),
    .D(_5197_),
    .Q(\genblk1[6].u_ce.Xin12b [5])
);

DFFPOSX1 _12775_ (
    .CLK(clk_bF$buf19),
    .D(_5198_),
    .Q(\genblk1[6].u_ce.Xin1 [0])
);

DFFPOSX1 _12776_ (
    .CLK(clk_bF$buf18),
    .D(_5199_),
    .Q(\genblk1[6].u_ce.Xin1 [1])
);

DFFPOSX1 _12777_ (
    .CLK(clk_bF$buf17),
    .D(_5200_),
    .Q(\genblk1[6].u_ce.Xin0 [0])
);

DFFPOSX1 _12778_ (
    .CLK(clk_bF$buf16),
    .D(_5201_),
    .Q(\genblk1[6].u_ce.Xin0 [1])
);

DFFPOSX1 _12779_ (
    .CLK(clk_bF$buf15),
    .D(_5202_),
    .Q(\genblk1[6].u_ce.Yin12b [10])
);

DFFPOSX1 _12780_ (
    .CLK(clk_bF$buf14),
    .D(_5203_),
    .Q(\genblk1[6].u_ce.Yin12b [11])
);

DFFPOSX1 _12781_ (
    .CLK(clk_bF$buf13),
    .D(_5204_),
    .Q(\genblk1[6].u_ce.Yin12b [8])
);

DFFPOSX1 _12782_ (
    .CLK(clk_bF$buf12),
    .D(_5205_),
    .Q(\genblk1[6].u_ce.Yin12b [9])
);

DFFPOSX1 _12783_ (
    .CLK(clk_bF$buf11),
    .D(_5206_),
    .Q(\genblk1[6].u_ce.Yin12b [6])
);

DFFPOSX1 _12784_ (
    .CLK(clk_bF$buf10),
    .D(_5207_),
    .Q(\genblk1[6].u_ce.Yin12b [7])
);

DFFPOSX1 _12785_ (
    .CLK(clk_bF$buf9),
    .D(_5208_),
    .Q(\genblk1[6].u_ce.Yin12b [4])
);

DFFPOSX1 _12786_ (
    .CLK(clk_bF$buf8),
    .D(_5209_),
    .Q(\genblk1[6].u_ce.Yin12b [5])
);

DFFPOSX1 _12787_ (
    .CLK(clk_bF$buf7),
    .D(_5210_),
    .Q(\genblk1[6].u_ce.Yin1 [0])
);

DFFPOSX1 _12788_ (
    .CLK(clk_bF$buf6),
    .D(_5211_),
    .Q(\genblk1[6].u_ce.Yin1 [1])
);

DFFPOSX1 _12789_ (
    .CLK(clk_bF$buf5),
    .D(_5212_),
    .Q(\genblk1[6].u_ce.Yin0 [0])
);

DFFPOSX1 _12790_ (
    .CLK(clk_bF$buf4),
    .D(_5213_),
    .Q(\genblk1[6].u_ce.Yin0 [1])
);

DFFPOSX1 _12791_ (
    .CLK(clk_bF$buf3),
    .D(_5214_),
    .Q(\genblk1[6].u_ce.Ain12b [11])
);

DFFPOSX1 _12792_ (
    .CLK(clk_bF$buf2),
    .D(\genblk1[5].u_ce.ISout ),
    .Q(\genblk1[6].u_ce.ISpipe [0])
);

DFFPOSX1 _12793_ (
    .CLK(clk_bF$buf1),
    .D(\genblk1[6].u_ce.ISpipe [0]),
    .Q(\genblk1[6].u_ce.ISpipe [1])
);

DFFPOSX1 _12794_ (
    .CLK(clk_bF$buf0),
    .D(\genblk1[6].u_ce.ISpipe [1]),
    .Q(\genblk1[6].u_ce.ISpipe [2])
);

DFFPOSX1 _12795_ (
    .CLK(clk_bF$buf75),
    .D(\genblk1[6].u_ce.ISpipe [2]),
    .Q(\genblk1[6].u_ce.ISpipe [3])
);

DFFPOSX1 _12796_ (
    .CLK(clk_bF$buf74),
    .D(\genblk1[6].u_ce.ISpipe [3]),
    .Q(\genblk1[6].u_ce.ISpipe [4])
);

DFFPOSX1 _12797_ (
    .CLK(clk_bF$buf73),
    .D(\genblk1[6].u_ce.ISpipe [4]),
    .Q(\genblk1[6].u_ce.ISpipe [5])
);

DFFPOSX1 _12798_ (
    .CLK(clk_bF$buf72),
    .D(\genblk1[6].u_ce.ISpipe [5]),
    .Q(\genblk1[6].u_ce.ISout )
);

DFFPOSX1 _12799_ (
    .CLK(clk_bF$buf71),
    .D(\genblk1[5].u_ce.Vld_bF$buf2 ),
    .Q(\genblk1[6].u_ce.LoadCtl [0])
);

DFFPOSX1 _12800_ (
    .CLK(clk_bF$buf70),
    .D(\genblk1[6].u_ce.LoadCtl_0_bF$buf1 ),
    .Q(\genblk1[6].u_ce.LoadCtl [1])
);

DFFPOSX1 _12801_ (
    .CLK(clk_bF$buf69),
    .D(\genblk1[6].u_ce.LoadCtl [1]),
    .Q(\genblk1[6].u_ce.LoadCtl [2])
);

DFFPOSX1 _12802_ (
    .CLK(clk_bF$buf68),
    .D(\genblk1[6].u_ce.LoadCtl [2]),
    .Q(\genblk1[6].u_ce.LoadCtl [3])
);

DFFPOSX1 _12803_ (
    .CLK(clk_bF$buf67),
    .D(\genblk1[6].u_ce.LoadCtl [3]),
    .Q(\genblk1[6].u_ce.LoadCtl [4])
);

DFFPOSX1 _12804_ (
    .CLK(clk_bF$buf66),
    .D(\genblk1[6].u_ce.LoadCtl [4]),
    .Q(\genblk1[6].u_ce.LoadCtl [5])
);

DFFPOSX1 _12805_ (
    .CLK(clk_bF$buf65),
    .D(\genblk1[6].u_ce.LoadCtl [5]),
    .Q(\genblk1[6].u_ce.Vld )
);

INVX1 _12806_ (
    .A(\u_ot.Ycalc [0]),
    .Y(_5871_)
);

NAND2X1 _12807_ (
    .A(\u_ot.Xcalc [0]),
    .B(selXY_bF$buf3),
    .Y(_5872_)
);

OAI21X1 _12808_ (
    .A(selXY_bF$buf2),
    .B(_5871_),
    .C(_5872_),
    .Y(_6348_[0])
);

INVX1 _12809_ (
    .A(\u_ot.Ycalc [1]),
    .Y(_5873_)
);

NAND2X1 _12810_ (
    .A(selXY_bF$buf1),
    .B(\u_ot.Xcalc [1]),
    .Y(_5874_)
);

OAI21X1 _12811_ (
    .A(selXY_bF$buf0),
    .B(_5873_),
    .C(_5874_),
    .Y(_6348_[1])
);

INVX1 _12812_ (
    .A(\u_ot.Ycalc [2]),
    .Y(_5875_)
);

NAND2X1 _12813_ (
    .A(selXY_bF$buf3),
    .B(\u_ot.Xcalc [2]),
    .Y(_5876_)
);

OAI21X1 _12814_ (
    .A(selXY_bF$buf2),
    .B(_5875_),
    .C(_5876_),
    .Y(_6348_[2])
);

INVX1 _12815_ (
    .A(\u_ot.Ycalc [3]),
    .Y(_5877_)
);

NAND2X1 _12816_ (
    .A(selXY_bF$buf1),
    .B(\u_ot.Xcalc [3]),
    .Y(_5878_)
);

OAI21X1 _12817_ (
    .A(selXY_bF$buf0),
    .B(_5877_),
    .C(_5878_),
    .Y(_6348_[3])
);

INVX1 _12818_ (
    .A(\u_ot.Ycalc [4]),
    .Y(_5879_)
);

NAND2X1 _12819_ (
    .A(selXY_bF$buf3),
    .B(\u_ot.Xcalc [4]),
    .Y(_5880_)
);

OAI21X1 _12820_ (
    .A(selXY_bF$buf2),
    .B(_5879_),
    .C(_5880_),
    .Y(_6348_[4])
);

INVX1 _12821_ (
    .A(\u_ot.Ycalc [5]),
    .Y(_5881_)
);

NAND2X1 _12822_ (
    .A(selXY_bF$buf1),
    .B(\u_ot.Xcalc [5]),
    .Y(_5882_)
);

OAI21X1 _12823_ (
    .A(selXY_bF$buf0),
    .B(_5881_),
    .C(_5882_),
    .Y(_6348_[5])
);

INVX1 _12824_ (
    .A(\u_ot.Ycalc [6]),
    .Y(_5883_)
);

NAND2X1 _12825_ (
    .A(selXY_bF$buf3),
    .B(\u_ot.Xcalc [6]),
    .Y(_5884_)
);

OAI21X1 _12826_ (
    .A(selXY_bF$buf2),
    .B(_5883_),
    .C(_5884_),
    .Y(_6348_[6])
);

INVX1 _12827_ (
    .A(\u_ot.Ycalc [7]),
    .Y(_5885_)
);

NAND2X1 _12828_ (
    .A(selXY_bF$buf1),
    .B(\u_ot.Xcalc [7]),
    .Y(_5886_)
);

OAI21X1 _12829_ (
    .A(selXY_bF$buf0),
    .B(_5885_),
    .C(_5886_),
    .Y(_6348_[7])
);

INVX1 _12830_ (
    .A(\u_ot.Ycalc [8]),
    .Y(_5887_)
);

NAND2X1 _12831_ (
    .A(selXY_bF$buf3),
    .B(\u_ot.Xcalc [8]),
    .Y(_5888_)
);

OAI21X1 _12832_ (
    .A(selXY_bF$buf2),
    .B(_5887_),
    .C(_5888_),
    .Y(_6348_[8])
);

INVX1 _12833_ (
    .A(\u_ot.Ycalc [9]),
    .Y(_5889_)
);

NAND2X1 _12834_ (
    .A(selXY_bF$buf1),
    .B(\u_ot.Xcalc [9]),
    .Y(_5890_)
);

OAI21X1 _12835_ (
    .A(selXY_bF$buf0),
    .B(_5889_),
    .C(_5890_),
    .Y(_6348_[9])
);

INVX1 _12836_ (
    .A(\u_ot.Ycalc [10]),
    .Y(_5891_)
);

NAND2X1 _12837_ (
    .A(selXY_bF$buf3),
    .B(\u_ot.Xcalc [10]),
    .Y(_5892_)
);

OAI21X1 _12838_ (
    .A(selXY_bF$buf2),
    .B(_5891_),
    .C(_5892_),
    .Y(_6348_[10])
);

INVX1 _12839_ (
    .A(\u_ot.Ycalc [11]),
    .Y(_5893_)
);

NAND2X1 _12840_ (
    .A(selXY_bF$buf1),
    .B(\u_ot.Xcalc [11]),
    .Y(_5894_)
);

OAI21X1 _12841_ (
    .A(selXY_bF$buf0),
    .B(_5893_),
    .C(_5894_),
    .Y(_6348_[11])
);

INVX1 _12842_ (
    .A(\u_ot.Yin0 [1]),
    .Y(_5895_)
);

INVX1 _12843_ (
    .A(\u_ot.Yin0 [0]),
    .Y(_5896_)
);

OAI21X1 _12844_ (
    .A(\u_ot.Yin0 [0]),
    .B(\u_ot.Yin0 [1]),
    .C(\u_ot.ISout_bF$buf4 ),
    .Y(_5897_)
);

INVX1 _12845_ (
    .A(_5897_),
    .Y(_5898_)
);

OAI21X1 _12846_ (
    .A(_5896_),
    .B(_5895_),
    .C(_5898_),
    .Y(_5899_)
);

OAI21X1 _12847_ (
    .A(_5895_),
    .B(\u_ot.ISout_bF$buf3 ),
    .C(_5899_),
    .Y(_5846_[1])
);

INVX2 _12848_ (
    .A(\u_ot.ISout_bF$buf2 ),
    .Y(_5900_)
);

NOR2X1 _12849_ (
    .A(\u_ot.Yin0 [0]),
    .B(\u_ot.Yin0 [1]),
    .Y(_5901_)
);

OAI21X1 _12850_ (
    .A(_5900_),
    .B(_5901_),
    .C(\u_ot.Yin1 [0]),
    .Y(_5902_)
);

INVX1 _12851_ (
    .A(\u_ot.Yin1 [0]),
    .Y(_5903_)
);

NAND2X1 _12852_ (
    .A(_5903_),
    .B(_5898_),
    .Y(_5904_)
);

NAND2X1 _12853_ (
    .A(_5902_),
    .B(_5904_),
    .Y(_5846_[2])
);

OAI21X1 _12854_ (
    .A(_5900_),
    .B(_5903_),
    .C(_5897_),
    .Y(_5905_)
);

NAND2X1 _12855_ (
    .A(\u_ot.Yin1 [1]),
    .B(_5905_),
    .Y(_5906_)
);

OR2X2 _12856_ (
    .A(_5905_),
    .B(\u_ot.Yin1 [1]),
    .Y(_5907_)
);

AND2X2 _12857_ (
    .A(_5907_),
    .B(_5906_),
    .Y(_5846_[3])
);

INVX1 _12858_ (
    .A(\u_ot.Yin12b [4]),
    .Y(_5908_)
);

NOR2X1 _12859_ (
    .A(\u_ot.Yin1 [0]),
    .B(\u_ot.Yin1 [1]),
    .Y(_5909_)
);

NAND2X1 _12860_ (
    .A(_5901_),
    .B(_5909_),
    .Y(_5910_)
);

NAND3X1 _12861_ (
    .A(\u_ot.ISout_bF$buf1 ),
    .B(_5908_),
    .C(_5910_),
    .Y(_5911_)
);

AND2X2 _12862_ (
    .A(_5901_),
    .B(_5909_),
    .Y(_5912_)
);

OAI21X1 _12863_ (
    .A(_5900_),
    .B(_5912_),
    .C(\u_ot.Yin12b [4]),
    .Y(_5913_)
);

NAND2X1 _12864_ (
    .A(_5911_),
    .B(_5913_),
    .Y(_5846_[4])
);

OAI21X1 _12865_ (
    .A(\u_ot.Yin12b [4]),
    .B(_5910_),
    .C(\u_ot.ISout_bF$buf0 ),
    .Y(_5914_)
);

NAND2X1 _12866_ (
    .A(\u_ot.Yin12b [5]),
    .B(_5914_),
    .Y(_5915_)
);

OR2X2 _12867_ (
    .A(_5914_),
    .B(\u_ot.Yin12b [5]),
    .Y(_5916_)
);

NAND2X1 _12868_ (
    .A(_5915_),
    .B(_5916_),
    .Y(_5846_[5])
);

INVX1 _12869_ (
    .A(\u_ot.Yin12b [6]),
    .Y(_5917_)
);

NOR2X1 _12870_ (
    .A(\u_ot.Yin12b [4]),
    .B(\u_ot.Yin12b [5]),
    .Y(_5918_)
);

NAND2X1 _12871_ (
    .A(_5918_),
    .B(_5912_),
    .Y(_5919_)
);

NAND3X1 _12872_ (
    .A(\u_ot.ISout_bF$buf4 ),
    .B(_5917_),
    .C(_5919_),
    .Y(_5920_)
);

NAND2X1 _12873_ (
    .A(\u_ot.ISout_bF$buf3 ),
    .B(_5919_),
    .Y(_5921_)
);

NAND2X1 _12874_ (
    .A(\u_ot.Yin12b [6]),
    .B(_5921_),
    .Y(_5922_)
);

NAND2X1 _12875_ (
    .A(_5920_),
    .B(_5922_),
    .Y(_5846_[6])
);

NAND2X1 _12876_ (
    .A(\u_ot.ISout_bF$buf2 ),
    .B(\u_ot.Yin12b [6]),
    .Y(_5923_)
);

NAND3X1 _12877_ (
    .A(\u_ot.Yin12b [7]),
    .B(_5923_),
    .C(_5921_),
    .Y(_5924_)
);

INVX1 _12878_ (
    .A(\u_ot.Yin12b [7]),
    .Y(_5925_)
);

NAND3X1 _12879_ (
    .A(_5917_),
    .B(_5918_),
    .C(_5912_),
    .Y(_5926_)
);

NAND3X1 _12880_ (
    .A(\u_ot.ISout_bF$buf1 ),
    .B(_5925_),
    .C(_5926_),
    .Y(_5927_)
);

NAND2X1 _12881_ (
    .A(_5927_),
    .B(_5924_),
    .Y(_5846_[7])
);

NOR2X1 _12882_ (
    .A(\u_ot.Yin12b [6]),
    .B(\u_ot.Yin12b [7]),
    .Y(_5928_)
);

NAND2X1 _12883_ (
    .A(_5918_),
    .B(_5928_),
    .Y(_5929_)
);

OAI21X1 _12884_ (
    .A(_5910_),
    .B(_5929_),
    .C(\u_ot.ISout_bF$buf0 ),
    .Y(_5930_)
);

NAND2X1 _12885_ (
    .A(\u_ot.Yin12b [8]),
    .B(_5930_),
    .Y(_5931_)
);

OR2X2 _12886_ (
    .A(_5930_),
    .B(\u_ot.Yin12b [8]),
    .Y(_5932_)
);

NAND2X1 _12887_ (
    .A(_5931_),
    .B(_5932_),
    .Y(_5846_[8])
);

NAND2X1 _12888_ (
    .A(\u_ot.ISout_bF$buf4 ),
    .B(\u_ot.Yin12b [8]),
    .Y(_5933_)
);

NAND3X1 _12889_ (
    .A(\u_ot.Yin12b [9]),
    .B(_5933_),
    .C(_5930_),
    .Y(_5934_)
);

INVX1 _12890_ (
    .A(\u_ot.Yin12b [9]),
    .Y(_5935_)
);

NAND2X1 _12891_ (
    .A(_5933_),
    .B(_5930_),
    .Y(_5936_)
);

NAND2X1 _12892_ (
    .A(_5935_),
    .B(_5936_),
    .Y(_5937_)
);

NAND2X1 _12893_ (
    .A(_5934_),
    .B(_5937_),
    .Y(_5846_[9])
);

INVX1 _12894_ (
    .A(\u_ot.Yin12b [10]),
    .Y(_5938_)
);

AND2X2 _12895_ (
    .A(_5918_),
    .B(_5928_),
    .Y(_5939_)
);

NOR2X1 _12896_ (
    .A(\u_ot.Yin12b [8]),
    .B(\u_ot.Yin12b [9]),
    .Y(_5940_)
);

NAND3X1 _12897_ (
    .A(_5940_),
    .B(_5912_),
    .C(_5939_),
    .Y(_5941_)
);

NAND3X1 _12898_ (
    .A(\u_ot.ISout_bF$buf3 ),
    .B(_5938_),
    .C(_5941_),
    .Y(_5942_)
);

NAND2X1 _12899_ (
    .A(\u_ot.ISout_bF$buf2 ),
    .B(_5941_),
    .Y(_5943_)
);

NAND2X1 _12900_ (
    .A(\u_ot.Yin12b [10]),
    .B(_5943_),
    .Y(_5944_)
);

NAND2X1 _12901_ (
    .A(_5942_),
    .B(_5944_),
    .Y(_5846_[10])
);

INVX1 _12902_ (
    .A(\u_ot.Yin12b [11]),
    .Y(_5945_)
);

NAND2X1 _12903_ (
    .A(\u_ot.ISout_bF$buf1 ),
    .B(\u_ot.Yin12b [10]),
    .Y(_5946_)
);

NAND3X1 _12904_ (
    .A(_5945_),
    .B(_5946_),
    .C(_5943_),
    .Y(_5947_)
);

OAI21X1 _12905_ (
    .A(\u_ot.Yin12b [8]),
    .B(\u_ot.Yin12b [9]),
    .C(\u_ot.ISout_bF$buf0 ),
    .Y(_5948_)
);

NAND3X1 _12906_ (
    .A(_5948_),
    .B(_5946_),
    .C(_5930_),
    .Y(_5949_)
);

NAND2X1 _12907_ (
    .A(\u_ot.Yin12b [11]),
    .B(_5949_),
    .Y(_5950_)
);

NAND2X1 _12908_ (
    .A(_5950_),
    .B(_5947_),
    .Y(_5846_[11])
);

INVX1 _12909_ (
    .A(\u_ot.Xin0 [1]),
    .Y(_5951_)
);

INVX1 _12910_ (
    .A(\u_ot.Xin0 [0]),
    .Y(_5952_)
);

OAI21X1 _12911_ (
    .A(\u_ot.Xin0 [0]),
    .B(\u_ot.Xin0 [1]),
    .C(\u_ot.ISout_bF$buf4 ),
    .Y(_5953_)
);

INVX1 _12912_ (
    .A(_5953_),
    .Y(_5954_)
);

OAI21X1 _12913_ (
    .A(_5952_),
    .B(_5951_),
    .C(_5954_),
    .Y(_5955_)
);

OAI21X1 _12914_ (
    .A(\u_ot.ISout_bF$buf3 ),
    .B(_5951_),
    .C(_5955_),
    .Y(_5845_[1])
);

NOR2X1 _12915_ (
    .A(\u_ot.Xin0 [0]),
    .B(\u_ot.Xin0 [1]),
    .Y(_5956_)
);

OAI21X1 _12916_ (
    .A(_5900_),
    .B(_5956_),
    .C(\u_ot.Xin1 [0]),
    .Y(_5957_)
);

INVX1 _12917_ (
    .A(\u_ot.Xin1 [0]),
    .Y(_5958_)
);

NAND2X1 _12918_ (
    .A(_5958_),
    .B(_5954_),
    .Y(_5959_)
);

NAND2X1 _12919_ (
    .A(_5957_),
    .B(_5959_),
    .Y(_5845_[2])
);

OAI21X1 _12920_ (
    .A(_5900_),
    .B(_5958_),
    .C(_5953_),
    .Y(_5960_)
);

NAND2X1 _12921_ (
    .A(\u_ot.Xin1 [1]),
    .B(_5960_),
    .Y(_5961_)
);

OR2X2 _12922_ (
    .A(_5960_),
    .B(\u_ot.Xin1 [1]),
    .Y(_5962_)
);

AND2X2 _12923_ (
    .A(_5962_),
    .B(_5961_),
    .Y(_5845_[3])
);

INVX1 _12924_ (
    .A(\u_ot.Xin12b [4]),
    .Y(_5963_)
);

NOR2X1 _12925_ (
    .A(\u_ot.Xin1 [0]),
    .B(\u_ot.Xin1 [1]),
    .Y(_5964_)
);

NAND2X1 _12926_ (
    .A(_5956_),
    .B(_5964_),
    .Y(_5965_)
);

NAND3X1 _12927_ (
    .A(\u_ot.ISout_bF$buf2 ),
    .B(_5963_),
    .C(_5965_),
    .Y(_5966_)
);

AND2X2 _12928_ (
    .A(_5956_),
    .B(_5964_),
    .Y(_5967_)
);

OAI21X1 _12929_ (
    .A(_5900_),
    .B(_5967_),
    .C(\u_ot.Xin12b [4]),
    .Y(_5968_)
);

NAND2X1 _12930_ (
    .A(_5966_),
    .B(_5968_),
    .Y(_5845_[4])
);

OAI21X1 _12931_ (
    .A(\u_ot.Xin12b [4]),
    .B(_5965_),
    .C(\u_ot.ISout_bF$buf1 ),
    .Y(_5969_)
);

NAND2X1 _12932_ (
    .A(\u_ot.Xin12b [5]),
    .B(_5969_),
    .Y(_5970_)
);

OR2X2 _12933_ (
    .A(_5969_),
    .B(\u_ot.Xin12b [5]),
    .Y(_5971_)
);

NAND2X1 _12934_ (
    .A(_5970_),
    .B(_5971_),
    .Y(_5845_[5])
);

INVX1 _12935_ (
    .A(\u_ot.Xin12b [6]),
    .Y(_5972_)
);

NOR2X1 _12936_ (
    .A(\u_ot.Xin12b [4]),
    .B(\u_ot.Xin12b [5]),
    .Y(_5973_)
);

NAND2X1 _12937_ (
    .A(_5973_),
    .B(_5967_),
    .Y(_5974_)
);

NAND3X1 _12938_ (
    .A(\u_ot.ISout_bF$buf0 ),
    .B(_5972_),
    .C(_5974_),
    .Y(_5975_)
);

NAND2X1 _12939_ (
    .A(\u_ot.ISout_bF$buf4 ),
    .B(_5974_),
    .Y(_5976_)
);

NAND2X1 _12940_ (
    .A(\u_ot.Xin12b [6]),
    .B(_5976_),
    .Y(_5977_)
);

NAND2X1 _12941_ (
    .A(_5975_),
    .B(_5977_),
    .Y(_5845_[6])
);

NAND2X1 _12942_ (
    .A(\u_ot.ISout_bF$buf3 ),
    .B(\u_ot.Xin12b [6]),
    .Y(_5978_)
);

NAND3X1 _12943_ (
    .A(\u_ot.Xin12b [7]),
    .B(_5978_),
    .C(_5976_),
    .Y(_5979_)
);

INVX1 _12944_ (
    .A(\u_ot.Xin12b [7]),
    .Y(_5980_)
);

NAND3X1 _12945_ (
    .A(_5972_),
    .B(_5973_),
    .C(_5967_),
    .Y(_5981_)
);

NAND3X1 _12946_ (
    .A(\u_ot.ISout_bF$buf2 ),
    .B(_5980_),
    .C(_5981_),
    .Y(_5982_)
);

NAND2X1 _12947_ (
    .A(_5982_),
    .B(_5979_),
    .Y(_5845_[7])
);

NOR2X1 _12948_ (
    .A(\u_ot.Xin12b [6]),
    .B(\u_ot.Xin12b [7]),
    .Y(_5983_)
);

NAND2X1 _12949_ (
    .A(_5973_),
    .B(_5983_),
    .Y(_5984_)
);

OAI21X1 _12950_ (
    .A(_5965_),
    .B(_5984_),
    .C(\u_ot.ISout_bF$buf1 ),
    .Y(_5985_)
);

NAND2X1 _12951_ (
    .A(\u_ot.Xin12b [8]),
    .B(_5985_),
    .Y(_5986_)
);

OR2X2 _12952_ (
    .A(_5985_),
    .B(\u_ot.Xin12b [8]),
    .Y(_5987_)
);

NAND2X1 _12953_ (
    .A(_5986_),
    .B(_5987_),
    .Y(_5845_[8])
);

NAND2X1 _12954_ (
    .A(\u_ot.ISout_bF$buf0 ),
    .B(\u_ot.Xin12b [8]),
    .Y(_5988_)
);

NAND3X1 _12955_ (
    .A(\u_ot.Xin12b [9]),
    .B(_5988_),
    .C(_5985_),
    .Y(_5989_)
);

INVX1 _12956_ (
    .A(\u_ot.Xin12b [9]),
    .Y(_5990_)
);

NAND2X1 _12957_ (
    .A(_5988_),
    .B(_5985_),
    .Y(_5991_)
);

NAND2X1 _12958_ (
    .A(_5990_),
    .B(_5991_),
    .Y(_5992_)
);

NAND2X1 _12959_ (
    .A(_5989_),
    .B(_5992_),
    .Y(_5845_[9])
);

INVX1 _12960_ (
    .A(\u_ot.Xin12b [10]),
    .Y(_5993_)
);

AND2X2 _12961_ (
    .A(_5973_),
    .B(_5983_),
    .Y(_5994_)
);

NOR2X1 _12962_ (
    .A(\u_ot.Xin12b [8]),
    .B(\u_ot.Xin12b [9]),
    .Y(_5995_)
);

NAND3X1 _12963_ (
    .A(_5995_),
    .B(_5967_),
    .C(_5994_),
    .Y(_5996_)
);

NAND3X1 _12964_ (
    .A(\u_ot.ISout_bF$buf4 ),
    .B(_5993_),
    .C(_5996_),
    .Y(_5997_)
);

NAND2X1 _12965_ (
    .A(\u_ot.ISout_bF$buf3 ),
    .B(_5996_),
    .Y(_5998_)
);

NAND2X1 _12966_ (
    .A(\u_ot.Xin12b [10]),
    .B(_5998_),
    .Y(_5999_)
);

NAND2X1 _12967_ (
    .A(_5997_),
    .B(_5999_),
    .Y(_5845_[10])
);

INVX1 _12968_ (
    .A(\u_ot.Xin12b [11]),
    .Y(_6000_)
);

NAND2X1 _12969_ (
    .A(\u_ot.ISout_bF$buf2 ),
    .B(\u_ot.Xin12b [10]),
    .Y(_6001_)
);

NAND3X1 _12970_ (
    .A(_6000_),
    .B(_6001_),
    .C(_5998_),
    .Y(_6002_)
);

OAI21X1 _12971_ (
    .A(\u_ot.Xin12b [8]),
    .B(\u_ot.Xin12b [9]),
    .C(\u_ot.ISout_bF$buf1 ),
    .Y(_6003_)
);

NAND3X1 _12972_ (
    .A(_6003_),
    .B(_6001_),
    .C(_5985_),
    .Y(_6004_)
);

NAND2X1 _12973_ (
    .A(\u_ot.Xin12b [11]),
    .B(_6004_),
    .Y(_6005_)
);

NAND2X1 _12974_ (
    .A(_6005_),
    .B(_6002_),
    .Y(_5845_[11])
);

INVX2 _12975_ (
    .A(\u_ot.LoadCtl [1]),
    .Y(_6006_)
);

NOR2X1 _12976_ (
    .A(\u_ot.LoadCtl [2]),
    .B(\u_ot.LoadCtl [0]),
    .Y(_6007_)
);

AND2X2 _12977_ (
    .A(_6007_),
    .B(_6006_),
    .Y(_6008_)
);

INVX1 _12978_ (
    .A(\u_ot.LoadCtl [4]),
    .Y(_6009_)
);

NAND2X1 _12979_ (
    .A(\u_ot.LoadCtl [5]),
    .B(_6009_),
    .Y(_6010_)
);

NOR2X1 _12980_ (
    .A(\u_ot.LoadCtl [3]),
    .B(_6010_),
    .Y(_6011_)
);

AND2X2 _12981_ (
    .A(_6011_),
    .B(_6008_),
    .Y(_6012_)
);

NAND2X1 _12982_ (
    .A(\genblk1[6].u_ce.X_ [0]),
    .B(_6012_),
    .Y(_6013_)
);

OAI21X1 _12983_ (
    .A(_5993_),
    .B(_6012_),
    .C(_6013_),
    .Y(_5847_)
);

NAND2X1 _12984_ (
    .A(\genblk1[6].u_ce.X_ [1]),
    .B(_6012_),
    .Y(_6014_)
);

OAI21X1 _12985_ (
    .A(_6000_),
    .B(_6012_),
    .C(_6014_),
    .Y(_5848_)
);

INVX1 _12986_ (
    .A(\genblk1[6].u_ce.X_ [0]),
    .Y(_6015_)
);

NOR2X1 _12987_ (
    .A(\u_ot.LoadCtl [3]),
    .B(_6009_),
    .Y(_6016_)
);

NAND2X1 _12988_ (
    .A(_6016_),
    .B(_6008_),
    .Y(_6017_)
);

NAND2X1 _12989_ (
    .A(\u_ot.Xin12b [8]),
    .B(_6017_),
    .Y(_6018_)
);

OAI21X1 _12990_ (
    .A(_6015_),
    .B(_6017_),
    .C(_6018_),
    .Y(_5849_)
);

INVX1 _12991_ (
    .A(\genblk1[6].u_ce.X_ [1]),
    .Y(_6019_)
);

NAND2X1 _12992_ (
    .A(\u_ot.Xin12b [9]),
    .B(_6017_),
    .Y(_6020_)
);

OAI21X1 _12993_ (
    .A(_6019_),
    .B(_6017_),
    .C(_6020_),
    .Y(_5850_)
);

NAND2X1 _12994_ (
    .A(\u_ot.LoadCtl [3]),
    .B(_6008_),
    .Y(_6021_)
);

NAND2X1 _12995_ (
    .A(\u_ot.Xin12b [6]),
    .B(_6021_),
    .Y(_6022_)
);

OAI21X1 _12996_ (
    .A(_6015_),
    .B(_6021_),
    .C(_6022_),
    .Y(_5851_)
);

NAND2X1 _12997_ (
    .A(\u_ot.Xin12b [7]),
    .B(_6021_),
    .Y(_6023_)
);

OAI21X1 _12998_ (
    .A(_6019_),
    .B(_6021_),
    .C(_6023_),
    .Y(_5852_)
);

INVX1 _12999_ (
    .A(\u_ot.LoadCtl [0]),
    .Y(_6024_)
);

NAND3X1 _13000_ (
    .A(\u_ot.LoadCtl [2]),
    .B(_6006_),
    .C(_6024_),
    .Y(_6025_)
);

NAND2X1 _13001_ (
    .A(\u_ot.Xin12b [4]),
    .B(_6025_),
    .Y(_6026_)
);

OAI21X1 _13002_ (
    .A(_6015_),
    .B(_6025_),
    .C(_6026_),
    .Y(_5853_)
);

NAND2X1 _13003_ (
    .A(\u_ot.Xin12b [5]),
    .B(_6025_),
    .Y(_6027_)
);

OAI21X1 _13004_ (
    .A(_6019_),
    .B(_6025_),
    .C(_6027_),
    .Y(_5854_)
);

NAND2X1 _13005_ (
    .A(\u_ot.LoadCtl [1]),
    .B(_6024_),
    .Y(_6028_)
);

OAI21X1 _13006_ (
    .A(\u_ot.LoadCtl [0]),
    .B(_6006_),
    .C(\u_ot.Xin1 [0]),
    .Y(_6029_)
);

OAI21X1 _13007_ (
    .A(_6015_),
    .B(_6028_),
    .C(_6029_),
    .Y(_5855_)
);

OAI21X1 _13008_ (
    .A(\u_ot.LoadCtl [0]),
    .B(_6006_),
    .C(\u_ot.Xin1 [1]),
    .Y(_6030_)
);

OAI21X1 _13009_ (
    .A(_6019_),
    .B(_6028_),
    .C(_6030_),
    .Y(_5856_)
);

NAND2X1 _13010_ (
    .A(\u_ot.LoadCtl [0]),
    .B(\genblk1[6].u_ce.X_ [0]),
    .Y(_6031_)
);

OAI21X1 _13011_ (
    .A(\u_ot.LoadCtl [0]),
    .B(_5952_),
    .C(_6031_),
    .Y(_5857_)
);

NAND2X1 _13012_ (
    .A(\u_ot.LoadCtl [0]),
    .B(\genblk1[6].u_ce.X_ [1]),
    .Y(_6032_)
);

OAI21X1 _13013_ (
    .A(\u_ot.LoadCtl [0]),
    .B(_5951_),
    .C(_6032_),
    .Y(_5858_)
);

NAND2X1 _13014_ (
    .A(\genblk1[6].u_ce.Y_ [0]),
    .B(_6012_),
    .Y(_6033_)
);

OAI21X1 _13015_ (
    .A(_5938_),
    .B(_6012_),
    .C(_6033_),
    .Y(_5859_)
);

NAND2X1 _13016_ (
    .A(\genblk1[6].u_ce.Y_ [1]),
    .B(_6012_),
    .Y(_6034_)
);

OAI21X1 _13017_ (
    .A(_5945_),
    .B(_6012_),
    .C(_6034_),
    .Y(_5860_)
);

INVX1 _13018_ (
    .A(\genblk1[6].u_ce.Y_ [0]),
    .Y(_6035_)
);

NAND2X1 _13019_ (
    .A(\u_ot.Yin12b [8]),
    .B(_6017_),
    .Y(_6036_)
);

OAI21X1 _13020_ (
    .A(_6035_),
    .B(_6017_),
    .C(_6036_),
    .Y(_5861_)
);

INVX1 _13021_ (
    .A(\genblk1[6].u_ce.Y_ [1]),
    .Y(_6037_)
);

NAND2X1 _13022_ (
    .A(\u_ot.Yin12b [9]),
    .B(_6017_),
    .Y(_6038_)
);

OAI21X1 _13023_ (
    .A(_6037_),
    .B(_6017_),
    .C(_6038_),
    .Y(_5862_)
);

NAND2X1 _13024_ (
    .A(\u_ot.Yin12b [6]),
    .B(_6021_),
    .Y(_6039_)
);

OAI21X1 _13025_ (
    .A(_6035_),
    .B(_6021_),
    .C(_6039_),
    .Y(_5863_)
);

NAND2X1 _13026_ (
    .A(\u_ot.Yin12b [7]),
    .B(_6021_),
    .Y(_6040_)
);

OAI21X1 _13027_ (
    .A(_6037_),
    .B(_6021_),
    .C(_6040_),
    .Y(_5864_)
);

NAND2X1 _13028_ (
    .A(\u_ot.Yin12b [4]),
    .B(_6025_),
    .Y(_6041_)
);

OAI21X1 _13029_ (
    .A(_6035_),
    .B(_6025_),
    .C(_6041_),
    .Y(_5865_)
);

NAND2X1 _13030_ (
    .A(\u_ot.Yin12b [5]),
    .B(_6025_),
    .Y(_6042_)
);

OAI21X1 _13031_ (
    .A(_6037_),
    .B(_6025_),
    .C(_6042_),
    .Y(_5866_)
);

OAI21X1 _13032_ (
    .A(\u_ot.LoadCtl [0]),
    .B(_6006_),
    .C(\u_ot.Yin1 [0]),
    .Y(_6043_)
);

OAI21X1 _13033_ (
    .A(_6035_),
    .B(_6028_),
    .C(_6043_),
    .Y(_5867_)
);

OAI21X1 _13034_ (
    .A(\u_ot.LoadCtl [0]),
    .B(_6006_),
    .C(\u_ot.Yin1 [1]),
    .Y(_6044_)
);

OAI21X1 _13035_ (
    .A(_6037_),
    .B(_6028_),
    .C(_6044_),
    .Y(_5868_)
);

NAND2X1 _13036_ (
    .A(\u_ot.LoadCtl [0]),
    .B(\genblk1[6].u_ce.Y_ [0]),
    .Y(_6045_)
);

OAI21X1 _13037_ (
    .A(\u_ot.LoadCtl [0]),
    .B(_5896_),
    .C(_6045_),
    .Y(_5869_)
);

NAND2X1 _13038_ (
    .A(\u_ot.LoadCtl [0]),
    .B(\genblk1[6].u_ce.Y_ [1]),
    .Y(_6046_)
);

OAI21X1 _13039_ (
    .A(\u_ot.LoadCtl [0]),
    .B(_5895_),
    .C(_6046_),
    .Y(_5870_)
);

DFFPOSX1 _13040_ (
    .CLK(clk_bF$buf64),
    .D(\u_ot.Xin0 [0]),
    .Q(\u_ot.Xcalc [0])
);

DFFPOSX1 _13041_ (
    .CLK(clk_bF$buf63),
    .D(_5845_[1]),
    .Q(\u_ot.Xcalc [1])
);

DFFPOSX1 _13042_ (
    .CLK(clk_bF$buf62),
    .D(_5845_[2]),
    .Q(\u_ot.Xcalc [2])
);

DFFPOSX1 _13043_ (
    .CLK(clk_bF$buf61),
    .D(_5845_[3]),
    .Q(\u_ot.Xcalc [3])
);

DFFPOSX1 _13044_ (
    .CLK(clk_bF$buf60),
    .D(_5845_[4]),
    .Q(\u_ot.Xcalc [4])
);

DFFPOSX1 _13045_ (
    .CLK(clk_bF$buf59),
    .D(_5845_[5]),
    .Q(\u_ot.Xcalc [5])
);

DFFPOSX1 _13046_ (
    .CLK(clk_bF$buf58),
    .D(_5845_[6]),
    .Q(\u_ot.Xcalc [6])
);

DFFPOSX1 _13047_ (
    .CLK(clk_bF$buf57),
    .D(_5845_[7]),
    .Q(\u_ot.Xcalc [7])
);

DFFPOSX1 _13048_ (
    .CLK(clk_bF$buf56),
    .D(_5845_[8]),
    .Q(\u_ot.Xcalc [8])
);

DFFPOSX1 _13049_ (
    .CLK(clk_bF$buf55),
    .D(_5845_[9]),
    .Q(\u_ot.Xcalc [9])
);

DFFPOSX1 _13050_ (
    .CLK(clk_bF$buf54),
    .D(_5845_[10]),
    .Q(\u_ot.Xcalc [10])
);

DFFPOSX1 _13051_ (
    .CLK(clk_bF$buf53),
    .D(_5845_[11]),
    .Q(\u_ot.Xcalc [11])
);

DFFPOSX1 _13052_ (
    .CLK(clk_bF$buf52),
    .D(\u_ot.Yin0 [0]),
    .Q(\u_ot.Ycalc [0])
);

DFFPOSX1 _13053_ (
    .CLK(clk_bF$buf51),
    .D(_5846_[1]),
    .Q(\u_ot.Ycalc [1])
);

DFFPOSX1 _13054_ (
    .CLK(clk_bF$buf50),
    .D(_5846_[2]),
    .Q(\u_ot.Ycalc [2])
);

DFFPOSX1 _13055_ (
    .CLK(clk_bF$buf49),
    .D(_5846_[3]),
    .Q(\u_ot.Ycalc [3])
);

DFFPOSX1 _13056_ (
    .CLK(clk_bF$buf48),
    .D(_5846_[4]),
    .Q(\u_ot.Ycalc [4])
);

DFFPOSX1 _13057_ (
    .CLK(clk_bF$buf47),
    .D(_5846_[5]),
    .Q(\u_ot.Ycalc [5])
);

DFFPOSX1 _13058_ (
    .CLK(clk_bF$buf46),
    .D(_5846_[6]),
    .Q(\u_ot.Ycalc [6])
);

DFFPOSX1 _13059_ (
    .CLK(clk_bF$buf45),
    .D(_5846_[7]),
    .Q(\u_ot.Ycalc [7])
);

DFFPOSX1 _13060_ (
    .CLK(clk_bF$buf44),
    .D(_5846_[8]),
    .Q(\u_ot.Ycalc [8])
);

DFFPOSX1 _13061_ (
    .CLK(clk_bF$buf43),
    .D(_5846_[9]),
    .Q(\u_ot.Ycalc [9])
);

DFFPOSX1 _13062_ (
    .CLK(clk_bF$buf42),
    .D(_5846_[10]),
    .Q(\u_ot.Ycalc [10])
);

DFFPOSX1 _13063_ (
    .CLK(clk_bF$buf41),
    .D(_5846_[11]),
    .Q(\u_ot.Ycalc [11])
);

DFFPOSX1 _13064_ (
    .CLK(clk_bF$buf40),
    .D(_5847_),
    .Q(\u_ot.Xin12b [10])
);

DFFPOSX1 _13065_ (
    .CLK(clk_bF$buf39),
    .D(_5848_),
    .Q(\u_ot.Xin12b [11])
);

DFFPOSX1 _13066_ (
    .CLK(clk_bF$buf38),
    .D(_5849_),
    .Q(\u_ot.Xin12b [8])
);

DFFPOSX1 _13067_ (
    .CLK(clk_bF$buf37),
    .D(_5850_),
    .Q(\u_ot.Xin12b [9])
);

DFFPOSX1 _13068_ (
    .CLK(clk_bF$buf36),
    .D(_5851_),
    .Q(\u_ot.Xin12b [6])
);

DFFPOSX1 _13069_ (
    .CLK(clk_bF$buf35),
    .D(_5852_),
    .Q(\u_ot.Xin12b [7])
);

DFFPOSX1 _13070_ (
    .CLK(clk_bF$buf34),
    .D(_5853_),
    .Q(\u_ot.Xin12b [4])
);

DFFPOSX1 _13071_ (
    .CLK(clk_bF$buf33),
    .D(_5854_),
    .Q(\u_ot.Xin12b [5])
);

DFFPOSX1 _13072_ (
    .CLK(clk_bF$buf32),
    .D(_5855_),
    .Q(\u_ot.Xin1 [0])
);

DFFPOSX1 _13073_ (
    .CLK(clk_bF$buf31),
    .D(_5856_),
    .Q(\u_ot.Xin1 [1])
);

DFFPOSX1 _13074_ (
    .CLK(clk_bF$buf30),
    .D(_5857_),
    .Q(\u_ot.Xin0 [0])
);

DFFPOSX1 _13075_ (
    .CLK(clk_bF$buf29),
    .D(_5858_),
    .Q(\u_ot.Xin0 [1])
);

DFFPOSX1 _13076_ (
    .CLK(clk_bF$buf28),
    .D(_5859_),
    .Q(\u_ot.Yin12b [10])
);

DFFPOSX1 _13077_ (
    .CLK(clk_bF$buf27),
    .D(_5860_),
    .Q(\u_ot.Yin12b [11])
);

DFFPOSX1 _13078_ (
    .CLK(clk_bF$buf26),
    .D(_5861_),
    .Q(\u_ot.Yin12b [8])
);

DFFPOSX1 _13079_ (
    .CLK(clk_bF$buf25),
    .D(_5862_),
    .Q(\u_ot.Yin12b [9])
);

DFFPOSX1 _13080_ (
    .CLK(clk_bF$buf24),
    .D(_5863_),
    .Q(\u_ot.Yin12b [6])
);

DFFPOSX1 _13081_ (
    .CLK(clk_bF$buf23),
    .D(_5864_),
    .Q(\u_ot.Yin12b [7])
);

DFFPOSX1 _13082_ (
    .CLK(clk_bF$buf22),
    .D(_5865_),
    .Q(\u_ot.Yin12b [4])
);

DFFPOSX1 _13083_ (
    .CLK(clk_bF$buf21),
    .D(_5866_),
    .Q(\u_ot.Yin12b [5])
);

DFFPOSX1 _13084_ (
    .CLK(clk_bF$buf20),
    .D(_5867_),
    .Q(\u_ot.Yin1 [0])
);

DFFPOSX1 _13085_ (
    .CLK(clk_bF$buf19),
    .D(_5868_),
    .Q(\u_ot.Yin1 [1])
);

DFFPOSX1 _13086_ (
    .CLK(clk_bF$buf18),
    .D(\genblk1[6].u_ce.ISout ),
    .Q(\u_ot.ISpipe [0])
);

DFFPOSX1 _13087_ (
    .CLK(clk_bF$buf17),
    .D(\u_ot.ISpipe [0]),
    .Q(\u_ot.ISpipe [1])
);

DFFPOSX1 _13088_ (
    .CLK(clk_bF$buf16),
    .D(\u_ot.ISpipe [1]),
    .Q(\u_ot.ISpipe [2])
);

DFFPOSX1 _13089_ (
    .CLK(clk_bF$buf15),
    .D(\u_ot.ISpipe [2]),
    .Q(\u_ot.ISpipe [3])
);

DFFPOSX1 _13090_ (
    .CLK(clk_bF$buf14),
    .D(\u_ot.ISpipe [3]),
    .Q(\u_ot.ISpipe [4])
);

DFFPOSX1 _13091_ (
    .CLK(clk_bF$buf13),
    .D(\u_ot.ISpipe [4]),
    .Q(\u_ot.ISpipe [5])
);

DFFPOSX1 _13092_ (
    .CLK(clk_bF$buf12),
    .D(\u_ot.ISpipe [5]),
    .Q(\u_ot.ISout )
);

DFFPOSX1 _13093_ (
    .CLK(clk_bF$buf11),
    .D(\genblk1[6].u_ce.Vld ),
    .Q(\u_ot.LoadCtl [0])
);

DFFPOSX1 _13094_ (
    .CLK(clk_bF$buf10),
    .D(\u_ot.LoadCtl [0]),
    .Q(\u_ot.LoadCtl [1])
);

DFFPOSX1 _13095_ (
    .CLK(clk_bF$buf9),
    .D(\u_ot.LoadCtl [1]),
    .Q(\u_ot.LoadCtl [2])
);

DFFPOSX1 _13096_ (
    .CLK(clk_bF$buf8),
    .D(\u_ot.LoadCtl [2]),
    .Q(\u_ot.LoadCtl [3])
);

DFFPOSX1 _13097_ (
    .CLK(clk_bF$buf7),
    .D(\u_ot.LoadCtl [3]),
    .Q(\u_ot.LoadCtl [4])
);

DFFPOSX1 _13098_ (
    .CLK(clk_bF$buf6),
    .D(\u_ot.LoadCtl [4]),
    .Q(\u_ot.LoadCtl [5])
);

DFFPOSX1 _13099_ (
    .CLK(clk_bF$buf5),
    .D(\u_ot.LoadCtl [5]),
    .Q(\u_ot.LoadCtl [6])
);

DFFPOSX1 _13100_ (
    .CLK(clk_bF$buf4),
    .D(_5869_),
    .Q(\u_ot.Yin0 [0])
);

DFFPOSX1 _13101_ (
    .CLK(clk_bF$buf3),
    .D(_5870_),
    .Q(\u_ot.Yin0 [1])
);

INVX1 _13102_ (
    .A(\u_pa.Atmp [4]),
    .Y(_6086_)
);

INVX1 _13103_ (
    .A(\u_pa.RdyCtl [2]),
    .Y(_6087_)
);

INVX1 _13104_ (
    .A(\u_pa.Atmp [6]),
    .Y(_6088_)
);

INVX1 _13105_ (
    .A(\u_pa.RdyCtl [3]),
    .Y(_6089_)
);

INVX1 _13106_ (
    .A(\u_pa.Atmp [8]),
    .Y(_6090_)
);

INVX1 _13107_ (
    .A(\u_pa.RdyCtl [4]),
    .Y(_6091_)
);

NAND2X1 _13108_ (
    .A(\u_pa.Atmp [11]),
    .B(_6091_),
    .Y(_6092_)
);

OAI21X1 _13109_ (
    .A(_6090_),
    .B(_6091_),
    .C(_6092_),
    .Y(_6093_)
);

NAND2X1 _13110_ (
    .A(_6089_),
    .B(_6093_),
    .Y(_6094_)
);

OAI21X1 _13111_ (
    .A(_6088_),
    .B(_6089_),
    .C(_6094_),
    .Y(_6095_)
);

NAND2X1 _13112_ (
    .A(_6087_),
    .B(_6095_),
    .Y(_6096_)
);

OAI21X1 _13113_ (
    .A(_6086_),
    .B(_6087_),
    .C(_6096_),
    .Y(_6097_)
);

INVX1 _13114_ (
    .A(\u_pa.Atmp [2]),
    .Y(_6098_)
);

NAND2X1 _13115_ (
    .A(\u_pa.RdyCtl [1]),
    .B(_6098_),
    .Y(_6099_)
);

OAI21X1 _13116_ (
    .A(\u_pa.RdyCtl [1]),
    .B(_6097_),
    .C(_6099_),
    .Y(_6100_)
);

NAND2X1 _13117_ (
    .A(\u_pa.Atmp [0]),
    .B(\u_pa.RdyCtl [0]),
    .Y(_6101_)
);

OAI21X1 _13118_ (
    .A(\u_pa.RdyCtl [0]),
    .B(_6100_),
    .C(_6101_),
    .Y(\a[0] [0])
);

INVX1 _13119_ (
    .A(\u_pa.Atmp [5]),
    .Y(_6102_)
);

INVX1 _13120_ (
    .A(\u_pa.Atmp [9]),
    .Y(_6103_)
);

OAI21X1 _13121_ (
    .A(_6091_),
    .B(_6103_),
    .C(_6092_),
    .Y(_6104_)
);

INVX1 _13122_ (
    .A(\u_pa.Atmp [7]),
    .Y(_6105_)
);

AOI21X1 _13123_ (
    .A(_6105_),
    .B(\u_pa.RdyCtl [3]),
    .C(\u_pa.RdyCtl [2]),
    .Y(_6106_)
);

OAI21X1 _13124_ (
    .A(\u_pa.RdyCtl [3]),
    .B(_6104_),
    .C(_6106_),
    .Y(_6107_)
);

OAI21X1 _13125_ (
    .A(_6087_),
    .B(_6102_),
    .C(_6107_),
    .Y(_6108_)
);

INVX1 _13126_ (
    .A(\u_pa.Atmp [3]),
    .Y(_6109_)
);

NAND2X1 _13127_ (
    .A(\u_pa.RdyCtl [1]),
    .B(_6109_),
    .Y(_6110_)
);

OAI21X1 _13128_ (
    .A(\u_pa.RdyCtl [1]),
    .B(_6108_),
    .C(_6110_),
    .Y(_6111_)
);

NAND2X1 _13129_ (
    .A(\u_pa.RdyCtl [0]),
    .B(\u_pa.Atmp [1]),
    .Y(_6112_)
);

OAI21X1 _13130_ (
    .A(\u_pa.RdyCtl [0]),
    .B(_6111_),
    .C(_6112_),
    .Y(\a[0] [1])
);

INVX2 _13131_ (
    .A(\genblk1[0].u_ce.Rdy ),
    .Y(_6113_)
);

NAND2X1 _13132_ (
    .A(En),
    .B(_6113_),
    .Y(_6047_)
);

AND2X2 _13133_ (
    .A(\u_pa.RdyCtl [0]),
    .B(En),
    .Y(_6048_)
);

AND2X2 _13134_ (
    .A(\u_pa.RdyCtl [1]),
    .B(En),
    .Y(_6049_)
);

INVX2 _13135_ (
    .A(En),
    .Y(_6114_)
);

NOR2X1 _13136_ (
    .A(_6087_),
    .B(_6114_),
    .Y(_6050_)
);

NOR2X1 _13137_ (
    .A(_6089_),
    .B(_6114_),
    .Y(_6051_)
);

NOR2X1 _13138_ (
    .A(_6091_),
    .B(_6114_),
    .Y(_6052_)
);

AND2X2 _13139_ (
    .A(En),
    .B(\u_pa.RdyCtl [5]),
    .Y(_6053_)
);

NAND2X1 _13140_ (
    .A(\u_pa.acc_reg [18]),
    .B(\u_pa.acc_reg [19]),
    .Y(_6115_)
);

INVX1 _13141_ (
    .A(\u_pa.acc_reg [18]),
    .Y(_6116_)
);

INVX1 _13142_ (
    .A(\u_pa.acc_reg [19]),
    .Y(_6117_)
);

NAND2X1 _13143_ (
    .A(_6116_),
    .B(_6117_),
    .Y(_6118_)
);

NAND2X1 _13144_ (
    .A(_6115_),
    .B(_6118_),
    .Y(_6119_)
);

OAI21X1 _13145_ (
    .A(\genblk1[0].u_ce.ISin ),
    .B(\genblk1[0].u_ce.Rdy ),
    .C(En),
    .Y(_6120_)
);

AOI21X1 _13146_ (
    .A(_6119_),
    .B(\genblk1[0].u_ce.Rdy ),
    .C(_6120_),
    .Y(_6054_)
);

NAND2X1 _13147_ (
    .A(FCW[0]),
    .B(\u_pa.acc_reg [0]),
    .Y(_6121_)
);

INVX1 _13148_ (
    .A(_6121_),
    .Y(_6122_)
);

INVX1 _13149_ (
    .A(FCW[0]),
    .Y(_6123_)
);

NOR2X1 _13150_ (
    .A(_6123_),
    .B(_6113_),
    .Y(_6124_)
);

OAI21X1 _13151_ (
    .A(\u_pa.acc_reg [0]),
    .B(_6124_),
    .C(En),
    .Y(_6125_)
);

AOI21X1 _13152_ (
    .A(\genblk1[0].u_ce.Rdy ),
    .B(_6122_),
    .C(_6125_),
    .Y(_6055_)
);

INVX1 _13153_ (
    .A(\u_pa.acc_reg [1]),
    .Y(_6126_)
);

NAND2X1 _13154_ (
    .A(FCW[1]),
    .B(\u_pa.acc_reg [1]),
    .Y(_6127_)
);

INVX1 _13155_ (
    .A(_6127_),
    .Y(_6128_)
);

NOR2X1 _13156_ (
    .A(FCW[1]),
    .B(\u_pa.acc_reg [1]),
    .Y(_6129_)
);

OR2X2 _13157_ (
    .A(_6128_),
    .B(_6129_),
    .Y(_6130_)
);

INVX1 _13158_ (
    .A(_6130_),
    .Y(_6131_)
);

NOR2X1 _13159_ (
    .A(_6113_),
    .B(_6114_),
    .Y(_6132_)
);

INVX4 _13160_ (
    .A(_6132_),
    .Y(_6133_)
);

AOI21X1 _13161_ (
    .A(_6131_),
    .B(_6122_),
    .C(_6133__bF$buf3),
    .Y(_6134_)
);

OAI21X1 _13162_ (
    .A(_6122_),
    .B(_6131_),
    .C(_6134_),
    .Y(_6135_)
);

OAI21X1 _13163_ (
    .A(_6126_),
    .B(_6047__bF$buf3),
    .C(_6135_),
    .Y(_6056_)
);

OAI21X1 _13164_ (
    .A(_6121_),
    .B(_6129_),
    .C(_6127_),
    .Y(_6136_)
);

AND2X2 _13165_ (
    .A(FCW[2]),
    .B(\u_pa.acc_reg [2]),
    .Y(_6137_)
);

NOR2X1 _13166_ (
    .A(FCW[2]),
    .B(\u_pa.acc_reg [2]),
    .Y(_6138_)
);

NOR2X1 _13167_ (
    .A(_6138_),
    .B(_6137_),
    .Y(_6139_)
);

NOR2X1 _13168_ (
    .A(_6136_),
    .B(_6139_),
    .Y(_6140_)
);

AND2X2 _13169_ (
    .A(_6139_),
    .B(_6136_),
    .Y(_6141_)
);

OR2X2 _13170_ (
    .A(_6141_),
    .B(_6140_),
    .Y(_6142_)
);

OAI21X1 _13171_ (
    .A(\u_pa.acc_reg [2]),
    .B(\genblk1[0].u_ce.Rdy ),
    .C(En),
    .Y(_6143_)
);

AOI21X1 _13172_ (
    .A(_6142_),
    .B(\genblk1[0].u_ce.Rdy ),
    .C(_6143_),
    .Y(_6057_)
);

OAI21X1 _13173_ (
    .A(\u_pa.acc_reg [3]),
    .B(\genblk1[0].u_ce.Rdy ),
    .C(En),
    .Y(_6144_)
);

AND2X2 _13174_ (
    .A(FCW[3]),
    .B(\u_pa.acc_reg [3]),
    .Y(_6145_)
);

NOR2X1 _13175_ (
    .A(FCW[3]),
    .B(\u_pa.acc_reg [3]),
    .Y(_6146_)
);

NOR2X1 _13176_ (
    .A(_6146_),
    .B(_6145_),
    .Y(_6147_)
);

OAI21X1 _13177_ (
    .A(_6137_),
    .B(_6141_),
    .C(_6147_),
    .Y(_6148_)
);

NOR2X1 _13178_ (
    .A(_6137_),
    .B(_6141_),
    .Y(_6149_)
);

OAI21X1 _13179_ (
    .A(_6145_),
    .B(_6146_),
    .C(_6149_),
    .Y(_6150_)
);

NAND2X1 _13180_ (
    .A(_6148_),
    .B(_6150_),
    .Y(_6151_)
);

AOI21X1 _13181_ (
    .A(_6151_),
    .B(\genblk1[0].u_ce.Rdy ),
    .C(_6144_),
    .Y(_6058_)
);

INVX1 _13182_ (
    .A(\u_pa.acc_reg [4]),
    .Y(_6152_)
);

NAND3X1 _13183_ (
    .A(_6136_),
    .B(_6139_),
    .C(_6147_),
    .Y(_6153_)
);

INVX1 _13184_ (
    .A(_6146_),
    .Y(_6154_)
);

AOI21X1 _13185_ (
    .A(_6154_),
    .B(_6137_),
    .C(_6145_),
    .Y(_6155_)
);

NAND2X1 _13186_ (
    .A(_6155_),
    .B(_6153_),
    .Y(_6156_)
);

AND2X2 _13187_ (
    .A(FCW[4]),
    .B(\u_pa.acc_reg [4]),
    .Y(_6157_)
);

NOR2X1 _13188_ (
    .A(FCW[4]),
    .B(\u_pa.acc_reg [4]),
    .Y(_6158_)
);

NOR2X1 _13189_ (
    .A(_6158_),
    .B(_6157_),
    .Y(_6159_)
);

AND2X2 _13190_ (
    .A(_6156_),
    .B(_6159_),
    .Y(_6160_)
);

NOR2X1 _13191_ (
    .A(_6133__bF$buf2),
    .B(_6160_),
    .Y(_6161_)
);

OAI21X1 _13192_ (
    .A(_6156_),
    .B(_6159_),
    .C(_6161_),
    .Y(_6162_)
);

OAI21X1 _13193_ (
    .A(_6152_),
    .B(_6047__bF$buf2),
    .C(_6162_),
    .Y(_6059_)
);

OAI21X1 _13194_ (
    .A(\u_pa.acc_reg [5]),
    .B(\genblk1[0].u_ce.Rdy ),
    .C(En),
    .Y(_6163_)
);

NOR2X1 _13195_ (
    .A(_6157_),
    .B(_6160_),
    .Y(_6164_)
);

AND2X2 _13196_ (
    .A(FCW[5]),
    .B(\u_pa.acc_reg [5]),
    .Y(_6165_)
);

NOR2X1 _13197_ (
    .A(FCW[5]),
    .B(\u_pa.acc_reg [5]),
    .Y(_6166_)
);

OAI21X1 _13198_ (
    .A(_6165_),
    .B(_6166_),
    .C(_6164_),
    .Y(_6167_)
);

NOR2X1 _13199_ (
    .A(_6166_),
    .B(_6165_),
    .Y(_6168_)
);

OAI21X1 _13200_ (
    .A(_6157_),
    .B(_6160_),
    .C(_6168_),
    .Y(_6169_)
);

NAND2X1 _13201_ (
    .A(_6169_),
    .B(_6167_),
    .Y(_6170_)
);

AOI21X1 _13202_ (
    .A(_6170_),
    .B(\genblk1[0].u_ce.Rdy ),
    .C(_6163_),
    .Y(_6060_)
);

INVX1 _13203_ (
    .A(\u_pa.acc_reg [6]),
    .Y(_6171_)
);

INVX1 _13204_ (
    .A(_6157_),
    .Y(_6172_)
);

INVX1 _13205_ (
    .A(_6165_),
    .Y(_6173_)
);

OAI21X1 _13206_ (
    .A(_6166_),
    .B(_6172_),
    .C(_6173_),
    .Y(_6174_)
);

AND2X2 _13207_ (
    .A(_6159_),
    .B(_6168_),
    .Y(_6175_)
);

AOI21X1 _13208_ (
    .A(_6156_),
    .B(_6175_),
    .C(_6174_),
    .Y(_6176_)
);

NAND2X1 _13209_ (
    .A(FCW[6]),
    .B(\u_pa.acc_reg [6]),
    .Y(_6177_)
);

OR2X2 _13210_ (
    .A(FCW[6]),
    .B(\u_pa.acc_reg [6]),
    .Y(_6178_)
);

NAND2X1 _13211_ (
    .A(_6177_),
    .B(_6178_),
    .Y(_6179_)
);

NAND2X1 _13212_ (
    .A(_6179_),
    .B(_6176_),
    .Y(_6180_)
);

OR2X2 _13213_ (
    .A(_6176_),
    .B(_6179_),
    .Y(_6181_)
);

NAND3X1 _13214_ (
    .A(_6132_),
    .B(_6180_),
    .C(_6181_),
    .Y(_6182_)
);

OAI21X1 _13215_ (
    .A(_6171_),
    .B(_6047__bF$buf1),
    .C(_6182_),
    .Y(_6061_)
);

OAI21X1 _13216_ (
    .A(\u_pa.acc_reg [7]),
    .B(\genblk1[0].u_ce.Rdy ),
    .C(En),
    .Y(_6183_)
);

AND2X2 _13217_ (
    .A(_6181_),
    .B(_6177_),
    .Y(_6184_)
);

AND2X2 _13218_ (
    .A(FCW[7]),
    .B(\u_pa.acc_reg [7]),
    .Y(_6185_)
);

NOR2X1 _13219_ (
    .A(FCW[7]),
    .B(\u_pa.acc_reg [7]),
    .Y(_6186_)
);

NOR2X1 _13220_ (
    .A(_6186_),
    .B(_6185_),
    .Y(_6187_)
);

OR2X2 _13221_ (
    .A(_6184_),
    .B(_6187_),
    .Y(_6188_)
);

AOI21X1 _13222_ (
    .A(_6184_),
    .B(_6187_),
    .C(_6113_),
    .Y(_6189_)
);

AOI21X1 _13223_ (
    .A(_6188_),
    .B(_6189_),
    .C(_6183_),
    .Y(_6062_)
);

INVX1 _13224_ (
    .A(\u_pa.acc_reg [8]),
    .Y(_6190_)
);

NAND2X1 _13225_ (
    .A(_6159_),
    .B(_6168_),
    .Y(_6191_)
);

NAND3X1 _13226_ (
    .A(_6177_),
    .B(_6178_),
    .C(_6187_),
    .Y(_6192_)
);

NOR2X1 _13227_ (
    .A(_6191_),
    .B(_6192_),
    .Y(_6193_)
);

INVX1 _13228_ (
    .A(_6166_),
    .Y(_6194_)
);

AOI21X1 _13229_ (
    .A(_6194_),
    .B(_6157_),
    .C(_6165_),
    .Y(_6195_)
);

NAND2X1 _13230_ (
    .A(FCW[7]),
    .B(\u_pa.acc_reg [7]),
    .Y(_6196_)
);

OAI21X1 _13231_ (
    .A(_6177_),
    .B(_6186_),
    .C(_6196_),
    .Y(_6197_)
);

INVX1 _13232_ (
    .A(_6197_),
    .Y(_6198_)
);

OAI21X1 _13233_ (
    .A(_6195_),
    .B(_6192_),
    .C(_6198_),
    .Y(_6199_)
);

AOI21X1 _13234_ (
    .A(_6193_),
    .B(_6156_),
    .C(_6199_),
    .Y(_6200_)
);

NAND2X1 _13235_ (
    .A(FCW[8]),
    .B(\u_pa.acc_reg [8]),
    .Y(_6201_)
);

OR2X2 _13236_ (
    .A(FCW[8]),
    .B(\u_pa.acc_reg [8]),
    .Y(_6202_)
);

NAND2X1 _13237_ (
    .A(_6201_),
    .B(_6202_),
    .Y(_6203_)
);

AND2X2 _13238_ (
    .A(_6200_),
    .B(_6203_),
    .Y(_6204_)
);

OAI21X1 _13239_ (
    .A(_6203_),
    .B(_6200_),
    .C(_6132_),
    .Y(_6205_)
);

OAI22X1 _13240_ (
    .A(_6190_),
    .B(_6047__bF$buf0),
    .C(_6205_),
    .D(_6204_),
    .Y(_6063_)
);

OAI21X1 _13241_ (
    .A(\u_pa.acc_reg [9]),
    .B(\genblk1[0].u_ce.Rdy ),
    .C(En),
    .Y(_6206_)
);

OAI21X1 _13242_ (
    .A(_6203_),
    .B(_6200_),
    .C(_6201_),
    .Y(_6207_)
);

NAND2X1 _13243_ (
    .A(FCW[9]),
    .B(\u_pa.acc_reg [9]),
    .Y(_6208_)
);

INVX1 _13244_ (
    .A(FCW[9]),
    .Y(_6209_)
);

INVX1 _13245_ (
    .A(\u_pa.acc_reg [9]),
    .Y(_6210_)
);

NAND2X1 _13246_ (
    .A(_6209_),
    .B(_6210_),
    .Y(_6211_)
);

NAND2X1 _13247_ (
    .A(_6208_),
    .B(_6211_),
    .Y(_6212_)
);

NAND2X1 _13248_ (
    .A(_6212_),
    .B(_6207_),
    .Y(_6213_)
);

NOR2X1 _13249_ (
    .A(_6212_),
    .B(_6207_),
    .Y(_6214_)
);

NOR2X1 _13250_ (
    .A(_6113_),
    .B(_6214_),
    .Y(_6215_)
);

AOI21X1 _13251_ (
    .A(_6215_),
    .B(_6213_),
    .C(_6206_),
    .Y(_6064_)
);

INVX1 _13252_ (
    .A(\u_pa.acc_reg [10]),
    .Y(_6216_)
);

AND2X2 _13253_ (
    .A(_6153_),
    .B(_6155_),
    .Y(_6217_)
);

OR2X2 _13254_ (
    .A(FCW[7]),
    .B(\u_pa.acc_reg [7]),
    .Y(_6218_)
);

NAND2X1 _13255_ (
    .A(_6196_),
    .B(_6218_),
    .Y(_6219_)
);

NOR2X1 _13256_ (
    .A(_6219_),
    .B(_6179_),
    .Y(_6220_)
);

NAND2X1 _13257_ (
    .A(_6220_),
    .B(_6175_),
    .Y(_6221_)
);

AOI21X1 _13258_ (
    .A(_6220_),
    .B(_6174_),
    .C(_6197_),
    .Y(_6222_)
);

OAI21X1 _13259_ (
    .A(_6221_),
    .B(_6217_),
    .C(_6222_),
    .Y(_6223_)
);

NOR2X1 _13260_ (
    .A(FCW[9]),
    .B(\u_pa.acc_reg [9]),
    .Y(_6224_)
);

OAI21X1 _13261_ (
    .A(_6201_),
    .B(_6224_),
    .C(_6208_),
    .Y(_6225_)
);

NOR2X1 _13262_ (
    .A(_6203_),
    .B(_6212_),
    .Y(_6226_)
);

AOI21X1 _13263_ (
    .A(_6223_),
    .B(_6226_),
    .C(_6225_),
    .Y(_6227_)
);

INVX1 _13264_ (
    .A(_6227_),
    .Y(_6228_)
);

AND2X2 _13265_ (
    .A(FCW[10]),
    .B(\u_pa.acc_reg [10]),
    .Y(_6229_)
);

NOR2X1 _13266_ (
    .A(FCW[10]),
    .B(\u_pa.acc_reg [10]),
    .Y(_6230_)
);

NOR2X1 _13267_ (
    .A(_6230_),
    .B(_6229_),
    .Y(_6231_)
);

AOI21X1 _13268_ (
    .A(_6228_),
    .B(_6231_),
    .C(_6133__bF$buf1),
    .Y(_6232_)
);

OAI21X1 _13269_ (
    .A(_6228_),
    .B(_6231_),
    .C(_6232_),
    .Y(_6233_)
);

OAI21X1 _13270_ (
    .A(_6216_),
    .B(_6047__bF$buf3),
    .C(_6233_),
    .Y(_6065_)
);

INVX1 _13271_ (
    .A(\u_pa.acc_reg [11]),
    .Y(_6234_)
);

OAI21X1 _13272_ (
    .A(_6234_),
    .B(_6114_),
    .C(_6133__bF$buf0),
    .Y(_6235_)
);

INVX1 _13273_ (
    .A(_6229_),
    .Y(_6236_)
);

OAI21X1 _13274_ (
    .A(_6230_),
    .B(_6227_),
    .C(_6236_),
    .Y(_6237_)
);

AND2X2 _13275_ (
    .A(FCW[11]),
    .B(\u_pa.acc_reg [11]),
    .Y(_6238_)
);

NOR2X1 _13276_ (
    .A(FCW[11]),
    .B(\u_pa.acc_reg [11]),
    .Y(_6239_)
);

NOR2X1 _13277_ (
    .A(_6239_),
    .B(_6238_),
    .Y(_6240_)
);

INVX1 _13278_ (
    .A(_6240_),
    .Y(_6241_)
);

AOI21X1 _13279_ (
    .A(_6237_),
    .B(_6241_),
    .C(_6113_),
    .Y(_6242_)
);

OAI21X1 _13280_ (
    .A(_6237_),
    .B(_6241_),
    .C(_6242_),
    .Y(_6243_)
);

AND2X2 _13281_ (
    .A(_6243_),
    .B(_6235_),
    .Y(_6066_)
);

INVX1 _13282_ (
    .A(\u_pa.acc_reg [12]),
    .Y(_6244_)
);

NAND3X1 _13283_ (
    .A(_6231_),
    .B(_6240_),
    .C(_6226_),
    .Y(_6245_)
);

NAND3X1 _13284_ (
    .A(_6225_),
    .B(_6231_),
    .C(_6240_),
    .Y(_6246_)
);

INVX1 _13285_ (
    .A(_6239_),
    .Y(_6247_)
);

AOI21X1 _13286_ (
    .A(_6247_),
    .B(_6229_),
    .C(_6238_),
    .Y(_6248_)
);

AND2X2 _13287_ (
    .A(_6246_),
    .B(_6248_),
    .Y(_6249_)
);

OAI21X1 _13288_ (
    .A(_6245_),
    .B(_6200_),
    .C(_6249_),
    .Y(_6250_)
);

NAND2X1 _13289_ (
    .A(FCW[12]),
    .B(\u_pa.acc_reg [12]),
    .Y(_6251_)
);

OR2X2 _13290_ (
    .A(FCW[12]),
    .B(\u_pa.acc_reg [12]),
    .Y(_6252_)
);

NAND2X1 _13291_ (
    .A(_6251_),
    .B(_6252_),
    .Y(_6253_)
);

INVX1 _13292_ (
    .A(_6253_),
    .Y(_6254_)
);

NOR2X1 _13293_ (
    .A(_6254_),
    .B(_6250_),
    .Y(_6255_)
);

INVX1 _13294_ (
    .A(_6245_),
    .Y(_6256_)
);

NAND2X1 _13295_ (
    .A(_6248_),
    .B(_6246_),
    .Y(_6257_)
);

AOI21X1 _13296_ (
    .A(_6223_),
    .B(_6256_),
    .C(_6257_),
    .Y(_6258_)
);

OAI21X1 _13297_ (
    .A(_6253_),
    .B(_6258_),
    .C(_6132_),
    .Y(_6259_)
);

OAI22X1 _13298_ (
    .A(_6244_),
    .B(_6047__bF$buf2),
    .C(_6255_),
    .D(_6259_),
    .Y(_6067_)
);

INVX1 _13299_ (
    .A(\u_pa.acc_reg [13]),
    .Y(_6260_)
);

OAI21X1 _13300_ (
    .A(_6260_),
    .B(_6114_),
    .C(_6133__bF$buf3),
    .Y(_6261_)
);

OAI21X1 _13301_ (
    .A(_6253_),
    .B(_6258_),
    .C(_6251_),
    .Y(_6262_)
);

NAND2X1 _13302_ (
    .A(FCW[13]),
    .B(\u_pa.acc_reg [13]),
    .Y(_6263_)
);

OR2X2 _13303_ (
    .A(FCW[13]),
    .B(\u_pa.acc_reg [13]),
    .Y(_6264_)
);

NAND2X1 _13304_ (
    .A(_6263_),
    .B(_6264_),
    .Y(_6265_)
);

AOI21X1 _13305_ (
    .A(_6262_),
    .B(_6265_),
    .C(_6113_),
    .Y(_6266_)
);

OAI21X1 _13306_ (
    .A(_6262_),
    .B(_6265_),
    .C(_6266_),
    .Y(_6267_)
);

AND2X2 _13307_ (
    .A(_6267_),
    .B(_6261_),
    .Y(_6068_)
);

INVX1 _13308_ (
    .A(\u_pa.acc_reg [14]),
    .Y(_6268_)
);

NOR2X1 _13309_ (
    .A(_6253_),
    .B(_6265_),
    .Y(_6269_)
);

NOR2X1 _13310_ (
    .A(FCW[13]),
    .B(\u_pa.acc_reg [13]),
    .Y(_6270_)
);

OAI21X1 _13311_ (
    .A(_6251_),
    .B(_6270_),
    .C(_6263_),
    .Y(_6271_)
);

AOI21X1 _13312_ (
    .A(_6250_),
    .B(_6269_),
    .C(_6271_),
    .Y(_6272_)
);

AND2X2 _13313_ (
    .A(FCW[14]),
    .B(\u_pa.acc_reg [14]),
    .Y(_6273_)
);

NOR2X1 _13314_ (
    .A(FCW[14]),
    .B(\u_pa.acc_reg [14]),
    .Y(_6274_)
);

OAI21X1 _13315_ (
    .A(_6273_),
    .B(_6274_),
    .C(_6272_),
    .Y(_6275_)
);

OR2X2 _13316_ (
    .A(_6273_),
    .B(_6274_),
    .Y(_6276_)
);

OR2X2 _13317_ (
    .A(_6272_),
    .B(_6276_),
    .Y(_6277_)
);

NAND3X1 _13318_ (
    .A(_6132_),
    .B(_6275_),
    .C(_6277_),
    .Y(_6278_)
);

OAI21X1 _13319_ (
    .A(_6268_),
    .B(_6047__bF$buf1),
    .C(_6278_),
    .Y(_6069_)
);

OAI21X1 _13320_ (
    .A(\u_pa.acc_reg [15]),
    .B(\genblk1[0].u_ce.Rdy ),
    .C(En),
    .Y(_6279_)
);

NAND2X1 _13321_ (
    .A(FCW[14]),
    .B(\u_pa.acc_reg [14]),
    .Y(_6280_)
);

NAND2X1 _13322_ (
    .A(FCW[15]),
    .B(\u_pa.acc_reg [15]),
    .Y(_6281_)
);

INVX1 _13323_ (
    .A(_6281_),
    .Y(_6282_)
);

NOR2X1 _13324_ (
    .A(FCW[15]),
    .B(\u_pa.acc_reg [15]),
    .Y(_6283_)
);

NOR2X1 _13325_ (
    .A(_6283_),
    .B(_6282_),
    .Y(_6284_)
);

NAND3X1 _13326_ (
    .A(_6280_),
    .B(_6284_),
    .C(_6277_),
    .Y(_6285_)
);

OAI21X1 _13327_ (
    .A(_6276_),
    .B(_6272_),
    .C(_6280_),
    .Y(_6286_)
);

INVX1 _13328_ (
    .A(_6283_),
    .Y(_6287_)
);

NAND2X1 _13329_ (
    .A(_6281_),
    .B(_6287_),
    .Y(_6288_)
);

AOI21X1 _13330_ (
    .A(_6286_),
    .B(_6288_),
    .C(_6113_),
    .Y(_6289_)
);

AOI21X1 _13331_ (
    .A(_6285_),
    .B(_6289_),
    .C(_6279_),
    .Y(_6070_)
);

INVX1 _13332_ (
    .A(\u_pa.acc_reg [16]),
    .Y(_6290_)
);

NOR2X1 _13333_ (
    .A(_6276_),
    .B(_6288_),
    .Y(_6291_)
);

AND2X2 _13334_ (
    .A(_6291_),
    .B(_6269_),
    .Y(_6292_)
);

NAND2X1 _13335_ (
    .A(_6292_),
    .B(_6256_),
    .Y(_6293_)
);

NOR2X1 _13336_ (
    .A(_6274_),
    .B(_6273_),
    .Y(_6294_)
);

NAND3X1 _13337_ (
    .A(_6271_),
    .B(_6294_),
    .C(_6284_),
    .Y(_6295_)
);

AOI21X1 _13338_ (
    .A(_6287_),
    .B(_6273_),
    .C(_6282_),
    .Y(_6296_)
);

NAND2X1 _13339_ (
    .A(_6296_),
    .B(_6295_),
    .Y(_6297_)
);

AOI21X1 _13340_ (
    .A(_6292_),
    .B(_6257_),
    .C(_6297_),
    .Y(_6298_)
);

OAI21X1 _13341_ (
    .A(_6200_),
    .B(_6293_),
    .C(_6298_),
    .Y(_6299_)
);

AND2X2 _13342_ (
    .A(FCW[16]),
    .B(\u_pa.acc_reg [16]),
    .Y(_6300_)
);

NOR2X1 _13343_ (
    .A(FCW[16]),
    .B(\u_pa.acc_reg [16]),
    .Y(_6301_)
);

NOR2X1 _13344_ (
    .A(_6301_),
    .B(_6300_),
    .Y(_6302_)
);

NAND3X1 _13345_ (
    .A(_6294_),
    .B(_6284_),
    .C(_6269_),
    .Y(_6303_)
);

NOR2X1 _13346_ (
    .A(_6245_),
    .B(_6303_),
    .Y(_6304_)
);

AND2X2 _13347_ (
    .A(_6295_),
    .B(_6296_),
    .Y(_6305_)
);

OAI21X1 _13348_ (
    .A(_6303_),
    .B(_6249_),
    .C(_6305_),
    .Y(_6306_)
);

AOI21X1 _13349_ (
    .A(_6223_),
    .B(_6304_),
    .C(_6306_),
    .Y(_6307_)
);

INVX1 _13350_ (
    .A(_6302_),
    .Y(_6308_)
);

NOR2X1 _13351_ (
    .A(_6308_),
    .B(_6307_),
    .Y(_6309_)
);

NOR2X1 _13352_ (
    .A(_6133__bF$buf2),
    .B(_6309_),
    .Y(_6310_)
);

OAI21X1 _13353_ (
    .A(_6299_),
    .B(_6302_),
    .C(_6310_),
    .Y(_6311_)
);

OAI21X1 _13354_ (
    .A(_6290_),
    .B(_6047__bF$buf0),
    .C(_6311_),
    .Y(_6071_)
);

NAND2X1 _13355_ (
    .A(\u_pa.acc_reg [17]),
    .B(En),
    .Y(_6312_)
);

AND2X2 _13356_ (
    .A(FCW[17]),
    .B(\u_pa.acc_reg [17]),
    .Y(_6313_)
);

NOR2X1 _13357_ (
    .A(FCW[17]),
    .B(\u_pa.acc_reg [17]),
    .Y(_6314_)
);

NOR2X1 _13358_ (
    .A(_6314_),
    .B(_6313_),
    .Y(_6315_)
);

INVX1 _13359_ (
    .A(_6315_),
    .Y(_6316_)
);

OAI21X1 _13360_ (
    .A(_6300_),
    .B(_6309_),
    .C(_6316_),
    .Y(_6317_)
);

NOR2X1 _13361_ (
    .A(_6300_),
    .B(_6309_),
    .Y(_6318_)
);

AOI21X1 _13362_ (
    .A(_6318_),
    .B(_6315_),
    .C(_6113_),
    .Y(_6319_)
);

AOI22X1 _13363_ (
    .A(_6133__bF$buf1),
    .B(_6312_),
    .C(_6319_),
    .D(_6317_),
    .Y(_6072_)
);

NAND2X1 _13364_ (
    .A(_6302_),
    .B(_6315_),
    .Y(_6320_)
);

AOI21X1 _13365_ (
    .A(_6315_),
    .B(_6300_),
    .C(_6313_),
    .Y(_6321_)
);

OAI21X1 _13366_ (
    .A(_6320_),
    .B(_6307_),
    .C(_6321_),
    .Y(_6322_)
);

INVX1 _13367_ (
    .A(FCW[18]),
    .Y(_6323_)
);

NOR2X1 _13368_ (
    .A(_6116_),
    .B(_6323_),
    .Y(_6324_)
);

NOR2X1 _13369_ (
    .A(\u_pa.acc_reg [18]),
    .B(FCW[18]),
    .Y(_6325_)
);

NOR2X1 _13370_ (
    .A(_6325_),
    .B(_6324_),
    .Y(_6326_)
);

NOR2X1 _13371_ (
    .A(_6326_),
    .B(_6322_),
    .Y(_6327_)
);

INVX1 _13372_ (
    .A(_6320_),
    .Y(_6328_)
);

INVX1 _13373_ (
    .A(_6321_),
    .Y(_6329_)
);

AOI21X1 _13374_ (
    .A(_6299_),
    .B(_6328_),
    .C(_6329_),
    .Y(_6330_)
);

INVX1 _13375_ (
    .A(_6326_),
    .Y(_6331_)
);

OAI21X1 _13376_ (
    .A(_6331_),
    .B(_6330_),
    .C(_6132_),
    .Y(_6332_)
);

OAI22X1 _13377_ (
    .A(_6116_),
    .B(_6047__bF$buf3),
    .C(_6327_),
    .D(_6332_),
    .Y(_6073_)
);

NAND2X1 _13378_ (
    .A(\u_pa.acc_reg [19]),
    .B(En),
    .Y(_6333_)
);

INVX1 _13379_ (
    .A(_6324_),
    .Y(_6334_)
);

OAI21X1 _13380_ (
    .A(_6331_),
    .B(_6330_),
    .C(_6334_),
    .Y(_6335_)
);

NAND2X1 _13381_ (
    .A(\u_pa.acc_reg [19]),
    .B(FCW[19]),
    .Y(_6336_)
);

OR2X2 _13382_ (
    .A(\u_pa.acc_reg [19]),
    .B(FCW[19]),
    .Y(_6337_)
);

NAND2X1 _13383_ (
    .A(_6336_),
    .B(_6337_),
    .Y(_6338_)
);

NAND2X1 _13384_ (
    .A(_6338_),
    .B(_6335_),
    .Y(_6339_)
);

AOI21X1 _13385_ (
    .A(_6322_),
    .B(_6326_),
    .C(_6324_),
    .Y(_6340_)
);

INVX1 _13386_ (
    .A(_6338_),
    .Y(_6341_)
);

AOI21X1 _13387_ (
    .A(_6340_),
    .B(_6341_),
    .C(_6113_),
    .Y(_6342_)
);

AOI22X1 _13388_ (
    .A(_6133__bF$buf0),
    .B(_6333_),
    .C(_6342_),
    .D(_6339_),
    .Y(_6074_)
);

INVX1 _13389_ (
    .A(\u_pa.Atmp [0]),
    .Y(_6343_)
);

OAI22X1 _13390_ (
    .A(_6343_),
    .B(_6047__bF$buf2),
    .C(_6190_),
    .D(_6133__bF$buf3),
    .Y(_6075_)
);

INVX1 _13391_ (
    .A(\u_pa.Atmp [1]),
    .Y(_6344_)
);

OAI22X1 _13392_ (
    .A(_6344_),
    .B(_6047__bF$buf1),
    .C(_6210_),
    .D(_6133__bF$buf2),
    .Y(_6076_)
);

OAI22X1 _13393_ (
    .A(_6098_),
    .B(_6047__bF$buf0),
    .C(_6216_),
    .D(_6133__bF$buf1),
    .Y(_6077_)
);

OAI22X1 _13394_ (
    .A(_6109_),
    .B(_6047__bF$buf3),
    .C(_6234_),
    .D(_6133__bF$buf0),
    .Y(_6078_)
);

OAI22X1 _13395_ (
    .A(_6086_),
    .B(_6047__bF$buf2),
    .C(_6244_),
    .D(_6133__bF$buf3),
    .Y(_6079_)
);

OAI22X1 _13396_ (
    .A(_6102_),
    .B(_6047__bF$buf1),
    .C(_6260_),
    .D(_6133__bF$buf2),
    .Y(_6080_)
);

OAI22X1 _13397_ (
    .A(_6088_),
    .B(_6047__bF$buf0),
    .C(_6268_),
    .D(_6133__bF$buf1),
    .Y(_6081_)
);

NAND2X1 _13398_ (
    .A(\u_pa.acc_reg [15]),
    .B(_6132_),
    .Y(_6345_)
);

OAI21X1 _13399_ (
    .A(_6105_),
    .B(_6047__bF$buf3),
    .C(_6345_),
    .Y(_6082_)
);

OAI22X1 _13400_ (
    .A(_6090_),
    .B(_6047__bF$buf2),
    .C(_6290_),
    .D(_6133__bF$buf0),
    .Y(_6083_)
);

NAND2X1 _13401_ (
    .A(\u_pa.acc_reg [17]),
    .B(_6132_),
    .Y(_6346_)
);

OAI21X1 _13402_ (
    .A(_6103_),
    .B(_6047__bF$buf1),
    .C(_6346_),
    .Y(_6084_)
);

INVX1 _13403_ (
    .A(\u_pa.Atmp [11]),
    .Y(_6347_)
);

OAI22X1 _13404_ (
    .A(_6347_),
    .B(_6047__bF$buf0),
    .C(_6116_),
    .D(_6133__bF$buf3),
    .Y(_6085_)
);

DFFPOSX1 _13405_ (
    .CLK(clk_bF$buf2),
    .D(_6047__bF$buf3),
    .Q(\u_pa.RdyCtl [0])
);

DFFPOSX1 _13406_ (
    .CLK(clk_bF$buf1),
    .D(_6048_),
    .Q(\u_pa.RdyCtl [1])
);

DFFPOSX1 _13407_ (
    .CLK(clk_bF$buf0),
    .D(_6049_),
    .Q(\u_pa.RdyCtl [2])
);

DFFPOSX1 _13408_ (
    .CLK(clk_bF$buf75),
    .D(_6050_),
    .Q(\u_pa.RdyCtl [3])
);

DFFPOSX1 _13409_ (
    .CLK(clk_bF$buf74),
    .D(_6051_),
    .Q(\u_pa.RdyCtl [4])
);

DFFPOSX1 _13410_ (
    .CLK(clk_bF$buf73),
    .D(_6052_),
    .Q(\u_pa.RdyCtl [5])
);

DFFPOSX1 _13411_ (
    .CLK(clk_bF$buf72),
    .D(_6053_),
    .Q(\genblk1[0].u_ce.Rdy )
);

DFFPOSX1 _13412_ (
    .CLK(clk_bF$buf71),
    .D(_6054_),
    .Q(\genblk1[0].u_ce.ISin )
);

DFFPOSX1 _13413_ (
    .CLK(clk_bF$buf70),
    .D(_6055_),
    .Q(\u_pa.acc_reg [0])
);

DFFPOSX1 _13414_ (
    .CLK(clk_bF$buf69),
    .D(_6056_),
    .Q(\u_pa.acc_reg [1])
);

DFFPOSX1 _13415_ (
    .CLK(clk_bF$buf68),
    .D(_6057_),
    .Q(\u_pa.acc_reg [2])
);

DFFPOSX1 _13416_ (
    .CLK(clk_bF$buf67),
    .D(_6058_),
    .Q(\u_pa.acc_reg [3])
);

DFFPOSX1 _13417_ (
    .CLK(clk_bF$buf66),
    .D(_6059_),
    .Q(\u_pa.acc_reg [4])
);

DFFPOSX1 _13418_ (
    .CLK(clk_bF$buf65),
    .D(_6060_),
    .Q(\u_pa.acc_reg [5])
);

DFFPOSX1 _13419_ (
    .CLK(clk_bF$buf64),
    .D(_6061_),
    .Q(\u_pa.acc_reg [6])
);

DFFPOSX1 _13420_ (
    .CLK(clk_bF$buf63),
    .D(_6062_),
    .Q(\u_pa.acc_reg [7])
);

DFFPOSX1 _13421_ (
    .CLK(clk_bF$buf62),
    .D(_6063_),
    .Q(\u_pa.acc_reg [8])
);

DFFPOSX1 _13422_ (
    .CLK(clk_bF$buf61),
    .D(_6064_),
    .Q(\u_pa.acc_reg [9])
);

DFFPOSX1 _13423_ (
    .CLK(clk_bF$buf60),
    .D(_6065_),
    .Q(\u_pa.acc_reg [10])
);

DFFPOSX1 _13424_ (
    .CLK(clk_bF$buf59),
    .D(_6066_),
    .Q(\u_pa.acc_reg [11])
);

DFFPOSX1 _13425_ (
    .CLK(clk_bF$buf58),
    .D(_6067_),
    .Q(\u_pa.acc_reg [12])
);

DFFPOSX1 _13426_ (
    .CLK(clk_bF$buf57),
    .D(_6068_),
    .Q(\u_pa.acc_reg [13])
);

DFFPOSX1 _13427_ (
    .CLK(clk_bF$buf56),
    .D(_6069_),
    .Q(\u_pa.acc_reg [14])
);

DFFPOSX1 _13428_ (
    .CLK(clk_bF$buf55),
    .D(_6070_),
    .Q(\u_pa.acc_reg [15])
);

DFFPOSX1 _13429_ (
    .CLK(clk_bF$buf54),
    .D(_6071_),
    .Q(\u_pa.acc_reg [16])
);

DFFPOSX1 _13430_ (
    .CLK(clk_bF$buf53),
    .D(_6072_),
    .Q(\u_pa.acc_reg [17])
);

DFFPOSX1 _13431_ (
    .CLK(clk_bF$buf52),
    .D(_6073_),
    .Q(\u_pa.acc_reg [18])
);

DFFPOSX1 _13432_ (
    .CLK(clk_bF$buf51),
    .D(_6074_),
    .Q(\u_pa.acc_reg [19])
);

DFFPOSX1 _13433_ (
    .CLK(clk_bF$buf50),
    .D(_6075_),
    .Q(\u_pa.Atmp [0])
);

DFFPOSX1 _13434_ (
    .CLK(clk_bF$buf49),
    .D(_6076_),
    .Q(\u_pa.Atmp [1])
);

DFFPOSX1 _13435_ (
    .CLK(clk_bF$buf48),
    .D(_6077_),
    .Q(\u_pa.Atmp [2])
);

DFFPOSX1 _13436_ (
    .CLK(clk_bF$buf47),
    .D(_6078_),
    .Q(\u_pa.Atmp [3])
);

DFFPOSX1 _13437_ (
    .CLK(clk_bF$buf46),
    .D(_6079_),
    .Q(\u_pa.Atmp [4])
);

DFFPOSX1 _13438_ (
    .CLK(clk_bF$buf45),
    .D(_6080_),
    .Q(\u_pa.Atmp [5])
);

DFFPOSX1 _13439_ (
    .CLK(clk_bF$buf44),
    .D(_6081_),
    .Q(\u_pa.Atmp [6])
);

DFFPOSX1 _13440_ (
    .CLK(clk_bF$buf43),
    .D(_6082_),
    .Q(\u_pa.Atmp [7])
);

DFFPOSX1 _13441_ (
    .CLK(clk_bF$buf42),
    .D(_6083_),
    .Q(\u_pa.Atmp [8])
);

DFFPOSX1 _13442_ (
    .CLK(clk_bF$buf41),
    .D(_6084_),
    .Q(\u_pa.Atmp [9])
);

DFFPOSX1 _13443_ (
    .CLK(clk_bF$buf40),
    .D(_6085_),
    .Q(\u_pa.Atmp [11])
);

BUFX2 _13444_ (
    .A(_6348_[0]),
    .Y(Dout[0])
);

BUFX2 _13445_ (
    .A(_6348_[1]),
    .Y(Dout[1])
);

BUFX2 _13446_ (
    .A(_6348_[10]),
    .Y(Dout[10])
);

BUFX2 _13447_ (
    .A(_6348_[11]),
    .Y(Dout[11])
);

BUFX2 _13448_ (
    .A(_6348_[2]),
    .Y(Dout[2])
);

BUFX2 _13449_ (
    .A(_6348_[3]),
    .Y(Dout[3])
);

BUFX2 _13450_ (
    .A(_6348_[4]),
    .Y(Dout[4])
);

BUFX2 _13451_ (
    .A(_6348_[5]),
    .Y(Dout[5])
);

BUFX2 _13452_ (
    .A(_6348_[6]),
    .Y(Dout[6])
);

BUFX2 _13453_ (
    .A(_6348_[7]),
    .Y(Dout[7])
);

BUFX2 _13454_ (
    .A(_6348_[8]),
    .Y(Dout[8])
);

BUFX2 _13455_ (
    .A(_6348_[9]),
    .Y(Dout[9])
);

BUFX2 _13456_ (
    .A(\u_ot.LoadCtl [6]),
    .Y(Vld)
);

NOR2X1 _6349_ (
    .A(\genblk1[0].u_ce.LoadCtl [3]),
    .B(\genblk1[0].u_ce.LoadCtl [2]),
    .Y(_92_)
);

INVX1 _6350_ (
    .A(\genblk1[0].u_ce.Acalc [10]),
    .Y(_93_)
);

NAND2X1 _6351_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(\genblk1[0].u_ce.Acalc [8]),
    .Y(_94_)
);

OAI21X1 _6352_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(_93_),
    .C(_94_),
    .Y(_95_)
);

INVX2 _6353_ (
    .A(\genblk1[0].u_ce.LoadCtl [2]),
    .Y(_96_)
);

INVX1 _6354_ (
    .A(\genblk1[0].u_ce.Acalc [4]),
    .Y(_97_)
);

INVX1 _6355_ (
    .A(\genblk1[0].u_ce.LoadCtl [3]),
    .Y(_98_)
);

NOR2X1 _6356_ (
    .A(\genblk1[0].u_ce.LoadCtl [2]),
    .B(_98_),
    .Y(_99_)
);

NAND2X1 _6357_ (
    .A(\genblk1[0].u_ce.Acalc [6]),
    .B(_99_),
    .Y(_100_)
);

OAI21X1 _6358_ (
    .A(_96_),
    .B(_97_),
    .C(_100_),
    .Y(_101_)
);

AOI21X1 _6359_ (
    .A(_92_),
    .B(_95_),
    .C(_101_),
    .Y(_102_)
);

NOR2X1 _6360_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[0].u_ce.LoadCtl [1]),
    .Y(_103_)
);

INVX4 _6361_ (
    .A(_103_),
    .Y(_104_)
);

INVX2 _6362_ (
    .A(\genblk1[0].u_ce.LoadCtl [1]),
    .Y(_105_)
);

NOR2X1 _6363_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_105_),
    .Y(_106_)
);

AOI22X1 _6364_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[0].u_ce.Acalc [0]),
    .C(_106_),
    .D(\genblk1[0].u_ce.Acalc [2]),
    .Y(_107_)
);

OAI21X1 _6365_ (
    .A(_104_),
    .B(_102_),
    .C(_107_),
    .Y(\a[1] [0])
);

INVX1 _6366_ (
    .A(\genblk1[0].u_ce.Acalc [11]),
    .Y(_108_)
);

NAND2X1 _6367_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(\genblk1[0].u_ce.Acalc [9]),
    .Y(_109_)
);

OAI21X1 _6368_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(_108_),
    .C(_109_),
    .Y(_110_)
);

INVX1 _6369_ (
    .A(\genblk1[0].u_ce.Acalc [7]),
    .Y(_111_)
);

INVX4 _6370_ (
    .A(_99_),
    .Y(_112_)
);

NAND2X1 _6371_ (
    .A(\genblk1[0].u_ce.LoadCtl [2]),
    .B(\genblk1[0].u_ce.Acalc [5]),
    .Y(_113_)
);

OAI21X1 _6372_ (
    .A(_111_),
    .B(_112_),
    .C(_113_),
    .Y(_114_)
);

AOI21X1 _6373_ (
    .A(_92_),
    .B(_110_),
    .C(_114_),
    .Y(_115_)
);

AOI22X1 _6374_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[0].u_ce.Acalc [1]),
    .C(_106_),
    .D(\genblk1[0].u_ce.Acalc [3]),
    .Y(_116_)
);

OAI21X1 _6375_ (
    .A(_104_),
    .B(_115_),
    .C(_116_),
    .Y(\a[1] [1])
);

INVX1 _6376_ (
    .A(\genblk1[0].u_ce.Ycalc [10]),
    .Y(_117_)
);

NAND2X1 _6377_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(\genblk1[0].u_ce.Ycalc [8]),
    .Y(_118_)
);

OAI21X1 _6378_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(_117_),
    .C(_118_),
    .Y(_119_)
);

INVX1 _6379_ (
    .A(\genblk1[0].u_ce.Ycalc [6]),
    .Y(_120_)
);

INVX1 _6380_ (
    .A(\genblk1[0].u_ce.Ycalc [4]),
    .Y(_121_)
);

OAI22X1 _6381_ (
    .A(_96_),
    .B(_121_),
    .C(_120_),
    .D(_112_),
    .Y(_122_)
);

AOI21X1 _6382_ (
    .A(_92_),
    .B(_119_),
    .C(_122_),
    .Y(_123_)
);

AOI22X1 _6383_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[0].u_ce.Ycalc [0]),
    .C(_106_),
    .D(\genblk1[0].u_ce.Ycalc [2]),
    .Y(_124_)
);

OAI21X1 _6384_ (
    .A(_104_),
    .B(_123_),
    .C(_124_),
    .Y(\genblk1[0].u_ce.Y_ [0])
);

INVX1 _6385_ (
    .A(\genblk1[0].u_ce.Ycalc [11]),
    .Y(_125_)
);

NAND2X1 _6386_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(\genblk1[0].u_ce.Ycalc [9]),
    .Y(_126_)
);

OAI21X1 _6387_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(_125_),
    .C(_126_),
    .Y(_127_)
);

INVX1 _6388_ (
    .A(\genblk1[0].u_ce.Ycalc [7]),
    .Y(_128_)
);

INVX1 _6389_ (
    .A(\genblk1[0].u_ce.Ycalc [5]),
    .Y(_129_)
);

OAI22X1 _6390_ (
    .A(_96_),
    .B(_129_),
    .C(_128_),
    .D(_112_),
    .Y(_130_)
);

AOI21X1 _6391_ (
    .A(_92_),
    .B(_127_),
    .C(_130_),
    .Y(_131_)
);

AOI22X1 _6392_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[0].u_ce.Ycalc [1]),
    .C(_106_),
    .D(\genblk1[0].u_ce.Ycalc [3]),
    .Y(_132_)
);

OAI21X1 _6393_ (
    .A(_104_),
    .B(_131_),
    .C(_132_),
    .Y(\genblk1[0].u_ce.Y_ [1])
);

INVX1 _6394_ (
    .A(\genblk1[0].u_ce.Xcalc [2]),
    .Y(_133_)
);

INVX2 _6395_ (
    .A(_106_),
    .Y(_134_)
);

INVX1 _6396_ (
    .A(\genblk1[0].u_ce.Xcalc [4]),
    .Y(_135_)
);

INVX1 _6397_ (
    .A(\genblk1[0].u_ce.Xcalc [6]),
    .Y(_136_)
);

NOR2X1 _6398_ (
    .A(_98_),
    .B(_136_),
    .Y(_137_)
);

INVX1 _6399_ (
    .A(\genblk1[0].u_ce.Xcalc [8]),
    .Y(_138_)
);

NAND2X1 _6400_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(_138_),
    .Y(_139_)
);

OAI21X1 _6401_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(\genblk1[0].u_ce.Xcalc [10]),
    .C(_139_),
    .Y(_140_)
);

NOR2X1 _6402_ (
    .A(\genblk1[0].u_ce.LoadCtl [3]),
    .B(_140_),
    .Y(_141_)
);

OAI21X1 _6403_ (
    .A(_137_),
    .B(_141_),
    .C(_96_),
    .Y(_142_)
);

OAI21X1 _6404_ (
    .A(_96_),
    .B(_135_),
    .C(_142_),
    .Y(_143_)
);

AOI22X1 _6405_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[0].u_ce.Xcalc [0]),
    .C(_143_),
    .D(_103_),
    .Y(_144_)
);

OAI21X1 _6406_ (
    .A(_133_),
    .B(_134_),
    .C(_144_),
    .Y(\genblk1[0].u_ce.X_ [0])
);

INVX1 _6407_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .Y(_145_)
);

INVX1 _6408_ (
    .A(\genblk1[0].u_ce.Xcalc [9]),
    .Y(_146_)
);

NAND2X1 _6409_ (
    .A(\genblk1[0].u_ce.Xcalc [11]),
    .B(_145_),
    .Y(_147_)
);

OAI21X1 _6410_ (
    .A(_145_),
    .B(_146_),
    .C(_147_),
    .Y(_148_)
);

INVX1 _6411_ (
    .A(\genblk1[0].u_ce.Xcalc [7]),
    .Y(_149_)
);

INVX1 _6412_ (
    .A(\genblk1[0].u_ce.Xcalc [5]),
    .Y(_150_)
);

OAI22X1 _6413_ (
    .A(_96_),
    .B(_150_),
    .C(_149_),
    .D(_112_),
    .Y(_151_)
);

AOI21X1 _6414_ (
    .A(_92_),
    .B(_148_),
    .C(_151_),
    .Y(_152_)
);

AOI22X1 _6415_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[0].u_ce.Xcalc [1]),
    .C(_106_),
    .D(\genblk1[0].u_ce.Xcalc [3]),
    .Y(_153_)
);

OAI21X1 _6416_ (
    .A(_104_),
    .B(_152_),
    .C(_153_),
    .Y(\genblk1[0].u_ce.X_ [1])
);

INVX1 _6417_ (
    .A(\genblk1[0].u_ce.Ain0 [0]),
    .Y(_154_)
);

NAND2X1 _6418_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\a[0] [0]),
    .Y(_155_)
);

OAI21X1 _6419_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_154_),
    .C(_155_),
    .Y(_0_)
);

INVX1 _6420_ (
    .A(\genblk1[0].u_ce.Ain0 [1]),
    .Y(_156_)
);

NAND2X1 _6421_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\a[0] [1]),
    .Y(_157_)
);

OAI21X1 _6422_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_156_),
    .C(_157_),
    .Y(_1_)
);

INVX8 _6423_ (
    .A(\genblk1[0].u_ce.Vld_bF$buf4 ),
    .Y(_158_)
);

NAND2X1 _6424_ (
    .A(\genblk1[0].u_ce.Ycalc [2]),
    .B(_158__bF$buf4),
    .Y(_159_)
);

INVX2 _6425_ (
    .A(1'h0),
    .Y(_160_)
);

NOR2X1 _6426_ (
    .A(1'h0),
    .B(1'h0),
    .Y(_161_)
);

NAND2X1 _6427_ (
    .A(_160_),
    .B(_161_),
    .Y(_162_)
);

INVX2 _6428_ (
    .A(_162_),
    .Y(_163_)
);

INVX8 _6429_ (
    .A(1'h0),
    .Y(_164_)
);

MUX2X1 _6430_ (
    .A(\genblk1[0].u_ce.Xin12b [4]),
    .B(\genblk1[0].u_ce.Xin1 [1]),
    .S(1'h0),
    .Y(_165_)
);

MUX2X1 _6431_ (
    .A(\genblk1[0].u_ce.Xin1 [0]),
    .B(\genblk1[0].u_ce.Xin0 [1]),
    .S(1'h0),
    .Y(_166_)
);

MUX2X1 _6432_ (
    .A(_166_),
    .B(_165_),
    .S(_164__bF$buf4),
    .Y(_167_)
);

MUX2X1 _6433_ (
    .A(\genblk1[0].u_ce.Xin12b [8]),
    .B(\genblk1[0].u_ce.Xin12b [7]),
    .S(1'h0),
    .Y(_168_)
);

MUX2X1 _6434_ (
    .A(\genblk1[0].u_ce.Xin12b [6]),
    .B(\genblk1[0].u_ce.Xin12b [5]),
    .S(1'h0),
    .Y(_169_)
);

MUX2X1 _6435_ (
    .A(_169_),
    .B(_168_),
    .S(_164__bF$buf3),
    .Y(_170_)
);

MUX2X1 _6436_ (
    .A(_170_),
    .B(_167_),
    .S(1'h0),
    .Y(_171_)
);

INVX1 _6437_ (
    .A(_171_),
    .Y(_172_)
);

MUX2X1 _6438_ (
    .A(\genblk1[0].u_ce.Xin1 [1]),
    .B(\genblk1[0].u_ce.Xin1 [0]),
    .S(1'h0),
    .Y(_173_)
);

MUX2X1 _6439_ (
    .A(\genblk1[0].u_ce.Xin0 [1]),
    .B(\genblk1[0].u_ce.Xin0 [0]),
    .S(1'h0),
    .Y(_174_)
);

MUX2X1 _6440_ (
    .A(_174_),
    .B(_173_),
    .S(_164__bF$buf2),
    .Y(_175_)
);

MUX2X1 _6441_ (
    .A(\genblk1[0].u_ce.Xin12b [7]),
    .B(\genblk1[0].u_ce.Xin12b [6]),
    .S(1'h0),
    .Y(_176_)
);

MUX2X1 _6442_ (
    .A(\genblk1[0].u_ce.Xin12b [5]),
    .B(\genblk1[0].u_ce.Xin12b [4]),
    .S(1'h0),
    .Y(_177_)
);

MUX2X1 _6443_ (
    .A(_177_),
    .B(_176_),
    .S(_164__bF$buf1),
    .Y(_178_)
);

MUX2X1 _6444_ (
    .A(_178_),
    .B(_175_),
    .S(1'h0),
    .Y(_179_)
);

OAI21X1 _6445_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf4 ),
    .B(_179_),
    .C(_172_),
    .Y(_180_)
);

NOR2X1 _6446_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .B(_179_),
    .Y(_181_)
);

NAND2X1 _6447_ (
    .A(_171_),
    .B(_181_),
    .Y(_182_)
);

NAND3X1 _6448_ (
    .A(\genblk1[0].u_ce.Yin0 [1]),
    .B(_180_),
    .C(_182_),
    .Y(_183_)
);

NOR2X1 _6449_ (
    .A(\genblk1[0].u_ce.Yin0 [0]),
    .B(_179_),
    .Y(_184_)
);

AOI21X1 _6450_ (
    .A(_182_),
    .B(_180_),
    .C(\genblk1[0].u_ce.Yin0 [1]),
    .Y(_185_)
);

OAI21X1 _6451_ (
    .A(_184_),
    .B(_185_),
    .C(_183_),
    .Y(_186_)
);

INVX1 _6452_ (
    .A(\genblk1[0].u_ce.Yin1 [0]),
    .Y(_187_)
);

MUX2X1 _6453_ (
    .A(\genblk1[0].u_ce.Xin12b [9]),
    .B(\genblk1[0].u_ce.Xin12b [8]),
    .S(1'h0),
    .Y(_188_)
);

MUX2X1 _6454_ (
    .A(_188_),
    .B(_176_),
    .S(1'h0),
    .Y(_189_)
);

AND2X2 _6455_ (
    .A(_189_),
    .B(1'h0),
    .Y(_190_)
);

INVX4 _6456_ (
    .A(1'h0),
    .Y(_191_)
);

NAND2X1 _6457_ (
    .A(_191__bF$buf3),
    .B(_164__bF$buf0),
    .Y(_192_)
);

NAND2X1 _6458_ (
    .A(1'h0),
    .B(_191__bF$buf2),
    .Y(_193_)
);

OAI22X1 _6459_ (
    .A(_192_),
    .B(_173_),
    .C(_177_),
    .D(_193_),
    .Y(_194_)
);

INVX1 _6460_ (
    .A(\genblk1[0].u_ce.Xin1 [1]),
    .Y(_195_)
);

NAND2X1 _6461_ (
    .A(_160_),
    .B(_195_),
    .Y(_196_)
);

INVX1 _6462_ (
    .A(\genblk1[0].u_ce.Xin12b [4]),
    .Y(_197_)
);

NAND2X1 _6463_ (
    .A(1'h0),
    .B(_197_),
    .Y(_198_)
);

NAND3X1 _6464_ (
    .A(1'h0),
    .B(_198_),
    .C(_196_),
    .Y(_199_)
);

INVX1 _6465_ (
    .A(\genblk1[0].u_ce.Xin0 [1]),
    .Y(_200_)
);

NAND2X1 _6466_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Xin1 [0]),
    .Y(_201_)
);

OAI21X1 _6467_ (
    .A(1'h0),
    .B(_200_),
    .C(_201_),
    .Y(_202_)
);

NAND2X1 _6468_ (
    .A(_164__bF$buf4),
    .B(_202_),
    .Y(_203_)
);

NAND3X1 _6469_ (
    .A(_191__bF$buf1),
    .B(_199_),
    .C(_203_),
    .Y(_204_)
);

INVX1 _6470_ (
    .A(\genblk1[0].u_ce.Xin12b [5]),
    .Y(_205_)
);

NAND2X1 _6471_ (
    .A(_160_),
    .B(_205_),
    .Y(_206_)
);

INVX1 _6472_ (
    .A(\genblk1[0].u_ce.Xin12b [6]),
    .Y(_207_)
);

NAND2X1 _6473_ (
    .A(1'h0),
    .B(_207_),
    .Y(_208_)
);

NAND3X1 _6474_ (
    .A(_164__bF$buf3),
    .B(_208_),
    .C(_206_),
    .Y(_209_)
);

INVX1 _6475_ (
    .A(\genblk1[0].u_ce.Xin12b [7]),
    .Y(_210_)
);

NAND2X1 _6476_ (
    .A(_160_),
    .B(_210_),
    .Y(_211_)
);

INVX1 _6477_ (
    .A(\genblk1[0].u_ce.Xin12b [8]),
    .Y(_212_)
);

NAND2X1 _6478_ (
    .A(1'h0),
    .B(_212_),
    .Y(_213_)
);

NAND3X1 _6479_ (
    .A(1'h0),
    .B(_213_),
    .C(_211_),
    .Y(_214_)
);

NAND3X1 _6480_ (
    .A(1'h0),
    .B(_209_),
    .C(_214_),
    .Y(_215_)
);

INVX1 _6481_ (
    .A(\genblk1[0].u_ce.Xin1 [0]),
    .Y(_216_)
);

NAND2X1 _6482_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Xin1 [1]),
    .Y(_217_)
);

OAI21X1 _6483_ (
    .A(1'h0),
    .B(_216_),
    .C(_217_),
    .Y(_218_)
);

NAND2X1 _6484_ (
    .A(1'h0),
    .B(_218_),
    .Y(_219_)
);

INVX1 _6485_ (
    .A(\genblk1[0].u_ce.Xin0 [0]),
    .Y(_220_)
);

NAND2X1 _6486_ (
    .A(\genblk1[0].u_ce.Xin0 [1]),
    .B(1'h0),
    .Y(_221_)
);

OAI21X1 _6487_ (
    .A(1'h0),
    .B(_220_),
    .C(_221_),
    .Y(_222_)
);

NAND2X1 _6488_ (
    .A(_164__bF$buf2),
    .B(_222_),
    .Y(_223_)
);

NAND3X1 _6489_ (
    .A(_191__bF$buf0),
    .B(_219_),
    .C(_223_),
    .Y(_224_)
);

NAND2X1 _6490_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Xin12b [5]),
    .Y(_225_)
);

OAI21X1 _6491_ (
    .A(1'h0),
    .B(_197_),
    .C(_225_),
    .Y(_226_)
);

NAND2X1 _6492_ (
    .A(_164__bF$buf1),
    .B(_226_),
    .Y(_227_)
);

NAND2X1 _6493_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Xin12b [7]),
    .Y(_228_)
);

OAI21X1 _6494_ (
    .A(1'h0),
    .B(_207_),
    .C(_228_),
    .Y(_229_)
);

NAND2X1 _6495_ (
    .A(1'h0),
    .B(_229_),
    .Y(_230_)
);

NAND3X1 _6496_ (
    .A(1'h0),
    .B(_227_),
    .C(_230_),
    .Y(_231_)
);

AOI22X1 _6497_ (
    .A(_204_),
    .B(_215_),
    .C(_224_),
    .D(_231_),
    .Y(_232_)
);

NOR2X1 _6498_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_232_),
    .Y(_233_)
);

OAI21X1 _6499_ (
    .A(_190_),
    .B(_194_),
    .C(_233_),
    .Y(_234_)
);

AOI21X1 _6500_ (
    .A(1'h0),
    .B(_189_),
    .C(_194_),
    .Y(_235_)
);

OAI21X1 _6501_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .B(_232_),
    .C(_235_),
    .Y(_236_)
);

NAND3X1 _6502_ (
    .A(_187_),
    .B(_236_),
    .C(_234_),
    .Y(_237_)
);

NAND2X1 _6503_ (
    .A(_235_),
    .B(_233_),
    .Y(_238_)
);

OAI22X1 _6504_ (
    .A(_190_),
    .B(_194_),
    .C(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .D(_232_),
    .Y(_239_)
);

NAND3X1 _6505_ (
    .A(\genblk1[0].u_ce.Yin1 [0]),
    .B(_239_),
    .C(_238_),
    .Y(_240_)
);

NAND3X1 _6506_ (
    .A(_237_),
    .B(_240_),
    .C(_186_),
    .Y(_241_)
);

INVX1 _6507_ (
    .A(\genblk1[0].u_ce.Yin0 [1]),
    .Y(_242_)
);

NAND2X1 _6508_ (
    .A(_172_),
    .B(_181_),
    .Y(_243_)
);

OAI21X1 _6509_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf4 ),
    .B(_179_),
    .C(_171_),
    .Y(_244_)
);

AOI21X1 _6510_ (
    .A(_243_),
    .B(_244_),
    .C(_242_),
    .Y(_245_)
);

INVX1 _6511_ (
    .A(_184_),
    .Y(_246_)
);

NAND3X1 _6512_ (
    .A(_242_),
    .B(_244_),
    .C(_243_),
    .Y(_247_)
);

AOI21X1 _6513_ (
    .A(_246_),
    .B(_247_),
    .C(_245_),
    .Y(_248_)
);

AOI21X1 _6514_ (
    .A(_238_),
    .B(_239_),
    .C(\genblk1[0].u_ce.Yin1 [0]),
    .Y(_249_)
);

AOI21X1 _6515_ (
    .A(_234_),
    .B(_236_),
    .C(_187_),
    .Y(_250_)
);

OAI21X1 _6516_ (
    .A(_249_),
    .B(_250_),
    .C(_248_),
    .Y(_251_)
);

AOI21X1 _6517_ (
    .A(_241_),
    .B(_251_),
    .C(_163_),
    .Y(_252_)
);

INVX8 _6518_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_253_)
);

NAND3X1 _6519_ (
    .A(_191__bF$buf3),
    .B(_160_),
    .C(_253__bF$buf5),
    .Y(_254_)
);

OAI21X1 _6520_ (
    .A(1'h0),
    .B(_254_),
    .C(\genblk1[0].u_ce.Vld_bF$buf3 ),
    .Y(_255_)
);

OAI21X1 _6521_ (
    .A(_255_),
    .B(_252_),
    .C(_159_),
    .Y(_2_)
);

INVX1 _6522_ (
    .A(\genblk1[0].u_ce.Ycalc [3]),
    .Y(_256_)
);

INVX1 _6523_ (
    .A(\genblk1[0].u_ce.Xin12b [9]),
    .Y(_257_)
);

NAND2X1 _6524_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Xin12b [10]),
    .Y(_258_)
);

OAI21X1 _6525_ (
    .A(1'h0),
    .B(_257_),
    .C(_258_),
    .Y(_259_)
);

NAND2X1 _6526_ (
    .A(1'h0),
    .B(_259_),
    .Y(_260_)
);

OAI21X1 _6527_ (
    .A(1'h0),
    .B(_168_),
    .C(_260_),
    .Y(_261_)
);

OAI22X1 _6528_ (
    .A(_192_),
    .B(_165_),
    .C(_169_),
    .D(_193_),
    .Y(_262_)
);

AOI21X1 _6529_ (
    .A(_261_),
    .B(1'h0),
    .C(_262_),
    .Y(_263_)
);

NAND3X1 _6530_ (
    .A(_235_),
    .B(_171_),
    .C(_179_),
    .Y(_264_)
);

INVX1 _6531_ (
    .A(_264_),
    .Y(_265_)
);

NOR2X1 _6532_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_265_),
    .Y(_266_)
);

NAND2X1 _6533_ (
    .A(_263_),
    .B(_266_),
    .Y(_267_)
);

INVX1 _6534_ (
    .A(_263_),
    .Y(_268_)
);

OAI21X1 _6535_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .B(_265_),
    .C(_268_),
    .Y(_269_)
);

AOI21X1 _6536_ (
    .A(_267_),
    .B(_269_),
    .C(\genblk1[0].u_ce.Yin1 [1]),
    .Y(_270_)
);

AOI21X1 _6537_ (
    .A(_186_),
    .B(_237_),
    .C(_250_),
    .Y(_271_)
);

NAND3X1 _6538_ (
    .A(\genblk1[0].u_ce.Yin1 [1]),
    .B(_269_),
    .C(_267_),
    .Y(_272_)
);

NAND2X1 _6539_ (
    .A(_272_),
    .B(_271_),
    .Y(_273_)
);

OAI21X1 _6540_ (
    .A(_249_),
    .B(_248_),
    .C(_240_),
    .Y(_274_)
);

INVX1 _6541_ (
    .A(\genblk1[0].u_ce.Yin1 [1]),
    .Y(_275_)
);

NAND2X1 _6542_ (
    .A(_268_),
    .B(_266_),
    .Y(_276_)
);

OAI21X1 _6543_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .B(_265_),
    .C(_263_),
    .Y(_277_)
);

AOI21X1 _6544_ (
    .A(_276_),
    .B(_277_),
    .C(_275_),
    .Y(_278_)
);

OAI21X1 _6545_ (
    .A(_270_),
    .B(_278_),
    .C(_274_),
    .Y(_279_)
);

OAI21X1 _6546_ (
    .A(_270_),
    .B(_273_),
    .C(_279_),
    .Y(_280_)
);

OAI21X1 _6547_ (
    .A(_253__bF$buf4),
    .B(_162_),
    .C(\genblk1[0].u_ce.Vld_bF$buf2 ),
    .Y(_281_)
);

INVX1 _6548_ (
    .A(_281_),
    .Y(_282_)
);

OAI21X1 _6549_ (
    .A(_163_),
    .B(_280_),
    .C(_282_),
    .Y(_283_)
);

OAI21X1 _6550_ (
    .A(_256_),
    .B(\genblk1[0].u_ce.Vld_bF$buf1 ),
    .C(_283_),
    .Y(_3_)
);

INVX1 _6551_ (
    .A(_255_),
    .Y(_284_)
);

INVX1 _6552_ (
    .A(\genblk1[0].u_ce.Yin12b [4]),
    .Y(_285_)
);

NAND3X1 _6553_ (
    .A(_235_),
    .B(_263_),
    .C(_232_),
    .Y(_286_)
);

INVX1 _6554_ (
    .A(\genblk1[0].u_ce.Xin12b [10]),
    .Y(_287_)
);

NAND2X1 _6555_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Xin12b [11]),
    .Y(_288_)
);

OAI21X1 _6556_ (
    .A(1'h0),
    .B(_287_),
    .C(_288_),
    .Y(_289_)
);

NAND2X1 _6557_ (
    .A(_164__bF$buf0),
    .B(_188_),
    .Y(_290_)
);

OAI21X1 _6558_ (
    .A(_164__bF$buf4),
    .B(_289_),
    .C(_290_),
    .Y(_291_)
);

NAND2X1 _6559_ (
    .A(_191__bF$buf2),
    .B(_178_),
    .Y(_292_)
);

OAI21X1 _6560_ (
    .A(_191__bF$buf1),
    .B(_291_),
    .C(_292_),
    .Y(_293_)
);

INVX1 _6561_ (
    .A(_293_),
    .Y(_294_)
);

NAND3X1 _6562_ (
    .A(_253__bF$buf3),
    .B(_294_),
    .C(_286_),
    .Y(_295_)
);

INVX1 _6563_ (
    .A(_295_),
    .Y(_296_)
);

AOI21X1 _6564_ (
    .A(_286_),
    .B(_253__bF$buf2),
    .C(_294_),
    .Y(_297_)
);

OAI21X1 _6565_ (
    .A(_297_),
    .B(_296_),
    .C(_285_),
    .Y(_298_)
);

OAI21X1 _6566_ (
    .A(_264_),
    .B(_268_),
    .C(_253__bF$buf1),
    .Y(_299_)
);

NAND2X1 _6567_ (
    .A(_293_),
    .B(_299_),
    .Y(_300_)
);

NAND3X1 _6568_ (
    .A(\genblk1[0].u_ce.Yin12b [4]),
    .B(_295_),
    .C(_300_),
    .Y(_301_)
);

NAND2X1 _6569_ (
    .A(_301_),
    .B(_298_),
    .Y(_302_)
);

INVX1 _6570_ (
    .A(_270_),
    .Y(_303_)
);

OAI21X1 _6571_ (
    .A(_278_),
    .B(_274_),
    .C(_303_),
    .Y(_304_)
);

AOI21X1 _6572_ (
    .A(_304_),
    .B(_302_),
    .C(_163_),
    .Y(_305_)
);

OAI21X1 _6573_ (
    .A(_302_),
    .B(_304_),
    .C(_305_),
    .Y(_306_)
);

AOI22X1 _6574_ (
    .A(_121_),
    .B(_158__bF$buf3),
    .C(_306_),
    .D(_284_),
    .Y(_4_)
);

INVX1 _6575_ (
    .A(_301_),
    .Y(_307_)
);

AOI21X1 _6576_ (
    .A(_271_),
    .B(_272_),
    .C(_270_),
    .Y(_308_)
);

AOI21X1 _6577_ (
    .A(_308_),
    .B(_298_),
    .C(_307_),
    .Y(_309_)
);

INVX1 _6578_ (
    .A(\genblk1[0].u_ce.Yin12b [5]),
    .Y(_310_)
);

NAND3X1 _6579_ (
    .A(_263_),
    .B(_294_),
    .C(_265_),
    .Y(_311_)
);

INVX1 _6580_ (
    .A(\genblk1[0].u_ce.Xin12b [11]),
    .Y(_312_)
);

NOR2X1 _6581_ (
    .A(_164__bF$buf3),
    .B(_312_),
    .Y(_313_)
);

AOI21X1 _6582_ (
    .A(_164__bF$buf2),
    .B(_259_),
    .C(_313_),
    .Y(_314_)
);

NAND2X1 _6583_ (
    .A(_191__bF$buf0),
    .B(_170_),
    .Y(_315_)
);

OAI21X1 _6584_ (
    .A(_191__bF$buf3),
    .B(_314_),
    .C(_315_),
    .Y(_316_)
);

NAND3X1 _6585_ (
    .A(_253__bF$buf0),
    .B(_316_),
    .C(_311_),
    .Y(_317_)
);

INVX1 _6586_ (
    .A(_316_),
    .Y(_318_)
);

OAI21X1 _6587_ (
    .A(_293_),
    .B(_286_),
    .C(_253__bF$buf5),
    .Y(_319_)
);

NAND2X1 _6588_ (
    .A(_318_),
    .B(_319_),
    .Y(_320_)
);

NAND3X1 _6589_ (
    .A(_310_),
    .B(_320_),
    .C(_317_),
    .Y(_321_)
);

NAND3X1 _6590_ (
    .A(_253__bF$buf4),
    .B(_318_),
    .C(_311_),
    .Y(_322_)
);

NAND2X1 _6591_ (
    .A(_316_),
    .B(_319_),
    .Y(_323_)
);

NAND3X1 _6592_ (
    .A(\genblk1[0].u_ce.Yin12b [5]),
    .B(_323_),
    .C(_322_),
    .Y(_324_)
);

NAND2X1 _6593_ (
    .A(_321_),
    .B(_324_),
    .Y(_325_)
);

INVX1 _6594_ (
    .A(_325_),
    .Y(_326_)
);

NOR2X1 _6595_ (
    .A(_326_),
    .B(_309_),
    .Y(_327_)
);

OAI21X1 _6596_ (
    .A(_302_),
    .B(_304_),
    .C(_301_),
    .Y(_328_)
);

OAI21X1 _6597_ (
    .A(_325_),
    .B(_328_),
    .C(_162_),
    .Y(_329_)
);

OAI21X1 _6598_ (
    .A(_329_),
    .B(_327_),
    .C(_284_),
    .Y(_330_)
);

OAI21X1 _6599_ (
    .A(_129_),
    .B(\genblk1[0].u_ce.Vld_bF$buf0 ),
    .C(_330_),
    .Y(_5_)
);

NOR2X1 _6600_ (
    .A(_302_),
    .B(_325_),
    .Y(_331_)
);

OAI21X1 _6601_ (
    .A(_301_),
    .B(_325_),
    .C(_324_),
    .Y(_332_)
);

AOI21X1 _6602_ (
    .A(_331_),
    .B(_308_),
    .C(_332_),
    .Y(_333_)
);

INVX1 _6603_ (
    .A(\genblk1[0].u_ce.Yin12b [6]),
    .Y(_334_)
);

NOR2X1 _6604_ (
    .A(_293_),
    .B(_286_),
    .Y(_335_)
);

NAND2X1 _6605_ (
    .A(_318_),
    .B(_335_),
    .Y(_336_)
);

AOI21X1 _6606_ (
    .A(_164__bF$buf1),
    .B(_289_),
    .C(_313_),
    .Y(_337_)
);

NAND2X1 _6607_ (
    .A(_191__bF$buf2),
    .B(_189_),
    .Y(_338_)
);

OAI21X1 _6608_ (
    .A(_191__bF$buf1),
    .B(_337_),
    .C(_338_),
    .Y(_339_)
);

NAND3X1 _6609_ (
    .A(_253__bF$buf3),
    .B(_339_),
    .C(_336_),
    .Y(_340_)
);

NOR3X1 _6610_ (
    .A(_293_),
    .B(_316_),
    .C(_286_),
    .Y(_341_)
);

INVX1 _6611_ (
    .A(_339_),
    .Y(_342_)
);

OAI21X1 _6612_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf4 ),
    .B(_341_),
    .C(_342_),
    .Y(_343_)
);

NAND3X1 _6613_ (
    .A(_334_),
    .B(_343_),
    .C(_340_),
    .Y(_344_)
);

NAND3X1 _6614_ (
    .A(_253__bF$buf2),
    .B(_342_),
    .C(_336_),
    .Y(_345_)
);

OAI21X1 _6615_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .B(_341_),
    .C(_339_),
    .Y(_346_)
);

NAND3X1 _6616_ (
    .A(\genblk1[0].u_ce.Yin12b [6]),
    .B(_346_),
    .C(_345_),
    .Y(_347_)
);

AND2X2 _6617_ (
    .A(_344_),
    .B(_347_),
    .Y(_348_)
);

INVX1 _6618_ (
    .A(_348_),
    .Y(_349_)
);

AOI21X1 _6619_ (
    .A(_333_),
    .B(_349_),
    .C(_163_),
    .Y(_350_)
);

OAI21X1 _6620_ (
    .A(_333_),
    .B(_349_),
    .C(_350_),
    .Y(_351_)
);

AOI22X1 _6621_ (
    .A(_120_),
    .B(_158__bF$buf2),
    .C(_351_),
    .D(_284_),
    .Y(_6_)
);

AND2X2 _6622_ (
    .A(_298_),
    .B(_301_),
    .Y(_352_)
);

NAND3X1 _6623_ (
    .A(_321_),
    .B(_324_),
    .C(_352_),
    .Y(_353_)
);

INVX1 _6624_ (
    .A(_324_),
    .Y(_354_)
);

AOI21X1 _6625_ (
    .A(_307_),
    .B(_321_),
    .C(_354_),
    .Y(_355_)
);

OAI21X1 _6626_ (
    .A(_304_),
    .B(_353_),
    .C(_355_),
    .Y(_356_)
);

INVX1 _6627_ (
    .A(_347_),
    .Y(_357_)
);

AOI21X1 _6628_ (
    .A(_356_),
    .B(_344_),
    .C(_357_),
    .Y(_358_)
);

INVX1 _6629_ (
    .A(\genblk1[0].u_ce.Yin12b [7]),
    .Y(_359_)
);

NAND2X1 _6630_ (
    .A(_342_),
    .B(_341_),
    .Y(_360_)
);

NOR2X1 _6631_ (
    .A(_191__bF$buf0),
    .B(_312_),
    .Y(_361_)
);

AOI21X1 _6632_ (
    .A(_261_),
    .B(_191__bF$buf3),
    .C(_361_),
    .Y(_362_)
);

INVX1 _6633_ (
    .A(_362_),
    .Y(_363_)
);

NAND3X1 _6634_ (
    .A(_253__bF$buf1),
    .B(_363_),
    .C(_360_),
    .Y(_364_)
);

AND2X2 _6635_ (
    .A(_341_),
    .B(_342_),
    .Y(_365_)
);

OAI21X1 _6636_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_365_),
    .C(_362_),
    .Y(_366_)
);

NAND3X1 _6637_ (
    .A(_359_),
    .B(_364_),
    .C(_366_),
    .Y(_367_)
);

NAND3X1 _6638_ (
    .A(_253__bF$buf0),
    .B(_362_),
    .C(_360_),
    .Y(_368_)
);

OAI21X1 _6639_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .B(_365_),
    .C(_363_),
    .Y(_369_)
);

NAND3X1 _6640_ (
    .A(\genblk1[0].u_ce.Yin12b [7]),
    .B(_368_),
    .C(_369_),
    .Y(_370_)
);

AND2X2 _6641_ (
    .A(_367_),
    .B(_370_),
    .Y(_371_)
);

NOR2X1 _6642_ (
    .A(_371_),
    .B(_358_),
    .Y(_372_)
);

NAND2X1 _6643_ (
    .A(_160_),
    .B(_164__bF$buf0),
    .Y(_373_)
);

NAND2X1 _6644_ (
    .A(_371_),
    .B(_358_),
    .Y(_374_)
);

OAI21X1 _6645_ (
    .A(1'h0),
    .B(_373_),
    .C(_374_),
    .Y(_375_)
);

OAI21X1 _6646_ (
    .A(_372_),
    .B(_375_),
    .C(_282_),
    .Y(_376_)
);

OAI21X1 _6647_ (
    .A(_128_),
    .B(\genblk1[0].u_ce.Vld_bF$buf4 ),
    .C(_376_),
    .Y(_7_)
);

INVX1 _6648_ (
    .A(\genblk1[0].u_ce.Ycalc [8]),
    .Y(_377_)
);

AOI21X1 _6649_ (
    .A(_366_),
    .B(_364_),
    .C(_359_),
    .Y(_378_)
);

OAI21X1 _6650_ (
    .A(_357_),
    .B(_378_),
    .C(_367_),
    .Y(_379_)
);

NAND3X1 _6651_ (
    .A(_348_),
    .B(_371_),
    .C(_356_),
    .Y(_380_)
);

INVX1 _6652_ (
    .A(\genblk1[0].u_ce.Yin12b [8]),
    .Y(_381_)
);

NAND3X1 _6653_ (
    .A(_342_),
    .B(_362_),
    .C(_341_),
    .Y(_382_)
);

INVX1 _6654_ (
    .A(_361_),
    .Y(_383_)
);

OAI21X1 _6655_ (
    .A(1'h0),
    .B(_291_),
    .C(_383_),
    .Y(_384_)
);

NAND3X1 _6656_ (
    .A(_253__bF$buf5),
    .B(_384_),
    .C(_382_),
    .Y(_385_)
);

INVX1 _6657_ (
    .A(_384_),
    .Y(_386_)
);

NAND2X1 _6658_ (
    .A(_253__bF$buf4),
    .B(_382_),
    .Y(_387_)
);

NAND2X1 _6659_ (
    .A(_386_),
    .B(_387_),
    .Y(_388_)
);

NAND3X1 _6660_ (
    .A(_381_),
    .B(_385_),
    .C(_388_),
    .Y(_389_)
);

NAND3X1 _6661_ (
    .A(_253__bF$buf3),
    .B(_386_),
    .C(_382_),
    .Y(_390_)
);

NAND2X1 _6662_ (
    .A(_384_),
    .B(_387_),
    .Y(_391_)
);

NAND3X1 _6663_ (
    .A(\genblk1[0].u_ce.Yin12b [8]),
    .B(_390_),
    .C(_391_),
    .Y(_392_)
);

AND2X2 _6664_ (
    .A(_389_),
    .B(_392_),
    .Y(_393_)
);

INVX1 _6665_ (
    .A(_393_),
    .Y(_394_)
);

AOI21X1 _6666_ (
    .A(_380_),
    .B(_379_),
    .C(_394_),
    .Y(_395_)
);

NAND3X1 _6667_ (
    .A(_367_),
    .B(_370_),
    .C(_348_),
    .Y(_396_)
);

OAI21X1 _6668_ (
    .A(_396_),
    .B(_333_),
    .C(_379_),
    .Y(_397_)
);

OAI21X1 _6669_ (
    .A(_393_),
    .B(_397_),
    .C(_162_),
    .Y(_398_)
);

OR2X2 _6670_ (
    .A(_398_),
    .B(_395_),
    .Y(_399_)
);

AOI22X1 _6671_ (
    .A(_377_),
    .B(_158__bF$buf1),
    .C(_399_),
    .D(_282_),
    .Y(_8_)
);

INVX1 _6672_ (
    .A(\genblk1[0].u_ce.Ycalc [9]),
    .Y(_400_)
);

INVX1 _6673_ (
    .A(_392_),
    .Y(_401_)
);

NOR2X1 _6674_ (
    .A(_401_),
    .B(_395_),
    .Y(_402_)
);

INVX1 _6675_ (
    .A(\genblk1[0].u_ce.Yin12b [9]),
    .Y(_403_)
);

OAI21X1 _6676_ (
    .A(1'h0),
    .B(_314_),
    .C(_383_),
    .Y(_404_)
);

INVX1 _6677_ (
    .A(_404_),
    .Y(_405_)
);

OAI21X1 _6678_ (
    .A(_384_),
    .B(_382_),
    .C(_253__bF$buf2),
    .Y(_406_)
);

NAND2X1 _6679_ (
    .A(_405_),
    .B(_406_),
    .Y(_407_)
);

NAND3X1 _6680_ (
    .A(_362_),
    .B(_386_),
    .C(_365_),
    .Y(_408_)
);

NAND3X1 _6681_ (
    .A(_253__bF$buf1),
    .B(_404_),
    .C(_408_),
    .Y(_409_)
);

NAND3X1 _6682_ (
    .A(_403_),
    .B(_407_),
    .C(_409_),
    .Y(_410_)
);

AND2X2 _6683_ (
    .A(_406_),
    .B(_405_),
    .Y(_411_)
);

NOR2X1 _6684_ (
    .A(_405_),
    .B(_406_),
    .Y(_412_)
);

OAI21X1 _6685_ (
    .A(_412_),
    .B(_411_),
    .C(\genblk1[0].u_ce.Yin12b [9]),
    .Y(_413_)
);

NAND2X1 _6686_ (
    .A(_410_),
    .B(_413_),
    .Y(_414_)
);

AOI21X1 _6687_ (
    .A(_402_),
    .B(_414_),
    .C(_163_),
    .Y(_415_)
);

OAI21X1 _6688_ (
    .A(_402_),
    .B(_414_),
    .C(_415_),
    .Y(_416_)
);

AOI22X1 _6689_ (
    .A(_400_),
    .B(_158__bF$buf0),
    .C(_416_),
    .D(_282_),
    .Y(_9_)
);

OAI21X1 _6690_ (
    .A(_392_),
    .B(_414_),
    .C(_413_),
    .Y(_417_)
);

NAND3X1 _6691_ (
    .A(_410_),
    .B(_413_),
    .C(_393_),
    .Y(_418_)
);

AOI21X1 _6692_ (
    .A(_379_),
    .B(_380_),
    .C(_418_),
    .Y(_419_)
);

INVX1 _6693_ (
    .A(\genblk1[0].u_ce.Yin12b [10]),
    .Y(_420_)
);

OAI21X1 _6694_ (
    .A(1'h0),
    .B(_337_),
    .C(_383_),
    .Y(_421_)
);

INVX1 _6695_ (
    .A(_421_),
    .Y(_422_)
);

OAI21X1 _6696_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .B(_405_),
    .C(_406_),
    .Y(_423_)
);

NAND2X1 _6697_ (
    .A(_422_),
    .B(_423_),
    .Y(_424_)
);

OAI21X1 _6698_ (
    .A(_404_),
    .B(_408_),
    .C(_253__bF$buf0),
    .Y(_425_)
);

NAND2X1 _6699_ (
    .A(_421_),
    .B(_425_),
    .Y(_426_)
);

NAND2X1 _6700_ (
    .A(_424_),
    .B(_426_),
    .Y(_427_)
);

NAND2X1 _6701_ (
    .A(_420_),
    .B(_427_),
    .Y(_428_)
);

NAND3X1 _6702_ (
    .A(\genblk1[0].u_ce.Yin12b [10]),
    .B(_424_),
    .C(_426_),
    .Y(_429_)
);

AND2X2 _6703_ (
    .A(_428_),
    .B(_429_),
    .Y(_430_)
);

OAI21X1 _6704_ (
    .A(_417_),
    .B(_419_),
    .C(_430_),
    .Y(_431_)
);

INVX1 _6705_ (
    .A(_413_),
    .Y(_432_)
);

AOI21X1 _6706_ (
    .A(_401_),
    .B(_410_),
    .C(_432_),
    .Y(_433_)
);

AND2X2 _6707_ (
    .A(_413_),
    .B(_410_),
    .Y(_434_)
);

NAND3X1 _6708_ (
    .A(_393_),
    .B(_434_),
    .C(_397_),
    .Y(_435_)
);

NAND2X1 _6709_ (
    .A(_429_),
    .B(_428_),
    .Y(_436_)
);

NAND3X1 _6710_ (
    .A(_433_),
    .B(_436_),
    .C(_435_),
    .Y(_437_)
);

NAND3X1 _6711_ (
    .A(_162_),
    .B(_437_),
    .C(_431_),
    .Y(_438_)
);

AOI22X1 _6712_ (
    .A(_117_),
    .B(_158__bF$buf4),
    .C(_438_),
    .D(_284_),
    .Y(_10_)
);

INVX1 _6713_ (
    .A(_429_),
    .Y(_439_)
);

AOI21X1 _6714_ (
    .A(_435_),
    .B(_433_),
    .C(_436_),
    .Y(_440_)
);

OAI21X1 _6715_ (
    .A(_421_),
    .B(_423_),
    .C(_253__bF$buf5),
    .Y(_441_)
);

INVX1 _6716_ (
    .A(_441_),
    .Y(_442_)
);

NAND2X1 _6717_ (
    .A(\genblk1[0].u_ce.Yin12b [11]),
    .B(_312_),
    .Y(_443_)
);

INVX1 _6718_ (
    .A(\genblk1[0].u_ce.Yin12b [11]),
    .Y(_444_)
);

NAND2X1 _6719_ (
    .A(\genblk1[0].u_ce.Xin12b [11]),
    .B(_444_),
    .Y(_445_)
);

NAND2X1 _6720_ (
    .A(_443_),
    .B(_445_),
    .Y(_446_)
);

OR2X2 _6721_ (
    .A(_442_),
    .B(_446_),
    .Y(_447_)
);

NAND2X1 _6722_ (
    .A(_446_),
    .B(_442_),
    .Y(_448_)
);

NAND2X1 _6723_ (
    .A(_448_),
    .B(_447_),
    .Y(_449_)
);

OAI21X1 _6724_ (
    .A(_439_),
    .B(_440_),
    .C(_449_),
    .Y(_450_)
);

INVX1 _6725_ (
    .A(_449_),
    .Y(_451_)
);

NAND3X1 _6726_ (
    .A(_429_),
    .B(_451_),
    .C(_431_),
    .Y(_452_)
);

NAND3X1 _6727_ (
    .A(_162_),
    .B(_452_),
    .C(_450_),
    .Y(_453_)
);

AOI22X1 _6728_ (
    .A(_125_),
    .B(_158__bF$buf3),
    .C(_453_),
    .D(_282_),
    .Y(_11_)
);

INVX1 _6729_ (
    .A(\genblk1[0].u_ce.Ycalc [0]),
    .Y(_454_)
);

OAI21X1 _6730_ (
    .A(1'h0),
    .B(_373_),
    .C(\genblk1[0].u_ce.Vld_bF$buf3 ),
    .Y(_455_)
);

INVX2 _6731_ (
    .A(_455_),
    .Y(_456_)
);

INVX1 _6732_ (
    .A(\genblk1[0].u_ce.Yin0 [0]),
    .Y(_457_)
);

AOI21X1 _6733_ (
    .A(_224_),
    .B(_231_),
    .C(_457_),
    .Y(_458_)
);

OAI21X1 _6734_ (
    .A(_458_),
    .B(_184_),
    .C(_456_),
    .Y(_459_)
);

OAI21X1 _6735_ (
    .A(_454_),
    .B(\genblk1[0].u_ce.Vld_bF$buf2 ),
    .C(_459_),
    .Y(_12_)
);

NAND2X1 _6736_ (
    .A(\genblk1[0].u_ce.Ycalc [1]),
    .B(_158__bF$buf2),
    .Y(_460_)
);

NAND3X1 _6737_ (
    .A(_246_),
    .B(_183_),
    .C(_247_),
    .Y(_461_)
);

OAI21X1 _6738_ (
    .A(_245_),
    .B(_185_),
    .C(_184_),
    .Y(_462_)
);

AOI21X1 _6739_ (
    .A(_462_),
    .B(_461_),
    .C(_163_),
    .Y(_463_)
);

OAI21X1 _6740_ (
    .A(_158__bF$buf1),
    .B(_463_),
    .C(_460_),
    .Y(_13_)
);

NAND2X1 _6741_ (
    .A(\genblk1[0].u_ce.Xcalc [0]),
    .B(_158__bF$buf0),
    .Y(_464_)
);

MUX2X1 _6742_ (
    .A(\genblk1[0].u_ce.Yin12b [7]),
    .B(\genblk1[0].u_ce.Yin12b [6]),
    .S(1'h0),
    .Y(_465_)
);

NAND2X1 _6743_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin12b [5]),
    .Y(_466_)
);

OAI21X1 _6744_ (
    .A(1'h0),
    .B(_285_),
    .C(_466_),
    .Y(_467_)
);

NAND2X1 _6745_ (
    .A(_164__bF$buf4),
    .B(_467_),
    .Y(_468_)
);

OAI21X1 _6746_ (
    .A(_164__bF$buf3),
    .B(_465_),
    .C(_468_),
    .Y(_469_)
);

NAND2X1 _6747_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin1 [1]),
    .Y(_470_)
);

OAI21X1 _6748_ (
    .A(1'h0),
    .B(_187_),
    .C(_470_),
    .Y(_471_)
);

NAND2X1 _6749_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin0 [1]),
    .Y(_472_)
);

OAI21X1 _6750_ (
    .A(1'h0),
    .B(_457_),
    .C(_472_),
    .Y(_473_)
);

MUX2X1 _6751_ (
    .A(_473_),
    .B(_471_),
    .S(_164__bF$buf2),
    .Y(_474_)
);

NAND2X1 _6752_ (
    .A(_191__bF$buf2),
    .B(_474_),
    .Y(_475_)
);

OAI21X1 _6753_ (
    .A(_191__bF$buf1),
    .B(_469_),
    .C(_475_),
    .Y(_476_)
);

INVX1 _6754_ (
    .A(_476_),
    .Y(_477_)
);

NOR2X1 _6755_ (
    .A(\genblk1[0].u_ce.Xin0 [0]),
    .B(_477_),
    .Y(_478_)
);

OAI21X1 _6756_ (
    .A(_220_),
    .B(_476_),
    .C(_456_),
    .Y(_479_)
);

OAI21X1 _6757_ (
    .A(_479_),
    .B(_478_),
    .C(_464_),
    .Y(_14_)
);

NAND2X1 _6758_ (
    .A(\genblk1[0].u_ce.Xcalc [1]),
    .B(_158__bF$buf4),
    .Y(_480_)
);

NOR2X1 _6759_ (
    .A(_220_),
    .B(_476_),
    .Y(_481_)
);

NAND2X1 _6760_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin12b [4]),
    .Y(_482_)
);

OAI21X1 _6761_ (
    .A(1'h0),
    .B(_275_),
    .C(_482_),
    .Y(_483_)
);

NAND2X1 _6762_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin1 [0]),
    .Y(_484_)
);

OAI21X1 _6763_ (
    .A(1'h0),
    .B(_242_),
    .C(_484_),
    .Y(_485_)
);

MUX2X1 _6764_ (
    .A(_485_),
    .B(_483_),
    .S(_164__bF$buf1),
    .Y(_486_)
);

NAND2X1 _6765_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin12b [8]),
    .Y(_487_)
);

OAI21X1 _6766_ (
    .A(1'h0),
    .B(_359_),
    .C(_487_),
    .Y(_488_)
);

NAND2X1 _6767_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin12b [6]),
    .Y(_489_)
);

OAI21X1 _6768_ (
    .A(1'h0),
    .B(_310_),
    .C(_489_),
    .Y(_490_)
);

MUX2X1 _6769_ (
    .A(_490_),
    .B(_488_),
    .S(_164__bF$buf0),
    .Y(_491_)
);

MUX2X1 _6770_ (
    .A(_491_),
    .B(_486_),
    .S(1'h0),
    .Y(_492_)
);

NOR2X1 _6771_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf4 ),
    .B(_476_),
    .Y(_493_)
);

NAND2X1 _6772_ (
    .A(_492_),
    .B(_493_),
    .Y(_494_)
);

NAND2X1 _6773_ (
    .A(_191__bF$buf0),
    .B(_486_),
    .Y(_495_)
);

NAND2X1 _6774_ (
    .A(1'h0),
    .B(_491_),
    .Y(_496_)
);

NAND2X1 _6775_ (
    .A(_495_),
    .B(_496_),
    .Y(_497_)
);

OAI21X1 _6776_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .B(_476_),
    .C(_497_),
    .Y(_498_)
);

NAND3X1 _6777_ (
    .A(\genblk1[0].u_ce.Xin0 [1]),
    .B(_498_),
    .C(_494_),
    .Y(_499_)
);

OAI21X1 _6778_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_476_),
    .C(_492_),
    .Y(_500_)
);

NAND2X1 _6779_ (
    .A(_497_),
    .B(_493_),
    .Y(_501_)
);

NAND3X1 _6780_ (
    .A(_200_),
    .B(_500_),
    .C(_501_),
    .Y(_502_)
);

NAND3X1 _6781_ (
    .A(_481_),
    .B(_499_),
    .C(_502_),
    .Y(_503_)
);

INVX1 _6782_ (
    .A(_481_),
    .Y(_504_)
);

AOI21X1 _6783_ (
    .A(_501_),
    .B(_500_),
    .C(_200_),
    .Y(_505_)
);

AOI21X1 _6784_ (
    .A(_494_),
    .B(_498_),
    .C(\genblk1[0].u_ce.Xin0 [1]),
    .Y(_506_)
);

OAI21X1 _6785_ (
    .A(_505_),
    .B(_506_),
    .C(_504_),
    .Y(_507_)
);

AOI21X1 _6786_ (
    .A(_507_),
    .B(_503_),
    .C(_163_),
    .Y(_508_)
);

OAI21X1 _6787_ (
    .A(_158__bF$buf3),
    .B(_508_),
    .C(_480_),
    .Y(_15_)
);

OAI21X1 _6788_ (
    .A(_504_),
    .B(_506_),
    .C(_499_),
    .Y(_509_)
);

MUX2X1 _6789_ (
    .A(\genblk1[0].u_ce.Yin12b [9]),
    .B(\genblk1[0].u_ce.Yin12b [8]),
    .S(1'h0),
    .Y(_510_)
);

MUX2X1 _6790_ (
    .A(_510_),
    .B(_465_),
    .S(1'h0),
    .Y(_511_)
);

NOR2X1 _6791_ (
    .A(1'h0),
    .B(_164__bF$buf4),
    .Y(_512_)
);

NAND2X1 _6792_ (
    .A(_467_),
    .B(_512_),
    .Y(_513_)
);

NAND2X1 _6793_ (
    .A(_161_),
    .B(_471_),
    .Y(_514_)
);

NAND2X1 _6794_ (
    .A(_514_),
    .B(_513_),
    .Y(_515_)
);

AOI21X1 _6795_ (
    .A(1'h0),
    .B(_511_),
    .C(_515_),
    .Y(_516_)
);

NAND2X1 _6796_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin12b [7]),
    .Y(_517_)
);

OAI21X1 _6797_ (
    .A(1'h0),
    .B(_334_),
    .C(_517_),
    .Y(_518_)
);

MUX2X1 _6798_ (
    .A(_467_),
    .B(_518_),
    .S(_164__bF$buf3),
    .Y(_519_)
);

NAND2X1 _6799_ (
    .A(1'h0),
    .B(_519_),
    .Y(_520_)
);

AOI21X1 _6800_ (
    .A(_475_),
    .B(_520_),
    .C(_492_),
    .Y(_521_)
);

NOR2X1 _6801_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .B(_521_),
    .Y(_522_)
);

NAND2X1 _6802_ (
    .A(_516_),
    .B(_522_),
    .Y(_523_)
);

INVX1 _6803_ (
    .A(_516_),
    .Y(_524_)
);

OAI21X1 _6804_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .B(_521_),
    .C(_524_),
    .Y(_525_)
);

AOI21X1 _6805_ (
    .A(_523_),
    .B(_525_),
    .C(_216_),
    .Y(_526_)
);

NAND3X1 _6806_ (
    .A(_216_),
    .B(_525_),
    .C(_523_),
    .Y(_527_)
);

INVX1 _6807_ (
    .A(_527_),
    .Y(_528_)
);

NOR2X1 _6808_ (
    .A(_526_),
    .B(_528_),
    .Y(_529_)
);

NOR2X1 _6809_ (
    .A(_509_),
    .B(_529_),
    .Y(_530_)
);

AOI21X1 _6810_ (
    .A(_481_),
    .B(_502_),
    .C(_505_),
    .Y(_531_)
);

INVX1 _6811_ (
    .A(_529_),
    .Y(_532_)
);

OAI21X1 _6812_ (
    .A(_531_),
    .B(_532_),
    .C(_456_),
    .Y(_533_)
);

OAI22X1 _6813_ (
    .A(_133_),
    .B(\genblk1[0].u_ce.Vld_bF$buf1 ),
    .C(_530_),
    .D(_533_),
    .Y(_16_)
);

NAND2X1 _6814_ (
    .A(\genblk1[0].u_ce.Xcalc [3]),
    .B(_158__bF$buf2),
    .Y(_534_)
);

AOI21X1 _6815_ (
    .A(_509_),
    .B(_527_),
    .C(_526_),
    .Y(_535_)
);

NAND2X1 _6816_ (
    .A(1'h0),
    .B(_420_),
    .Y(_536_)
);

OAI21X1 _6817_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin12b [9]),
    .C(_536_),
    .Y(_537_)
);

NAND2X1 _6818_ (
    .A(_164__bF$buf2),
    .B(_488_),
    .Y(_538_)
);

OAI21X1 _6819_ (
    .A(_164__bF$buf1),
    .B(_537_),
    .C(_538_),
    .Y(_539_)
);

NAND2X1 _6820_ (
    .A(_490_),
    .B(_512_),
    .Y(_540_)
);

NAND2X1 _6821_ (
    .A(_161_),
    .B(_483_),
    .Y(_541_)
);

NAND2X1 _6822_ (
    .A(_541_),
    .B(_540_),
    .Y(_542_)
);

AOI21X1 _6823_ (
    .A(_539_),
    .B(1'h0),
    .C(_542_),
    .Y(_543_)
);

NAND3X1 _6824_ (
    .A(_516_),
    .B(_497_),
    .C(_476_),
    .Y(_544_)
);

NAND2X1 _6825_ (
    .A(_253__bF$buf4),
    .B(_544_),
    .Y(_545_)
);

OR2X2 _6826_ (
    .A(_545_),
    .B(_543_),
    .Y(_546_)
);

INVX1 _6827_ (
    .A(_544_),
    .Y(_547_)
);

OAI21X1 _6828_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf4 ),
    .B(_547_),
    .C(_543_),
    .Y(_548_)
);

NAND3X1 _6829_ (
    .A(\genblk1[0].u_ce.Xin1 [1]),
    .B(_548_),
    .C(_546_),
    .Y(_549_)
);

INVX1 _6830_ (
    .A(_543_),
    .Y(_550_)
);

OR2X2 _6831_ (
    .A(_545_),
    .B(_550_),
    .Y(_551_)
);

OAI21X1 _6832_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .B(_547_),
    .C(_550_),
    .Y(_552_)
);

NAND3X1 _6833_ (
    .A(_195_),
    .B(_552_),
    .C(_551_),
    .Y(_553_)
);

NAND2X1 _6834_ (
    .A(_549_),
    .B(_553_),
    .Y(_554_)
);

OR2X2 _6835_ (
    .A(_535_),
    .B(_554_),
    .Y(_555_)
);

NAND2X1 _6836_ (
    .A(_554_),
    .B(_535_),
    .Y(_556_)
);

AOI21X1 _6837_ (
    .A(_555_),
    .B(_556_),
    .C(_163_),
    .Y(_557_)
);

OAI21X1 _6838_ (
    .A(_158__bF$buf1),
    .B(_557_),
    .C(_534_),
    .Y(_17_)
);

OAI21X1 _6839_ (
    .A(_554_),
    .B(_535_),
    .C(_549_),
    .Y(_558_)
);

NAND2X1 _6840_ (
    .A(1'h0),
    .B(\genblk1[0].u_ce.Yin12b [11]),
    .Y(_559_)
);

OAI21X1 _6841_ (
    .A(1'h0),
    .B(_420_),
    .C(_559_),
    .Y(_560_)
);

NAND2X1 _6842_ (
    .A(1'h0),
    .B(_560_),
    .Y(_561_)
);

OAI21X1 _6843_ (
    .A(1'h0),
    .B(_510_),
    .C(_561_),
    .Y(_562_)
);

NAND2X1 _6844_ (
    .A(1'h0),
    .B(_562_),
    .Y(_563_)
);

OAI21X1 _6845_ (
    .A(1'h0),
    .B(_519_),
    .C(_563_),
    .Y(_564_)
);

INVX1 _6846_ (
    .A(_564_),
    .Y(_565_)
);

OAI21X1 _6847_ (
    .A(_550_),
    .B(_544_),
    .C(_253__bF$buf3),
    .Y(_566_)
);

OR2X2 _6848_ (
    .A(_566_),
    .B(_565_),
    .Y(_567_)
);

NAND2X1 _6849_ (
    .A(_565_),
    .B(_566_),
    .Y(_568_)
);

NAND3X1 _6850_ (
    .A(\genblk1[0].u_ce.Xin12b [4]),
    .B(_568_),
    .C(_567_),
    .Y(_569_)
);

OR2X2 _6851_ (
    .A(_566_),
    .B(_564_),
    .Y(_570_)
);

NAND2X1 _6852_ (
    .A(_564_),
    .B(_566_),
    .Y(_571_)
);

NAND3X1 _6853_ (
    .A(_197_),
    .B(_571_),
    .C(_570_),
    .Y(_572_)
);

AND2X2 _6854_ (
    .A(_569_),
    .B(_572_),
    .Y(_573_)
);

NAND2X1 _6855_ (
    .A(_573_),
    .B(_558_),
    .Y(_574_)
);

INVX1 _6856_ (
    .A(_526_),
    .Y(_575_)
);

OAI21X1 _6857_ (
    .A(_528_),
    .B(_531_),
    .C(_575_),
    .Y(_576_)
);

INVX1 _6858_ (
    .A(_549_),
    .Y(_577_)
);

AOI21X1 _6859_ (
    .A(_576_),
    .B(_553_),
    .C(_577_),
    .Y(_578_)
);

NAND2X1 _6860_ (
    .A(_572_),
    .B(_569_),
    .Y(_579_)
);

NAND2X1 _6861_ (
    .A(_579_),
    .B(_578_),
    .Y(_580_)
);

NAND2X1 _6862_ (
    .A(_574_),
    .B(_580_),
    .Y(_581_)
);

AOI22X1 _6863_ (
    .A(_135_),
    .B(_158__bF$buf0),
    .C(_581_),
    .D(_456_),
    .Y(_18_)
);

NAND3X1 _6864_ (
    .A(_543_),
    .B(_565_),
    .C(_547_),
    .Y(_582_)
);

NOR2X1 _6865_ (
    .A(1'h0),
    .B(_537_),
    .Y(_583_)
);

NOR2X1 _6866_ (
    .A(_164__bF$buf0),
    .B(_444_),
    .Y(_584_)
);

OAI21X1 _6867_ (
    .A(_584_),
    .B(_583_),
    .C(1'h0),
    .Y(_585_)
);

OAI21X1 _6868_ (
    .A(1'h0),
    .B(_491_),
    .C(_585_),
    .Y(_586_)
);

NAND3X1 _6869_ (
    .A(_253__bF$buf2),
    .B(_586_),
    .C(_582_),
    .Y(_587_)
);

INVX1 _6870_ (
    .A(_586_),
    .Y(_588_)
);

NAND3X1 _6871_ (
    .A(_516_),
    .B(_543_),
    .C(_521_),
    .Y(_589_)
);

OAI21X1 _6872_ (
    .A(_564_),
    .B(_589_),
    .C(_253__bF$buf1),
    .Y(_590_)
);

NAND2X1 _6873_ (
    .A(_588_),
    .B(_590_),
    .Y(_591_)
);

NAND3X1 _6874_ (
    .A(\genblk1[0].u_ce.Xin12b [5]),
    .B(_591_),
    .C(_587_),
    .Y(_592_)
);

NAND3X1 _6875_ (
    .A(_253__bF$buf0),
    .B(_588_),
    .C(_582_),
    .Y(_593_)
);

NAND2X1 _6876_ (
    .A(_586_),
    .B(_590_),
    .Y(_594_)
);

NAND3X1 _6877_ (
    .A(_205_),
    .B(_594_),
    .C(_593_),
    .Y(_595_)
);

NAND2X1 _6878_ (
    .A(_592_),
    .B(_595_),
    .Y(_596_)
);

AOI21X1 _6879_ (
    .A(_574_),
    .B(_569_),
    .C(_596_),
    .Y(_597_)
);

OAI21X1 _6880_ (
    .A(_579_),
    .B(_578_),
    .C(_569_),
    .Y(_598_)
);

AND2X2 _6881_ (
    .A(_592_),
    .B(_595_),
    .Y(_599_)
);

OAI21X1 _6882_ (
    .A(_599_),
    .B(_598_),
    .C(_456_),
    .Y(_600_)
);

OAI22X1 _6883_ (
    .A(_150_),
    .B(\genblk1[0].u_ce.Vld_bF$buf0 ),
    .C(_597_),
    .D(_600_),
    .Y(_19_)
);

NOR2X1 _6884_ (
    .A(_564_),
    .B(_589_),
    .Y(_601_)
);

NAND2X1 _6885_ (
    .A(_588_),
    .B(_601_),
    .Y(_602_)
);

AOI21X1 _6886_ (
    .A(_164__bF$buf4),
    .B(_560_),
    .C(_584_),
    .Y(_603_)
);

NAND2X1 _6887_ (
    .A(_191__bF$buf3),
    .B(_511_),
    .Y(_604_)
);

OAI21X1 _6888_ (
    .A(_191__bF$buf2),
    .B(_603_),
    .C(_604_),
    .Y(_605_)
);

NAND3X1 _6889_ (
    .A(_253__bF$buf5),
    .B(_605_),
    .C(_602_),
    .Y(_606_)
);

NOR3X1 _6890_ (
    .A(_564_),
    .B(_586_),
    .C(_589_),
    .Y(_607_)
);

INVX1 _6891_ (
    .A(_605_),
    .Y(_608_)
);

OAI21X1 _6892_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_607_),
    .C(_608_),
    .Y(_609_)
);

NAND3X1 _6893_ (
    .A(\genblk1[0].u_ce.Xin12b [6]),
    .B(_609_),
    .C(_606_),
    .Y(_610_)
);

NAND3X1 _6894_ (
    .A(_253__bF$buf4),
    .B(_608_),
    .C(_602_),
    .Y(_611_)
);

OAI21X1 _6895_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .B(_607_),
    .C(_605_),
    .Y(_612_)
);

NAND3X1 _6896_ (
    .A(_207_),
    .B(_612_),
    .C(_611_),
    .Y(_613_)
);

AND2X2 _6897_ (
    .A(_610_),
    .B(_613_),
    .Y(_614_)
);

NAND2X1 _6898_ (
    .A(_573_),
    .B(_599_),
    .Y(_615_)
);

INVX1 _6899_ (
    .A(_569_),
    .Y(_616_)
);

INVX1 _6900_ (
    .A(_592_),
    .Y(_617_)
);

AOI21X1 _6901_ (
    .A(_616_),
    .B(_595_),
    .C(_617_),
    .Y(_618_)
);

OAI21X1 _6902_ (
    .A(_578_),
    .B(_615_),
    .C(_618_),
    .Y(_619_)
);

AND2X2 _6903_ (
    .A(_619_),
    .B(_614_),
    .Y(_620_)
);

NOR2X1 _6904_ (
    .A(_614_),
    .B(_619_),
    .Y(_621_)
);

OAI21X1 _6905_ (
    .A(_621_),
    .B(_620_),
    .C(_162_),
    .Y(_622_)
);

NAND2X1 _6906_ (
    .A(\genblk1[0].u_ce.Vld_bF$buf4 ),
    .B(_622_),
    .Y(_623_)
);

OAI21X1 _6907_ (
    .A(_136_),
    .B(\genblk1[0].u_ce.Vld_bF$buf3 ),
    .C(_623_),
    .Y(_20_)
);

INVX1 _6908_ (
    .A(_610_),
    .Y(_624_)
);

NOR2X1 _6909_ (
    .A(_624_),
    .B(_620_),
    .Y(_625_)
);

NAND2X1 _6910_ (
    .A(_608_),
    .B(_607_),
    .Y(_626_)
);

NOR2X1 _6911_ (
    .A(_191__bF$buf1),
    .B(_444_),
    .Y(_627_)
);

AOI21X1 _6912_ (
    .A(_539_),
    .B(_191__bF$buf0),
    .C(_627_),
    .Y(_628_)
);

NAND3X1 _6913_ (
    .A(_253__bF$buf3),
    .B(_628_),
    .C(_626_),
    .Y(_629_)
);

INVX1 _6914_ (
    .A(_629_),
    .Y(_630_)
);

AOI21X1 _6915_ (
    .A(_626_),
    .B(_253__bF$buf2),
    .C(_628_),
    .Y(_631_)
);

OAI21X1 _6916_ (
    .A(_631_),
    .B(_630_),
    .C(\genblk1[0].u_ce.Xin12b [7]),
    .Y(_632_)
);

INVX1 _6917_ (
    .A(_631_),
    .Y(_633_)
);

NAND3X1 _6918_ (
    .A(_210_),
    .B(_629_),
    .C(_633_),
    .Y(_634_)
);

AND2X2 _6919_ (
    .A(_634_),
    .B(_632_),
    .Y(_635_)
);

OR2X2 _6920_ (
    .A(_625_),
    .B(_635_),
    .Y(_636_)
);

AOI21X1 _6921_ (
    .A(_625_),
    .B(_635_),
    .C(_455_),
    .Y(_637_)
);

AOI22X1 _6922_ (
    .A(_149_),
    .B(_158__bF$buf4),
    .C(_636_),
    .D(_637_),
    .Y(_21_)
);

NOR2X1 _6923_ (
    .A(_579_),
    .B(_596_),
    .Y(_638_)
);

OAI21X1 _6924_ (
    .A(_569_),
    .B(_596_),
    .C(_592_),
    .Y(_639_)
);

AOI21X1 _6925_ (
    .A(_638_),
    .B(_558_),
    .C(_639_),
    .Y(_640_)
);

AOI21X1 _6926_ (
    .A(_633_),
    .B(_629_),
    .C(_210_),
    .Y(_641_)
);

AOI21X1 _6927_ (
    .A(_624_),
    .B(_634_),
    .C(_641_),
    .Y(_642_)
);

NAND3X1 _6928_ (
    .A(_614_),
    .B(_632_),
    .C(_634_),
    .Y(_643_)
);

OAI21X1 _6929_ (
    .A(_643_),
    .B(_640_),
    .C(_642_),
    .Y(_644_)
);

NAND3X1 _6930_ (
    .A(_608_),
    .B(_628_),
    .C(_607_),
    .Y(_645_)
);

INVX1 _6931_ (
    .A(_562_),
    .Y(_646_)
);

INVX1 _6932_ (
    .A(_627_),
    .Y(_647_)
);

OAI21X1 _6933_ (
    .A(1'h0),
    .B(_646_),
    .C(_647_),
    .Y(_648_)
);

INVX1 _6934_ (
    .A(_648_),
    .Y(_649_)
);

NAND3X1 _6935_ (
    .A(_253__bF$buf1),
    .B(_649_),
    .C(_645_),
    .Y(_650_)
);

INVX1 _6936_ (
    .A(_650_),
    .Y(_651_)
);

AOI21X1 _6937_ (
    .A(_645_),
    .B(_253__bF$buf0),
    .C(_649_),
    .Y(_652_)
);

OAI21X1 _6938_ (
    .A(_652_),
    .B(_651_),
    .C(\genblk1[0].u_ce.Xin12b [8]),
    .Y(_653_)
);

INVX1 _6939_ (
    .A(_652_),
    .Y(_654_)
);

NAND3X1 _6940_ (
    .A(_212_),
    .B(_650_),
    .C(_654_),
    .Y(_655_)
);

AND2X2 _6941_ (
    .A(_655_),
    .B(_653_),
    .Y(_656_)
);

OR2X2 _6942_ (
    .A(_644_),
    .B(_656_),
    .Y(_657_)
);

INVX1 _6943_ (
    .A(_657_),
    .Y(_658_)
);

NAND2X1 _6944_ (
    .A(_656_),
    .B(_644_),
    .Y(_659_)
);

NAND2X1 _6945_ (
    .A(_456_),
    .B(_659_),
    .Y(_660_)
);

OAI22X1 _6946_ (
    .A(_138_),
    .B(\genblk1[0].u_ce.Vld_bF$buf2 ),
    .C(_660_),
    .D(_658_),
    .Y(_22_)
);

NOR3X1 _6947_ (
    .A(_586_),
    .B(_605_),
    .C(_582_),
    .Y(_661_)
);

NAND3X1 _6948_ (
    .A(_628_),
    .B(_649_),
    .C(_661_),
    .Y(_662_)
);

OR2X2 _6949_ (
    .A(_583_),
    .B(_584_),
    .Y(_663_)
);

AOI21X1 _6950_ (
    .A(_663_),
    .B(_191__bF$buf3),
    .C(_627_),
    .Y(_664_)
);

INVX1 _6951_ (
    .A(_664_),
    .Y(_665_)
);

NAND3X1 _6952_ (
    .A(_253__bF$buf5),
    .B(_665_),
    .C(_662_),
    .Y(_666_)
);

OAI21X1 _6953_ (
    .A(_648_),
    .B(_645_),
    .C(_253__bF$buf4),
    .Y(_667_)
);

NAND2X1 _6954_ (
    .A(_664_),
    .B(_667_),
    .Y(_668_)
);

NAND3X1 _6955_ (
    .A(\genblk1[0].u_ce.Xin12b [9]),
    .B(_668_),
    .C(_666_),
    .Y(_669_)
);

NAND3X1 _6956_ (
    .A(_253__bF$buf3),
    .B(_664_),
    .C(_662_),
    .Y(_670_)
);

NAND2X1 _6957_ (
    .A(_665_),
    .B(_667_),
    .Y(_671_)
);

NAND3X1 _6958_ (
    .A(_257_),
    .B(_671_),
    .C(_670_),
    .Y(_672_)
);

NAND2X1 _6959_ (
    .A(_669_),
    .B(_672_),
    .Y(_673_)
);

AOI21X1 _6960_ (
    .A(_659_),
    .B(_653_),
    .C(_673_),
    .Y(_674_)
);

NAND3X1 _6961_ (
    .A(_653_),
    .B(_673_),
    .C(_659_),
    .Y(_675_)
);

NAND2X1 _6962_ (
    .A(_456_),
    .B(_675_),
    .Y(_676_)
);

OAI22X1 _6963_ (
    .A(_146_),
    .B(\genblk1[0].u_ce.Vld_bF$buf1 ),
    .C(_674_),
    .D(_676_),
    .Y(_23_)
);

NAND2X1 _6964_ (
    .A(\genblk1[0].u_ce.Xcalc [10]),
    .B(_158__bF$buf3),
    .Y(_677_)
);

OAI21X1 _6965_ (
    .A(1'h0),
    .B(_603_),
    .C(_647_),
    .Y(_678_)
);

OAI21X1 _6966_ (
    .A(_665_),
    .B(_662_),
    .C(_253__bF$buf2),
    .Y(_679_)
);

NOR2X1 _6967_ (
    .A(_678_),
    .B(_679_),
    .Y(_680_)
);

NAND2X1 _6968_ (
    .A(_678_),
    .B(_679_),
    .Y(_681_)
);

INVX1 _6969_ (
    .A(_681_),
    .Y(_682_)
);

OAI21X1 _6970_ (
    .A(_680_),
    .B(_682_),
    .C(\genblk1[0].u_ce.Xin12b [10]),
    .Y(_683_)
);

INVX1 _6971_ (
    .A(_680_),
    .Y(_684_)
);

NAND3X1 _6972_ (
    .A(_287_),
    .B(_681_),
    .C(_684_),
    .Y(_685_)
);

AND2X2 _6973_ (
    .A(_685_),
    .B(_683_),
    .Y(_686_)
);

OAI21X1 _6974_ (
    .A(_653_),
    .B(_673_),
    .C(_669_),
    .Y(_687_)
);

NAND3X1 _6975_ (
    .A(_614_),
    .B(_619_),
    .C(_635_),
    .Y(_688_)
);

NAND3X1 _6976_ (
    .A(_669_),
    .B(_672_),
    .C(_656_),
    .Y(_689_)
);

AOI21X1 _6977_ (
    .A(_688_),
    .B(_642_),
    .C(_689_),
    .Y(_690_)
);

OAI21X1 _6978_ (
    .A(_687_),
    .B(_690_),
    .C(_686_),
    .Y(_691_)
);

NAND2X1 _6979_ (
    .A(_683_),
    .B(_685_),
    .Y(_692_)
);

NAND2X1 _6980_ (
    .A(_653_),
    .B(_655_),
    .Y(_693_)
);

NOR2X1 _6981_ (
    .A(_693_),
    .B(_673_),
    .Y(_694_)
);

AOI21X1 _6982_ (
    .A(_644_),
    .B(_694_),
    .C(_687_),
    .Y(_695_)
);

NAND2X1 _6983_ (
    .A(_692_),
    .B(_695_),
    .Y(_696_)
);

AOI21X1 _6984_ (
    .A(_691_),
    .B(_696_),
    .C(_163_),
    .Y(_697_)
);

OAI21X1 _6985_ (
    .A(_158__bF$buf2),
    .B(_697_),
    .C(_677_),
    .Y(_24_)
);

NAND2X1 _6986_ (
    .A(\genblk1[0].u_ce.Xcalc [11]),
    .B(_158__bF$buf1),
    .Y(_698_)
);

OR2X2 _6987_ (
    .A(_662_),
    .B(_665_),
    .Y(_699_)
);

OAI21X1 _6988_ (
    .A(_678_),
    .B(_699_),
    .C(_253__bF$buf1),
    .Y(_700_)
);

OR2X2 _6989_ (
    .A(_700_),
    .B(_446_),
    .Y(_701_)
);

NAND2X1 _6990_ (
    .A(_446_),
    .B(_700_),
    .Y(_702_)
);

AOI22X1 _6991_ (
    .A(_701_),
    .B(_702_),
    .C(_691_),
    .D(_683_),
    .Y(_703_)
);

OAI21X1 _6992_ (
    .A(_692_),
    .B(_695_),
    .C(_683_),
    .Y(_704_)
);

NAND2X1 _6993_ (
    .A(_702_),
    .B(_701_),
    .Y(_705_)
);

OAI21X1 _6994_ (
    .A(_705_),
    .B(_704_),
    .C(_456_),
    .Y(_706_)
);

OAI21X1 _6995_ (
    .A(_703_),
    .B(_706_),
    .C(_698_),
    .Y(_25_)
);

NAND2X1 _6996_ (
    .A(1'h0),
    .B(1'h0),
    .Y(_707_)
);

OAI21X1 _6997_ (
    .A(_191__bF$buf2),
    .B(_373_),
    .C(_707_),
    .Y(_708_)
);

NOR2X1 _6998_ (
    .A(_154_),
    .B(_708_),
    .Y(_709_)
);

AND2X2 _6999_ (
    .A(_708_),
    .B(_154_),
    .Y(_710_)
);

OR2X2 _7000_ (
    .A(_710_),
    .B(_709_),
    .Y(_711_)
);

NAND2X1 _7001_ (
    .A(\genblk1[0].u_ce.Acalc [0]),
    .B(_158__bF$buf0),
    .Y(_712_)
);

OAI21X1 _7002_ (
    .A(_158__bF$buf4),
    .B(_711_),
    .C(_712_),
    .Y(_26_)
);

NAND2X1 _7003_ (
    .A(\genblk1[0].u_ce.Acalc [1]),
    .B(_158__bF$buf3),
    .Y(_713_)
);

OAI21X1 _7004_ (
    .A(1'h0),
    .B(_160_),
    .C(1'h0),
    .Y(_714_)
);

OAI21X1 _7005_ (
    .A(1'h0),
    .B(_160_),
    .C(_714_),
    .Y(_715_)
);

OAI21X1 _7006_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .B(_708_),
    .C(_715_),
    .Y(_716_)
);

OAI21X1 _7007_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf4 ),
    .B(_715_),
    .C(_716_),
    .Y(_717_)
);

OR2X2 _7008_ (
    .A(_717_),
    .B(\genblk1[0].u_ce.Ain0 [1]),
    .Y(_718_)
);

NAND2X1 _7009_ (
    .A(\genblk1[0].u_ce.Ain0 [1]),
    .B(_717_),
    .Y(_719_)
);

NAND2X1 _7010_ (
    .A(_719_),
    .B(_718_),
    .Y(_720_)
);

NOR2X1 _7011_ (
    .A(_709_),
    .B(_720_),
    .Y(_721_)
);

NAND2X1 _7012_ (
    .A(_709_),
    .B(_720_),
    .Y(_722_)
);

NAND2X1 _7013_ (
    .A(\genblk1[0].u_ce.Vld_bF$buf0 ),
    .B(_722_),
    .Y(_723_)
);

OAI21X1 _7014_ (
    .A(_721_),
    .B(_723_),
    .C(_713_),
    .Y(_27_)
);

NAND2X1 _7015_ (
    .A(\genblk1[0].u_ce.Acalc [2]),
    .B(_158__bF$buf2),
    .Y(_724_)
);

OAI21X1 _7016_ (
    .A(_156_),
    .B(_717_),
    .C(_722_),
    .Y(_725_)
);

OAI21X1 _7017_ (
    .A(_160_),
    .B(_164__bF$buf3),
    .C(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_726_)
);

NAND3X1 _7018_ (
    .A(1'h0),
    .B(_373_),
    .C(_726_),
    .Y(_727_)
);

OAI21X1 _7019_ (
    .A(1'h0),
    .B(_726_),
    .C(_727_),
    .Y(_728_)
);

NAND2X1 _7020_ (
    .A(\genblk1[0].u_ce.Ain1 [0]),
    .B(_728_),
    .Y(_729_)
);

OR2X2 _7021_ (
    .A(_728_),
    .B(\genblk1[0].u_ce.Ain1 [0]),
    .Y(_730_)
);

NAND2X1 _7022_ (
    .A(_729_),
    .B(_730_),
    .Y(_731_)
);

INVX1 _7023_ (
    .A(_731_),
    .Y(_732_)
);

NOR2X1 _7024_ (
    .A(_732_),
    .B(_725_),
    .Y(_733_)
);

NAND2X1 _7025_ (
    .A(_732_),
    .B(_725_),
    .Y(_734_)
);

NAND2X1 _7026_ (
    .A(\genblk1[0].u_ce.Vld_bF$buf4 ),
    .B(_734_),
    .Y(_735_)
);

OAI21X1 _7027_ (
    .A(_733_),
    .B(_735_),
    .C(_724_),
    .Y(_28_)
);

NAND2X1 _7028_ (
    .A(_729_),
    .B(_734_),
    .Y(_736_)
);

INVX1 _7029_ (
    .A(_736_),
    .Y(_737_)
);

INVX1 _7030_ (
    .A(\genblk1[0].u_ce.Ain1 [1]),
    .Y(_738_)
);

OAI21X1 _7031_ (
    .A(1'h0),
    .B(_164__bF$buf2),
    .C(1'h0),
    .Y(_739_)
);

NAND2X1 _7032_ (
    .A(_253__bF$buf0),
    .B(_739_),
    .Y(_740_)
);

OAI21X1 _7033_ (
    .A(1'h0),
    .B(1'h0),
    .C(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .Y(_741_)
);

OAI21X1 _7034_ (
    .A(_160_),
    .B(_741_),
    .C(_740_),
    .Y(_742_)
);

NOR2X1 _7035_ (
    .A(_738_),
    .B(_742_),
    .Y(_743_)
);

NAND2X1 _7036_ (
    .A(_738_),
    .B(_742_),
    .Y(_744_)
);

INVX1 _7037_ (
    .A(_744_),
    .Y(_745_)
);

OAI21X1 _7038_ (
    .A(_743_),
    .B(_745_),
    .C(_737_),
    .Y(_746_)
);

INVX1 _7039_ (
    .A(_743_),
    .Y(_747_)
);

NAND3X1 _7040_ (
    .A(_747_),
    .B(_744_),
    .C(_736_),
    .Y(_748_)
);

NAND2X1 _7041_ (
    .A(_748_),
    .B(_746_),
    .Y(_749_)
);

NAND2X1 _7042_ (
    .A(\genblk1[0].u_ce.Acalc [3]),
    .B(_158__bF$buf1),
    .Y(_750_)
);

OAI21X1 _7043_ (
    .A(_158__bF$buf0),
    .B(_749_),
    .C(_750_),
    .Y(_29_)
);

NOR2X1 _7044_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf1 ),
    .B(_715_),
    .Y(_751_)
);

NAND3X1 _7045_ (
    .A(1'h0),
    .B(_191__bF$buf1),
    .C(_164__bF$buf1),
    .Y(_752_)
);

AOI21X1 _7046_ (
    .A(_714_),
    .B(_752_),
    .C(_253__bF$buf5),
    .Y(_753_)
);

NOR2X1 _7047_ (
    .A(_753_),
    .B(_751_),
    .Y(_754_)
);

NAND2X1 _7048_ (
    .A(\genblk1[0].u_ce.Ain12b [4]),
    .B(_754_),
    .Y(_755_)
);

INVX1 _7049_ (
    .A(\genblk1[0].u_ce.Ain12b [4]),
    .Y(_756_)
);

OAI21X1 _7050_ (
    .A(_753_),
    .B(_751_),
    .C(_756_),
    .Y(_757_)
);

NAND2X1 _7051_ (
    .A(_757_),
    .B(_755_),
    .Y(_758_)
);

AOI21X1 _7052_ (
    .A(_736_),
    .B(_744_),
    .C(_743_),
    .Y(_759_)
);

AND2X2 _7053_ (
    .A(_759_),
    .B(_758_),
    .Y(_760_)
);

OAI21X1 _7054_ (
    .A(_758_),
    .B(_759_),
    .C(\genblk1[0].u_ce.Vld_bF$buf3 ),
    .Y(_761_)
);

OAI22X1 _7055_ (
    .A(_97_),
    .B(\genblk1[0].u_ce.Vld_bF$buf2 ),
    .C(_761_),
    .D(_760_),
    .Y(_30_)
);

NAND2X1 _7056_ (
    .A(\genblk1[0].u_ce.Acalc [5]),
    .B(_158__bF$buf4),
    .Y(_762_)
);

OAI21X1 _7057_ (
    .A(_758_),
    .B(_759_),
    .C(_755_),
    .Y(_763_)
);

OAI21X1 _7058_ (
    .A(1'h0),
    .B(1'h0),
    .C(_192_),
    .Y(_764_)
);

NAND2X1 _7059_ (
    .A(_253__bF$buf4),
    .B(_764_),
    .Y(_765_)
);

INVX1 _7060_ (
    .A(_765_),
    .Y(_766_)
);

NOR2X1 _7061_ (
    .A(_253__bF$buf3),
    .B(_764_),
    .Y(_767_)
);

NOR2X1 _7062_ (
    .A(_767_),
    .B(_766_),
    .Y(_768_)
);

NAND2X1 _7063_ (
    .A(\genblk1[0].u_ce.Ain12b [5]),
    .B(_768_),
    .Y(_769_)
);

INVX1 _7064_ (
    .A(\genblk1[0].u_ce.Ain12b [5]),
    .Y(_770_)
);

OAI21X1 _7065_ (
    .A(_767_),
    .B(_766_),
    .C(_770_),
    .Y(_771_)
);

NAND2X1 _7066_ (
    .A(_771_),
    .B(_769_),
    .Y(_772_)
);

INVX1 _7067_ (
    .A(_772_),
    .Y(_773_)
);

NOR2X1 _7068_ (
    .A(_773_),
    .B(_763_),
    .Y(_774_)
);

NAND2X1 _7069_ (
    .A(_773_),
    .B(_763_),
    .Y(_775_)
);

NAND2X1 _7070_ (
    .A(\genblk1[0].u_ce.Vld_bF$buf1 ),
    .B(_775_),
    .Y(_776_)
);

OAI21X1 _7071_ (
    .A(_774_),
    .B(_776_),
    .C(_762_),
    .Y(_31_)
);

NAND2X1 _7072_ (
    .A(\genblk1[0].u_ce.Acalc [6]),
    .B(_158__bF$buf3),
    .Y(_777_)
);

INVX1 _7073_ (
    .A(_759_),
    .Y(_778_)
);

NOR2X1 _7074_ (
    .A(_758_),
    .B(_772_),
    .Y(_779_)
);

OAI21X1 _7075_ (
    .A(_755_),
    .B(_772_),
    .C(_769_),
    .Y(_780_)
);

AOI21X1 _7076_ (
    .A(_778_),
    .B(_779_),
    .C(_780_),
    .Y(_781_)
);

OAI21X1 _7077_ (
    .A(1'h0),
    .B(_707_),
    .C(_162_),
    .Y(_782_)
);

NOR2X1 _7078_ (
    .A(_253__bF$buf2),
    .B(_782_),
    .Y(_783_)
);

NAND2X1 _7079_ (
    .A(_253__bF$buf1),
    .B(_782_),
    .Y(_784_)
);

INVX1 _7080_ (
    .A(_784_),
    .Y(_785_)
);

NOR2X1 _7081_ (
    .A(_783_),
    .B(_785_),
    .Y(_786_)
);

NAND2X1 _7082_ (
    .A(\genblk1[0].u_ce.Ain12b [6]),
    .B(_786_),
    .Y(_787_)
);

OR2X2 _7083_ (
    .A(_786_),
    .B(\genblk1[0].u_ce.Ain12b [6]),
    .Y(_788_)
);

AND2X2 _7084_ (
    .A(_788_),
    .B(_787_),
    .Y(_789_)
);

INVX1 _7085_ (
    .A(_789_),
    .Y(_790_)
);

AND2X2 _7086_ (
    .A(_781_),
    .B(_790_),
    .Y(_791_)
);

OAI21X1 _7087_ (
    .A(_790_),
    .B(_781_),
    .C(\genblk1[0].u_ce.Vld_bF$buf0 ),
    .Y(_792_)
);

OAI21X1 _7088_ (
    .A(_792_),
    .B(_791_),
    .C(_777_),
    .Y(_32_)
);

OAI21X1 _7089_ (
    .A(_790_),
    .B(_781_),
    .C(_787_),
    .Y(_793_)
);

OAI21X1 _7090_ (
    .A(1'h0),
    .B(1'h0),
    .C(\genblk1[0].u_ce.Ain12b_11_bF$buf0 ),
    .Y(_794_)
);

NAND2X1 _7091_ (
    .A(_794_),
    .B(_254_),
    .Y(_795_)
);

INVX1 _7092_ (
    .A(_795_),
    .Y(_796_)
);

NAND2X1 _7093_ (
    .A(\genblk1[0].u_ce.Ain12b [7]),
    .B(_796_),
    .Y(_797_)
);

INVX1 _7094_ (
    .A(_797_),
    .Y(_798_)
);

NOR2X1 _7095_ (
    .A(\genblk1[0].u_ce.Ain12b [7]),
    .B(_796_),
    .Y(_799_)
);

NOR2X1 _7096_ (
    .A(_799_),
    .B(_798_),
    .Y(_800_)
);

INVX1 _7097_ (
    .A(_800_),
    .Y(_801_)
);

OR2X2 _7098_ (
    .A(_793_),
    .B(_801_),
    .Y(_802_)
);

AOI21X1 _7099_ (
    .A(_793_),
    .B(_801_),
    .C(_158__bF$buf2),
    .Y(_803_)
);

AOI22X1 _7100_ (
    .A(_111_),
    .B(_158__bF$buf1),
    .C(_802_),
    .D(_803_),
    .Y(_33_)
);

NAND2X1 _7101_ (
    .A(\genblk1[0].u_ce.Acalc [8]),
    .B(_158__bF$buf0),
    .Y(_804_)
);

OAI21X1 _7102_ (
    .A(_799_),
    .B(_787_),
    .C(_797_),
    .Y(_805_)
);

NAND2X1 _7103_ (
    .A(_800_),
    .B(_789_),
    .Y(_806_)
);

INVX1 _7104_ (
    .A(_806_),
    .Y(_807_)
);

AOI21X1 _7105_ (
    .A(_807_),
    .B(_780_),
    .C(_805_),
    .Y(_808_)
);

NAND2X1 _7106_ (
    .A(_779_),
    .B(_807_),
    .Y(_809_)
);

OAI21X1 _7107_ (
    .A(_809_),
    .B(_759_),
    .C(_808_),
    .Y(_810_)
);

INVX1 _7108_ (
    .A(\genblk1[0].u_ce.Ain12b [8]),
    .Y(_811_)
);

NAND2X1 _7109_ (
    .A(_253__bF$buf0),
    .B(_161_),
    .Y(_812_)
);

NAND2X1 _7110_ (
    .A(_741_),
    .B(_812_),
    .Y(_813_)
);

OR2X2 _7111_ (
    .A(_813_),
    .B(_811_),
    .Y(_814_)
);

NAND2X1 _7112_ (
    .A(_811_),
    .B(_813_),
    .Y(_815_)
);

AND2X2 _7113_ (
    .A(_814_),
    .B(_815_),
    .Y(_816_)
);

NOR2X1 _7114_ (
    .A(_816_),
    .B(_810_),
    .Y(_817_)
);

NAND2X1 _7115_ (
    .A(_816_),
    .B(_810_),
    .Y(_818_)
);

NAND2X1 _7116_ (
    .A(\genblk1[0].u_ce.Vld_bF$buf4 ),
    .B(_818_),
    .Y(_819_)
);

OAI21X1 _7117_ (
    .A(_817_),
    .B(_819_),
    .C(_804_),
    .Y(_34_)
);

NAND2X1 _7118_ (
    .A(\genblk1[0].u_ce.Acalc [9]),
    .B(_158__bF$buf4),
    .Y(_820_)
);

OAI21X1 _7119_ (
    .A(_811_),
    .B(_813_),
    .C(_818_),
    .Y(_821_)
);

INVX1 _7120_ (
    .A(\genblk1[0].u_ce.Ain12b [9]),
    .Y(_822_)
);

NAND2X1 _7121_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf4 ),
    .B(_822_),
    .Y(_823_)
);

NOR2X1 _7122_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf3 ),
    .B(_822_),
    .Y(_824_)
);

INVX1 _7123_ (
    .A(_824_),
    .Y(_825_)
);

NAND2X1 _7124_ (
    .A(_823_),
    .B(_825_),
    .Y(_826_)
);

INVX1 _7125_ (
    .A(_826_),
    .Y(_827_)
);

NOR2X1 _7126_ (
    .A(_827_),
    .B(_821_),
    .Y(_828_)
);

NAND2X1 _7127_ (
    .A(_827_),
    .B(_821_),
    .Y(_829_)
);

NAND2X1 _7128_ (
    .A(\genblk1[0].u_ce.Vld_bF$buf3 ),
    .B(_829_),
    .Y(_830_)
);

OAI21X1 _7129_ (
    .A(_828_),
    .B(_830_),
    .C(_820_),
    .Y(_35_)
);

AOI21X1 _7130_ (
    .A(_821_),
    .B(_823_),
    .C(_824_),
    .Y(_831_)
);

INVX1 _7131_ (
    .A(\genblk1[0].u_ce.Ain12b [10]),
    .Y(_832_)
);

NAND2X1 _7132_ (
    .A(\genblk1[0].u_ce.Ain12b_11_bF$buf2 ),
    .B(_832_),
    .Y(_833_)
);

NAND2X1 _7133_ (
    .A(\genblk1[0].u_ce.Ain12b [10]),
    .B(_253__bF$buf5),
    .Y(_834_)
);

NAND2X1 _7134_ (
    .A(_833_),
    .B(_834_),
    .Y(_835_)
);

AND2X2 _7135_ (
    .A(_831_),
    .B(_835_),
    .Y(_836_)
);

OAI21X1 _7136_ (
    .A(_835_),
    .B(_831_),
    .C(\genblk1[0].u_ce.Vld_bF$buf2 ),
    .Y(_837_)
);

OAI22X1 _7137_ (
    .A(_93_),
    .B(\genblk1[0].u_ce.Vld_bF$buf1 ),
    .C(_837_),
    .D(_836_),
    .Y(_36_)
);

NAND2X1 _7138_ (
    .A(\genblk1[0].u_ce.Acalc [11]),
    .B(_158__bF$buf3),
    .Y(_838_)
);

OAI21X1 _7139_ (
    .A(_835_),
    .B(_831_),
    .C(_834_),
    .Y(_839_)
);

OAI21X1 _7140_ (
    .A(_158__bF$buf2),
    .B(_839_),
    .C(_838_),
    .Y(_37_)
);

INVX1 _7141_ (
    .A(_92_),
    .Y(_840_)
);

NAND3X1 _7142_ (
    .A(_145_),
    .B(\genblk1[0].u_ce.LoadCtl [5]),
    .C(_103_),
    .Y(_841_)
);

NOR2X1 _7143_ (
    .A(_840_),
    .B(_841_),
    .Y(_842_)
);

NAND2X1 _7144_ (
    .A(1'h0),
    .B(_842_),
    .Y(_843_)
);

OAI21X1 _7145_ (
    .A(_287_),
    .B(_842_),
    .C(_843_),
    .Y(_38_)
);

NAND2X1 _7146_ (
    .A(1'h0),
    .B(_842_),
    .Y(_844_)
);

OAI21X1 _7147_ (
    .A(_312_),
    .B(_842_),
    .C(_844_),
    .Y(_39_)
);

INVX1 _7148_ (
    .A(1'h0),
    .Y(_845_)
);

NAND3X1 _7149_ (
    .A(\genblk1[0].u_ce.LoadCtl [4]),
    .B(_92_),
    .C(_103_),
    .Y(_846_)
);

NAND2X1 _7150_ (
    .A(\genblk1[0].u_ce.Xin12b [8]),
    .B(_846_),
    .Y(_847_)
);

OAI21X1 _7151_ (
    .A(_845_),
    .B(_846_),
    .C(_847_),
    .Y(_40_)
);

INVX1 _7152_ (
    .A(1'h0),
    .Y(_848_)
);

NAND2X1 _7153_ (
    .A(\genblk1[0].u_ce.Xin12b [9]),
    .B(_846_),
    .Y(_849_)
);

OAI21X1 _7154_ (
    .A(_848_),
    .B(_846_),
    .C(_849_),
    .Y(_41_)
);

NAND2X1 _7155_ (
    .A(_103_),
    .B(_99_),
    .Y(_850_)
);

OAI21X1 _7156_ (
    .A(_104_),
    .B(_112_),
    .C(\genblk1[0].u_ce.Xin12b [6]),
    .Y(_851_)
);

OAI21X1 _7157_ (
    .A(_845_),
    .B(_850_),
    .C(_851_),
    .Y(_42_)
);

OAI21X1 _7158_ (
    .A(_104_),
    .B(_112_),
    .C(\genblk1[0].u_ce.Xin12b [7]),
    .Y(_852_)
);

OAI21X1 _7159_ (
    .A(_848_),
    .B(_850_),
    .C(_852_),
    .Y(_43_)
);

NOR2X1 _7160_ (
    .A(_96_),
    .B(_104_),
    .Y(_853_)
);

NAND2X1 _7161_ (
    .A(1'h0),
    .B(_853_),
    .Y(_854_)
);

OAI21X1 _7162_ (
    .A(_197_),
    .B(_853_),
    .C(_854_),
    .Y(_44_)
);

NAND2X1 _7163_ (
    .A(1'h0),
    .B(_853_),
    .Y(_855_)
);

OAI21X1 _7164_ (
    .A(_205_),
    .B(_853_),
    .C(_855_),
    .Y(_45_)
);

OAI21X1 _7165_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_105_),
    .C(\genblk1[0].u_ce.Xin1 [0]),
    .Y(_856_)
);

OAI21X1 _7166_ (
    .A(_845_),
    .B(_134_),
    .C(_856_),
    .Y(_46_)
);

OAI21X1 _7167_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_105_),
    .C(\genblk1[0].u_ce.Xin1 [1]),
    .Y(_857_)
);

OAI21X1 _7168_ (
    .A(_848_),
    .B(_134_),
    .C(_857_),
    .Y(_47_)
);

NAND2X1 _7169_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 ),
    .B(1'h0),
    .Y(_858_)
);

OAI21X1 _7170_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_220_),
    .C(_858_),
    .Y(_48_)
);

NAND2X1 _7171_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .B(1'h0),
    .Y(_859_)
);

OAI21X1 _7172_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_200_),
    .C(_859_),
    .Y(_49_)
);

NAND2X1 _7173_ (
    .A(1'h0),
    .B(_842_),
    .Y(_860_)
);

OAI21X1 _7174_ (
    .A(_420_),
    .B(_842_),
    .C(_860_),
    .Y(_50_)
);

NAND2X1 _7175_ (
    .A(1'h0),
    .B(_842_),
    .Y(_861_)
);

OAI21X1 _7176_ (
    .A(_444_),
    .B(_842_),
    .C(_861_),
    .Y(_51_)
);

INVX1 _7177_ (
    .A(1'h0),
    .Y(_862_)
);

NAND2X1 _7178_ (
    .A(\genblk1[0].u_ce.Yin12b [8]),
    .B(_846_),
    .Y(_863_)
);

OAI21X1 _7179_ (
    .A(_862_),
    .B(_846_),
    .C(_863_),
    .Y(_52_)
);

INVX1 _7180_ (
    .A(1'h0),
    .Y(_864_)
);

NAND2X1 _7181_ (
    .A(\genblk1[0].u_ce.Yin12b [9]),
    .B(_846_),
    .Y(_865_)
);

OAI21X1 _7182_ (
    .A(_864_),
    .B(_846_),
    .C(_865_),
    .Y(_53_)
);

OAI21X1 _7183_ (
    .A(_104_),
    .B(_112_),
    .C(\genblk1[0].u_ce.Yin12b [6]),
    .Y(_72_)
);

OAI21X1 _7184_ (
    .A(_862_),
    .B(_850_),
    .C(_72_),
    .Y(_54_)
);

OAI21X1 _7185_ (
    .A(_104_),
    .B(_112_),
    .C(\genblk1[0].u_ce.Yin12b [7]),
    .Y(_73_)
);

OAI21X1 _7186_ (
    .A(_864_),
    .B(_850_),
    .C(_73_),
    .Y(_55_)
);

NAND2X1 _7187_ (
    .A(1'h0),
    .B(_853_),
    .Y(_74_)
);

OAI21X1 _7188_ (
    .A(_285_),
    .B(_853_),
    .C(_74_),
    .Y(_56_)
);

NAND2X1 _7189_ (
    .A(1'h0),
    .B(_853_),
    .Y(_75_)
);

OAI21X1 _7190_ (
    .A(_310_),
    .B(_853_),
    .C(_75_),
    .Y(_57_)
);

OAI21X1 _7191_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_105_),
    .C(\genblk1[0].u_ce.Yin1 [0]),
    .Y(_76_)
);

OAI21X1 _7192_ (
    .A(_862_),
    .B(_134_),
    .C(_76_),
    .Y(_58_)
);

OAI21X1 _7193_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_105_),
    .C(\genblk1[0].u_ce.Yin1 [1]),
    .Y(_77_)
);

OAI21X1 _7194_ (
    .A(_864_),
    .B(_134_),
    .C(_77_),
    .Y(_59_)
);

NAND2X1 _7195_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(1'h0),
    .Y(_78_)
);

OAI21X1 _7196_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_457_),
    .C(_78_),
    .Y(_60_)
);

NAND2X1 _7197_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf2 ),
    .B(1'h0),
    .Y(_79_)
);

OAI21X1 _7198_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_242_),
    .C(_79_),
    .Y(_61_)
);

NAND2X1 _7199_ (
    .A(\a[0] [0]),
    .B(_842_),
    .Y(_80_)
);

OAI21X1 _7200_ (
    .A(_832_),
    .B(_842_),
    .C(_80_),
    .Y(_62_)
);

NAND2X1 _7201_ (
    .A(\a[0] [1]),
    .B(_842_),
    .Y(_81_)
);

OAI21X1 _7202_ (
    .A(_253__bF$buf4),
    .B(_842_),
    .C(_81_),
    .Y(_63_)
);

INVX1 _7203_ (
    .A(\a[0] [0]),
    .Y(_82_)
);

NAND2X1 _7204_ (
    .A(\genblk1[0].u_ce.Ain12b [8]),
    .B(_846_),
    .Y(_83_)
);

OAI21X1 _7205_ (
    .A(_82_),
    .B(_846_),
    .C(_83_),
    .Y(_64_)
);

INVX1 _7206_ (
    .A(\a[0] [1]),
    .Y(_84_)
);

NAND2X1 _7207_ (
    .A(\genblk1[0].u_ce.Ain12b [9]),
    .B(_846_),
    .Y(_85_)
);

OAI21X1 _7208_ (
    .A(_84_),
    .B(_846_),
    .C(_85_),
    .Y(_65_)
);

OAI21X1 _7209_ (
    .A(_104_),
    .B(_112_),
    .C(\genblk1[0].u_ce.Ain12b [6]),
    .Y(_86_)
);

OAI21X1 _7210_ (
    .A(_82_),
    .B(_850_),
    .C(_86_),
    .Y(_66_)
);

OAI21X1 _7211_ (
    .A(_104_),
    .B(_112_),
    .C(\genblk1[0].u_ce.Ain12b [7]),
    .Y(_87_)
);

OAI21X1 _7212_ (
    .A(_84_),
    .B(_850_),
    .C(_87_),
    .Y(_67_)
);

NAND2X1 _7213_ (
    .A(\a[0] [0]),
    .B(_853_),
    .Y(_88_)
);

OAI21X1 _7214_ (
    .A(_756_),
    .B(_853_),
    .C(_88_),
    .Y(_68_)
);

NAND2X1 _7215_ (
    .A(\a[0] [1]),
    .B(_853_),
    .Y(_89_)
);

OAI21X1 _7216_ (
    .A(_770_),
    .B(_853_),
    .C(_89_),
    .Y(_69_)
);

OAI21X1 _7217_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_105_),
    .C(\genblk1[0].u_ce.Ain1 [0]),
    .Y(_90_)
);

OAI21X1 _7218_ (
    .A(_82_),
    .B(_134_),
    .C(_90_),
    .Y(_70_)
);

OAI21X1 _7219_ (
    .A(\genblk1[0].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_105_),
    .C(\genblk1[0].u_ce.Ain1 [1]),
    .Y(_91_)
);

OAI21X1 _7220_ (
    .A(_84_),
    .B(_134_),
    .C(_91_),
    .Y(_71_)
);

DFFPOSX1 _7221_ (
    .CLK(clk_bF$buf39),
    .D(_0_),
    .Q(\genblk1[0].u_ce.Ain0 [0])
);

DFFPOSX1 _7222_ (
    .CLK(clk_bF$buf38),
    .D(_1_),
    .Q(\genblk1[0].u_ce.Ain0 [1])
);

DFFPOSX1 _7223_ (
    .CLK(clk_bF$buf37),
    .D(_2_),
    .Q(\genblk1[0].u_ce.Ycalc [2])
);

DFFPOSX1 _7224_ (
    .CLK(clk_bF$buf36),
    .D(_3_),
    .Q(\genblk1[0].u_ce.Ycalc [3])
);

DFFPOSX1 _7225_ (
    .CLK(clk_bF$buf35),
    .D(_4_),
    .Q(\genblk1[0].u_ce.Ycalc [4])
);

DFFPOSX1 _7226_ (
    .CLK(clk_bF$buf34),
    .D(_5_),
    .Q(\genblk1[0].u_ce.Ycalc [5])
);

DFFPOSX1 _7227_ (
    .CLK(clk_bF$buf33),
    .D(_6_),
    .Q(\genblk1[0].u_ce.Ycalc [6])
);

DFFPOSX1 _7228_ (
    .CLK(clk_bF$buf32),
    .D(_7_),
    .Q(\genblk1[0].u_ce.Ycalc [7])
);

DFFPOSX1 _7229_ (
    .CLK(clk_bF$buf31),
    .D(_8_),
    .Q(\genblk1[0].u_ce.Ycalc [8])
);

DFFPOSX1 _7230_ (
    .CLK(clk_bF$buf30),
    .D(_9_),
    .Q(\genblk1[0].u_ce.Ycalc [9])
);

DFFPOSX1 _7231_ (
    .CLK(clk_bF$buf29),
    .D(_10_),
    .Q(\genblk1[0].u_ce.Ycalc [10])
);

DFFPOSX1 _7232_ (
    .CLK(clk_bF$buf28),
    .D(_11_),
    .Q(\genblk1[0].u_ce.Ycalc [11])
);

DFFPOSX1 _7233_ (
    .CLK(clk_bF$buf27),
    .D(_12_),
    .Q(\genblk1[0].u_ce.Ycalc [0])
);

DFFPOSX1 _7234_ (
    .CLK(clk_bF$buf26),
    .D(_13_),
    .Q(\genblk1[0].u_ce.Ycalc [1])
);

DFFPOSX1 _7235_ (
    .CLK(clk_bF$buf25),
    .D(_14_),
    .Q(\genblk1[0].u_ce.Xcalc [0])
);

DFFPOSX1 _7236_ (
    .CLK(clk_bF$buf24),
    .D(_15_),
    .Q(\genblk1[0].u_ce.Xcalc [1])
);

DFFPOSX1 _7237_ (
    .CLK(clk_bF$buf23),
    .D(_16_),
    .Q(\genblk1[0].u_ce.Xcalc [2])
);

DFFPOSX1 _7238_ (
    .CLK(clk_bF$buf22),
    .D(_17_),
    .Q(\genblk1[0].u_ce.Xcalc [3])
);

DFFPOSX1 _7239_ (
    .CLK(clk_bF$buf21),
    .D(_18_),
    .Q(\genblk1[0].u_ce.Xcalc [4])
);

DFFPOSX1 _7240_ (
    .CLK(clk_bF$buf20),
    .D(_19_),
    .Q(\genblk1[0].u_ce.Xcalc [5])
);

DFFPOSX1 _7241_ (
    .CLK(clk_bF$buf19),
    .D(_20_),
    .Q(\genblk1[0].u_ce.Xcalc [6])
);

DFFPOSX1 _7242_ (
    .CLK(clk_bF$buf18),
    .D(_21_),
    .Q(\genblk1[0].u_ce.Xcalc [7])
);

DFFPOSX1 _7243_ (
    .CLK(clk_bF$buf17),
    .D(_22_),
    .Q(\genblk1[0].u_ce.Xcalc [8])
);

DFFPOSX1 _7244_ (
    .CLK(clk_bF$buf16),
    .D(_23_),
    .Q(\genblk1[0].u_ce.Xcalc [9])
);

DFFPOSX1 _7245_ (
    .CLK(clk_bF$buf15),
    .D(_24_),
    .Q(\genblk1[0].u_ce.Xcalc [10])
);

DFFPOSX1 _7246_ (
    .CLK(clk_bF$buf14),
    .D(_25_),
    .Q(\genblk1[0].u_ce.Xcalc [11])
);

DFFPOSX1 _7247_ (
    .CLK(clk_bF$buf13),
    .D(_26_),
    .Q(\genblk1[0].u_ce.Acalc [0])
);

DFFPOSX1 _7248_ (
    .CLK(clk_bF$buf12),
    .D(_27_),
    .Q(\genblk1[0].u_ce.Acalc [1])
);

DFFPOSX1 _7249_ (
    .CLK(clk_bF$buf11),
    .D(_28_),
    .Q(\genblk1[0].u_ce.Acalc [2])
);

DFFPOSX1 _7250_ (
    .CLK(clk_bF$buf10),
    .D(_29_),
    .Q(\genblk1[0].u_ce.Acalc [3])
);

DFFPOSX1 _7251_ (
    .CLK(clk_bF$buf9),
    .D(_30_),
    .Q(\genblk1[0].u_ce.Acalc [4])
);

DFFPOSX1 _7252_ (
    .CLK(clk_bF$buf8),
    .D(_31_),
    .Q(\genblk1[0].u_ce.Acalc [5])
);

DFFPOSX1 _7253_ (
    .CLK(clk_bF$buf7),
    .D(_32_),
    .Q(\genblk1[0].u_ce.Acalc [6])
);

DFFPOSX1 _7254_ (
    .CLK(clk_bF$buf6),
    .D(_33_),
    .Q(\genblk1[0].u_ce.Acalc [7])
);

DFFPOSX1 _7255_ (
    .CLK(clk_bF$buf5),
    .D(_34_),
    .Q(\genblk1[0].u_ce.Acalc [8])
);

DFFPOSX1 _7256_ (
    .CLK(clk_bF$buf4),
    .D(_35_),
    .Q(\genblk1[0].u_ce.Acalc [9])
);

DFFPOSX1 _7257_ (
    .CLK(clk_bF$buf3),
    .D(_36_),
    .Q(\genblk1[0].u_ce.Acalc [10])
);

DFFPOSX1 _7258_ (
    .CLK(clk_bF$buf2),
    .D(_37_),
    .Q(\genblk1[0].u_ce.Acalc [11])
);

DFFPOSX1 _7259_ (
    .CLK(clk_bF$buf1),
    .D(_38_),
    .Q(\genblk1[0].u_ce.Xin12b [10])
);

DFFPOSX1 _7260_ (
    .CLK(clk_bF$buf0),
    .D(_39_),
    .Q(\genblk1[0].u_ce.Xin12b [11])
);

DFFPOSX1 _7261_ (
    .CLK(clk_bF$buf75),
    .D(_40_),
    .Q(\genblk1[0].u_ce.Xin12b [8])
);

DFFPOSX1 _7262_ (
    .CLK(clk_bF$buf74),
    .D(_41_),
    .Q(\genblk1[0].u_ce.Xin12b [9])
);

DFFPOSX1 _7263_ (
    .CLK(clk_bF$buf73),
    .D(_42_),
    .Q(\genblk1[0].u_ce.Xin12b [6])
);

DFFPOSX1 _7264_ (
    .CLK(clk_bF$buf72),
    .D(_43_),
    .Q(\genblk1[0].u_ce.Xin12b [7])
);

DFFPOSX1 _7265_ (
    .CLK(clk_bF$buf71),
    .D(_44_),
    .Q(\genblk1[0].u_ce.Xin12b [4])
);

DFFPOSX1 _7266_ (
    .CLK(clk_bF$buf70),
    .D(_45_),
    .Q(\genblk1[0].u_ce.Xin12b [5])
);

DFFPOSX1 _7267_ (
    .CLK(clk_bF$buf69),
    .D(_46_),
    .Q(\genblk1[0].u_ce.Xin1 [0])
);

DFFPOSX1 _7268_ (
    .CLK(clk_bF$buf68),
    .D(_47_),
    .Q(\genblk1[0].u_ce.Xin1 [1])
);

DFFPOSX1 _7269_ (
    .CLK(clk_bF$buf67),
    .D(_48_),
    .Q(\genblk1[0].u_ce.Xin0 [0])
);

DFFPOSX1 _7270_ (
    .CLK(clk_bF$buf66),
    .D(_49_),
    .Q(\genblk1[0].u_ce.Xin0 [1])
);

DFFPOSX1 _7271_ (
    .CLK(clk_bF$buf65),
    .D(_50_),
    .Q(\genblk1[0].u_ce.Yin12b [10])
);

DFFPOSX1 _7272_ (
    .CLK(clk_bF$buf64),
    .D(_51_),
    .Q(\genblk1[0].u_ce.Yin12b [11])
);

DFFPOSX1 _7273_ (
    .CLK(clk_bF$buf63),
    .D(_52_),
    .Q(\genblk1[0].u_ce.Yin12b [8])
);

DFFPOSX1 _7274_ (
    .CLK(clk_bF$buf62),
    .D(_53_),
    .Q(\genblk1[0].u_ce.Yin12b [9])
);

DFFPOSX1 _7275_ (
    .CLK(clk_bF$buf61),
    .D(_54_),
    .Q(\genblk1[0].u_ce.Yin12b [6])
);

DFFPOSX1 _7276_ (
    .CLK(clk_bF$buf60),
    .D(_55_),
    .Q(\genblk1[0].u_ce.Yin12b [7])
);

DFFPOSX1 _7277_ (
    .CLK(clk_bF$buf59),
    .D(_56_),
    .Q(\genblk1[0].u_ce.Yin12b [4])
);

DFFPOSX1 _7278_ (
    .CLK(clk_bF$buf58),
    .D(_57_),
    .Q(\genblk1[0].u_ce.Yin12b [5])
);

DFFPOSX1 _7279_ (
    .CLK(clk_bF$buf57),
    .D(_58_),
    .Q(\genblk1[0].u_ce.Yin1 [0])
);

DFFPOSX1 _7280_ (
    .CLK(clk_bF$buf56),
    .D(_59_),
    .Q(\genblk1[0].u_ce.Yin1 [1])
);

DFFPOSX1 _7281_ (
    .CLK(clk_bF$buf55),
    .D(_60_),
    .Q(\genblk1[0].u_ce.Yin0 [0])
);

DFFPOSX1 _7282_ (
    .CLK(clk_bF$buf54),
    .D(_61_),
    .Q(\genblk1[0].u_ce.Yin0 [1])
);

DFFPOSX1 _7283_ (
    .CLK(clk_bF$buf53),
    .D(_62_),
    .Q(\genblk1[0].u_ce.Ain12b [10])
);

DFFPOSX1 _7284_ (
    .CLK(clk_bF$buf52),
    .D(_63_),
    .Q(\genblk1[0].u_ce.Ain12b [11])
);

DFFPOSX1 _7285_ (
    .CLK(clk_bF$buf51),
    .D(_64_),
    .Q(\genblk1[0].u_ce.Ain12b [8])
);

DFFPOSX1 _7286_ (
    .CLK(clk_bF$buf50),
    .D(_65_),
    .Q(\genblk1[0].u_ce.Ain12b [9])
);

DFFPOSX1 _7287_ (
    .CLK(clk_bF$buf49),
    .D(_66_),
    .Q(\genblk1[0].u_ce.Ain12b [6])
);

DFFPOSX1 _7288_ (
    .CLK(clk_bF$buf48),
    .D(_67_),
    .Q(\genblk1[0].u_ce.Ain12b [7])
);

DFFPOSX1 _7289_ (
    .CLK(clk_bF$buf47),
    .D(_68_),
    .Q(\genblk1[0].u_ce.Ain12b [4])
);

DFFPOSX1 _7290_ (
    .CLK(clk_bF$buf46),
    .D(_69_),
    .Q(\genblk1[0].u_ce.Ain12b [5])
);

DFFPOSX1 _7291_ (
    .CLK(clk_bF$buf45),
    .D(_70_),
    .Q(\genblk1[0].u_ce.Ain1 [0])
);

DFFPOSX1 _7292_ (
    .CLK(clk_bF$buf44),
    .D(_71_),
    .Q(\genblk1[0].u_ce.Ain1 [1])
);

DFFPOSX1 _7293_ (
    .CLK(clk_bF$buf43),
    .D(\genblk1[0].u_ce.ISin ),
    .Q(\genblk1[0].u_ce.ISpipe [0])
);

DFFPOSX1 _7294_ (
    .CLK(clk_bF$buf42),
    .D(\genblk1[0].u_ce.ISpipe [0]),
    .Q(\genblk1[0].u_ce.ISpipe [1])
);

DFFPOSX1 _7295_ (
    .CLK(clk_bF$buf41),
    .D(\genblk1[0].u_ce.ISpipe [1]),
    .Q(\genblk1[0].u_ce.ISpipe [2])
);

DFFPOSX1 _7296_ (
    .CLK(clk_bF$buf40),
    .D(\genblk1[0].u_ce.ISpipe [2]),
    .Q(\genblk1[0].u_ce.ISpipe [3])
);

DFFPOSX1 _7297_ (
    .CLK(clk_bF$buf39),
    .D(\genblk1[0].u_ce.ISpipe [3]),
    .Q(\genblk1[0].u_ce.ISpipe [4])
);

DFFPOSX1 _7298_ (
    .CLK(clk_bF$buf38),
    .D(\genblk1[0].u_ce.ISpipe [4]),
    .Q(\genblk1[0].u_ce.ISpipe [5])
);

DFFPOSX1 _7299_ (
    .CLK(clk_bF$buf37),
    .D(\genblk1[0].u_ce.ISpipe [5]),
    .Q(\genblk1[0].u_ce.ISout )
);

DFFPOSX1 _7300_ (
    .CLK(clk_bF$buf36),
    .D(\genblk1[0].u_ce.Rdy ),
    .Q(\genblk1[0].u_ce.LoadCtl [0])
);

DFFPOSX1 _7301_ (
    .CLK(clk_bF$buf35),
    .D(\genblk1[0].u_ce.LoadCtl_0_bF$buf3 ),
    .Q(\genblk1[0].u_ce.LoadCtl [1])
);

DFFPOSX1 _7302_ (
    .CLK(clk_bF$buf34),
    .D(\genblk1[0].u_ce.LoadCtl [1]),
    .Q(\genblk1[0].u_ce.LoadCtl [2])
);

DFFPOSX1 _7303_ (
    .CLK(clk_bF$buf33),
    .D(\genblk1[0].u_ce.LoadCtl [2]),
    .Q(\genblk1[0].u_ce.LoadCtl [3])
);

DFFPOSX1 _7304_ (
    .CLK(clk_bF$buf32),
    .D(\genblk1[0].u_ce.LoadCtl [3]),
    .Q(\genblk1[0].u_ce.LoadCtl [4])
);

DFFPOSX1 _7305_ (
    .CLK(clk_bF$buf31),
    .D(\genblk1[0].u_ce.LoadCtl [4]),
    .Q(\genblk1[0].u_ce.LoadCtl [5])
);

DFFPOSX1 _7306_ (
    .CLK(clk_bF$buf30),
    .D(\genblk1[0].u_ce.LoadCtl [5]),
    .Q(\genblk1[0].u_ce.Vld )
);

NOR2X1 _7307_ (
    .A(\genblk1[1].u_ce.LoadCtl [3]),
    .B(\genblk1[1].u_ce.LoadCtl [2]),
    .Y(_958_)
);

INVX1 _7308_ (
    .A(\genblk1[1].u_ce.Acalc [10]),
    .Y(_959_)
);

NAND2X1 _7309_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(\genblk1[1].u_ce.Acalc [8]),
    .Y(_960_)
);

OAI21X1 _7310_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(_959_),
    .C(_960_),
    .Y(_961_)
);

INVX2 _7311_ (
    .A(\genblk1[1].u_ce.LoadCtl [2]),
    .Y(_962_)
);

INVX1 _7312_ (
    .A(\genblk1[1].u_ce.Acalc [4]),
    .Y(_963_)
);

INVX1 _7313_ (
    .A(\genblk1[1].u_ce.LoadCtl [3]),
    .Y(_964_)
);

NOR2X1 _7314_ (
    .A(\genblk1[1].u_ce.LoadCtl [2]),
    .B(_964_),
    .Y(_965_)
);

NAND2X1 _7315_ (
    .A(\genblk1[1].u_ce.Acalc [6]),
    .B(_965_),
    .Y(_966_)
);

OAI21X1 _7316_ (
    .A(_962_),
    .B(_963_),
    .C(_966_),
    .Y(_967_)
);

AOI21X1 _7317_ (
    .A(_958_),
    .B(_961_),
    .C(_967_),
    .Y(_968_)
);

NOR2X1 _7318_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[1].u_ce.LoadCtl [1]),
    .Y(_969_)
);

INVX4 _7319_ (
    .A(_969_),
    .Y(_970_)
);

INVX2 _7320_ (
    .A(\genblk1[1].u_ce.LoadCtl [1]),
    .Y(_971_)
);

NOR2X1 _7321_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_971_),
    .Y(_972_)
);

AOI22X1 _7322_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[1].u_ce.Acalc [0]),
    .C(_972_),
    .D(\genblk1[1].u_ce.Acalc [2]),
    .Y(_973_)
);

OAI21X1 _7323_ (
    .A(_970_),
    .B(_968_),
    .C(_973_),
    .Y(\a[2] [0])
);

INVX1 _7324_ (
    .A(\genblk1[1].u_ce.Acalc [11]),
    .Y(_974_)
);

NAND2X1 _7325_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(\genblk1[1].u_ce.Acalc [9]),
    .Y(_975_)
);

OAI21X1 _7326_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(_974_),
    .C(_975_),
    .Y(_976_)
);

INVX1 _7327_ (
    .A(\genblk1[1].u_ce.Acalc [7]),
    .Y(_977_)
);

INVX4 _7328_ (
    .A(_965_),
    .Y(_978_)
);

NAND2X1 _7329_ (
    .A(\genblk1[1].u_ce.LoadCtl [2]),
    .B(\genblk1[1].u_ce.Acalc [5]),
    .Y(_979_)
);

OAI21X1 _7330_ (
    .A(_977_),
    .B(_978_),
    .C(_979_),
    .Y(_980_)
);

AOI21X1 _7331_ (
    .A(_958_),
    .B(_976_),
    .C(_980_),
    .Y(_981_)
);

AOI22X1 _7332_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[1].u_ce.Acalc [1]),
    .C(_972_),
    .D(\genblk1[1].u_ce.Acalc [3]),
    .Y(_982_)
);

OAI21X1 _7333_ (
    .A(_970_),
    .B(_981_),
    .C(_982_),
    .Y(\a[2] [1])
);

INVX1 _7334_ (
    .A(\genblk1[1].u_ce.Ycalc [10]),
    .Y(_983_)
);

NAND2X1 _7335_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(\genblk1[1].u_ce.Ycalc [8]),
    .Y(_984_)
);

OAI21X1 _7336_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(_983_),
    .C(_984_),
    .Y(_985_)
);

INVX1 _7337_ (
    .A(\genblk1[1].u_ce.Ycalc [6]),
    .Y(_986_)
);

INVX1 _7338_ (
    .A(\genblk1[1].u_ce.Ycalc [4]),
    .Y(_987_)
);

OAI22X1 _7339_ (
    .A(_962_),
    .B(_987_),
    .C(_986_),
    .D(_978_),
    .Y(_988_)
);

AOI21X1 _7340_ (
    .A(_958_),
    .B(_985_),
    .C(_988_),
    .Y(_989_)
);

AOI22X1 _7341_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[1].u_ce.Ycalc [0]),
    .C(_972_),
    .D(\genblk1[1].u_ce.Ycalc [2]),
    .Y(_990_)
);

OAI21X1 _7342_ (
    .A(_970_),
    .B(_989_),
    .C(_990_),
    .Y(\genblk1[1].u_ce.Y_ [0])
);

INVX1 _7343_ (
    .A(\genblk1[1].u_ce.Ycalc [11]),
    .Y(_991_)
);

NAND2X1 _7344_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(\genblk1[1].u_ce.Ycalc [9]),
    .Y(_992_)
);

OAI21X1 _7345_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(_991_),
    .C(_992_),
    .Y(_993_)
);

INVX1 _7346_ (
    .A(\genblk1[1].u_ce.Ycalc [7]),
    .Y(_994_)
);

INVX1 _7347_ (
    .A(\genblk1[1].u_ce.Ycalc [5]),
    .Y(_995_)
);

OAI22X1 _7348_ (
    .A(_962_),
    .B(_995_),
    .C(_994_),
    .D(_978_),
    .Y(_996_)
);

AOI21X1 _7349_ (
    .A(_958_),
    .B(_993_),
    .C(_996_),
    .Y(_997_)
);

AOI22X1 _7350_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[1].u_ce.Ycalc [1]),
    .C(_972_),
    .D(\genblk1[1].u_ce.Ycalc [3]),
    .Y(_998_)
);

OAI21X1 _7351_ (
    .A(_970_),
    .B(_997_),
    .C(_998_),
    .Y(\genblk1[1].u_ce.Y_ [1])
);

INVX1 _7352_ (
    .A(\genblk1[1].u_ce.Xcalc [2]),
    .Y(_999_)
);

INVX2 _7353_ (
    .A(_972_),
    .Y(_1000_)
);

INVX1 _7354_ (
    .A(\genblk1[1].u_ce.Xcalc [4]),
    .Y(_1001_)
);

INVX1 _7355_ (
    .A(\genblk1[1].u_ce.Xcalc [6]),
    .Y(_1002_)
);

NOR2X1 _7356_ (
    .A(_964_),
    .B(_1002_),
    .Y(_1003_)
);

INVX1 _7357_ (
    .A(\genblk1[1].u_ce.Xcalc [8]),
    .Y(_1004_)
);

NAND2X1 _7358_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(_1004_),
    .Y(_1005_)
);

OAI21X1 _7359_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(\genblk1[1].u_ce.Xcalc [10]),
    .C(_1005_),
    .Y(_1006_)
);

NOR2X1 _7360_ (
    .A(\genblk1[1].u_ce.LoadCtl [3]),
    .B(_1006_),
    .Y(_1007_)
);

OAI21X1 _7361_ (
    .A(_1003_),
    .B(_1007_),
    .C(_962_),
    .Y(_1008_)
);

OAI21X1 _7362_ (
    .A(_962_),
    .B(_1001_),
    .C(_1008_),
    .Y(_1009_)
);

AOI22X1 _7363_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[1].u_ce.Xcalc [0]),
    .C(_1009_),
    .D(_969_),
    .Y(_1010_)
);

OAI21X1 _7364_ (
    .A(_999_),
    .B(_1000_),
    .C(_1010_),
    .Y(\genblk1[1].u_ce.X_ [0])
);

INVX1 _7365_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .Y(_1011_)
);

INVX1 _7366_ (
    .A(\genblk1[1].u_ce.Xcalc [9]),
    .Y(_1012_)
);

NAND2X1 _7367_ (
    .A(\genblk1[1].u_ce.Xcalc [11]),
    .B(_1011_),
    .Y(_1013_)
);

OAI21X1 _7368_ (
    .A(_1011_),
    .B(_1012_),
    .C(_1013_),
    .Y(_1014_)
);

INVX1 _7369_ (
    .A(\genblk1[1].u_ce.Xcalc [7]),
    .Y(_1015_)
);

INVX1 _7370_ (
    .A(\genblk1[1].u_ce.Xcalc [5]),
    .Y(_1016_)
);

OAI22X1 _7371_ (
    .A(_962_),
    .B(_1016_),
    .C(_1015_),
    .D(_978_),
    .Y(_1017_)
);

AOI21X1 _7372_ (
    .A(_958_),
    .B(_1014_),
    .C(_1017_),
    .Y(_1018_)
);

AOI22X1 _7373_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[1].u_ce.Xcalc [1]),
    .C(_972_),
    .D(\genblk1[1].u_ce.Xcalc [3]),
    .Y(_1019_)
);

OAI21X1 _7374_ (
    .A(_970_),
    .B(_1018_),
    .C(_1019_),
    .Y(\genblk1[1].u_ce.X_ [1])
);

INVX1 _7375_ (
    .A(\genblk1[1].u_ce.Ain0 [0]),
    .Y(_1020_)
);

NAND2X1 _7376_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\a[1] [0]),
    .Y(_1021_)
);

OAI21X1 _7377_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_1020_),
    .C(_1021_),
    .Y(_866_)
);

INVX1 _7378_ (
    .A(\genblk1[1].u_ce.Ain0 [1]),
    .Y(_1022_)
);

NAND2X1 _7379_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\a[1] [1]),
    .Y(_1023_)
);

OAI21X1 _7380_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_1022_),
    .C(_1023_),
    .Y(_867_)
);

INVX8 _7381_ (
    .A(\genblk1[1].u_ce.Vld_bF$buf4 ),
    .Y(_1024_)
);

NAND2X1 _7382_ (
    .A(\genblk1[1].u_ce.Ycalc [2]),
    .B(_1024__bF$buf4),
    .Y(_1025_)
);

INVX2 _7383_ (
    .A(1'h1),
    .Y(_1026_)
);

NOR2X1 _7384_ (
    .A(1'h0),
    .B(1'h0),
    .Y(_1027_)
);

NAND2X1 _7385_ (
    .A(_1026_),
    .B(_1027_),
    .Y(_1028_)
);

INVX2 _7386_ (
    .A(_1028_),
    .Y(_1029_)
);

INVX8 _7387_ (
    .A(1'h0),
    .Y(_1030_)
);

MUX2X1 _7388_ (
    .A(\genblk1[1].u_ce.Xin12b [4]),
    .B(\genblk1[1].u_ce.Xin1 [1]),
    .S(1'h1),
    .Y(_1031_)
);

MUX2X1 _7389_ (
    .A(\genblk1[1].u_ce.Xin1 [0]),
    .B(\genblk1[1].u_ce.Xin0 [1]),
    .S(1'h1),
    .Y(_1032_)
);

MUX2X1 _7390_ (
    .A(_1032_),
    .B(_1031_),
    .S(_1030__bF$buf4),
    .Y(_1033_)
);

MUX2X1 _7391_ (
    .A(\genblk1[1].u_ce.Xin12b [8]),
    .B(\genblk1[1].u_ce.Xin12b [7]),
    .S(1'h1),
    .Y(_1034_)
);

MUX2X1 _7392_ (
    .A(\genblk1[1].u_ce.Xin12b [6]),
    .B(\genblk1[1].u_ce.Xin12b [5]),
    .S(1'h1),
    .Y(_1035_)
);

MUX2X1 _7393_ (
    .A(_1035_),
    .B(_1034_),
    .S(_1030__bF$buf3),
    .Y(_1036_)
);

MUX2X1 _7394_ (
    .A(_1036_),
    .B(_1033_),
    .S(1'h0),
    .Y(_1037_)
);

INVX1 _7395_ (
    .A(_1037_),
    .Y(_1038_)
);

MUX2X1 _7396_ (
    .A(\genblk1[1].u_ce.Xin1 [1]),
    .B(\genblk1[1].u_ce.Xin1 [0]),
    .S(1'h1),
    .Y(_1039_)
);

MUX2X1 _7397_ (
    .A(\genblk1[1].u_ce.Xin0 [1]),
    .B(\genblk1[1].u_ce.Xin0 [0]),
    .S(1'h1),
    .Y(_1040_)
);

MUX2X1 _7398_ (
    .A(_1040_),
    .B(_1039_),
    .S(_1030__bF$buf2),
    .Y(_1041_)
);

MUX2X1 _7399_ (
    .A(\genblk1[1].u_ce.Xin12b [7]),
    .B(\genblk1[1].u_ce.Xin12b [6]),
    .S(1'h1),
    .Y(_1042_)
);

MUX2X1 _7400_ (
    .A(\genblk1[1].u_ce.Xin12b [5]),
    .B(\genblk1[1].u_ce.Xin12b [4]),
    .S(1'h1),
    .Y(_1043_)
);

MUX2X1 _7401_ (
    .A(_1043_),
    .B(_1042_),
    .S(_1030__bF$buf1),
    .Y(_1044_)
);

MUX2X1 _7402_ (
    .A(_1044_),
    .B(_1041_),
    .S(1'h0),
    .Y(_1045_)
);

OAI21X1 _7403_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf4 ),
    .B(_1045_),
    .C(_1038_),
    .Y(_1046_)
);

NOR2X1 _7404_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1045_),
    .Y(_1047_)
);

NAND2X1 _7405_ (
    .A(_1037_),
    .B(_1047_),
    .Y(_1048_)
);

NAND3X1 _7406_ (
    .A(\genblk1[1].u_ce.Yin0 [1]),
    .B(_1046_),
    .C(_1048_),
    .Y(_1049_)
);

NOR2X1 _7407_ (
    .A(\genblk1[1].u_ce.Yin0 [0]),
    .B(_1045_),
    .Y(_1050_)
);

AOI21X1 _7408_ (
    .A(_1048_),
    .B(_1046_),
    .C(\genblk1[1].u_ce.Yin0 [1]),
    .Y(_1051_)
);

OAI21X1 _7409_ (
    .A(_1050_),
    .B(_1051_),
    .C(_1049_),
    .Y(_1052_)
);

INVX1 _7410_ (
    .A(\genblk1[1].u_ce.Yin1 [0]),
    .Y(_1053_)
);

MUX2X1 _7411_ (
    .A(\genblk1[1].u_ce.Xin12b [9]),
    .B(\genblk1[1].u_ce.Xin12b [8]),
    .S(1'h1),
    .Y(_1054_)
);

MUX2X1 _7412_ (
    .A(_1054_),
    .B(_1042_),
    .S(1'h0),
    .Y(_1055_)
);

AND2X2 _7413_ (
    .A(_1055_),
    .B(1'h0),
    .Y(_1056_)
);

INVX4 _7414_ (
    .A(1'h0),
    .Y(_1057_)
);

NAND2X1 _7415_ (
    .A(_1057__bF$buf3),
    .B(_1030__bF$buf0),
    .Y(_1058_)
);

NAND2X1 _7416_ (
    .A(1'h0),
    .B(_1057__bF$buf2),
    .Y(_1059_)
);

OAI22X1 _7417_ (
    .A(_1058_),
    .B(_1039_),
    .C(_1043_),
    .D(_1059_),
    .Y(_1060_)
);

INVX1 _7418_ (
    .A(\genblk1[1].u_ce.Xin1 [1]),
    .Y(_1061_)
);

NAND2X1 _7419_ (
    .A(_1026_),
    .B(_1061_),
    .Y(_1062_)
);

INVX1 _7420_ (
    .A(\genblk1[1].u_ce.Xin12b [4]),
    .Y(_1063_)
);

NAND2X1 _7421_ (
    .A(1'h1),
    .B(_1063_),
    .Y(_1064_)
);

NAND3X1 _7422_ (
    .A(1'h0),
    .B(_1064_),
    .C(_1062_),
    .Y(_1065_)
);

INVX1 _7423_ (
    .A(\genblk1[1].u_ce.Xin0 [1]),
    .Y(_1066_)
);

NAND2X1 _7424_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Xin1 [0]),
    .Y(_1067_)
);

OAI21X1 _7425_ (
    .A(1'h1),
    .B(_1066_),
    .C(_1067_),
    .Y(_1068_)
);

NAND2X1 _7426_ (
    .A(_1030__bF$buf4),
    .B(_1068_),
    .Y(_1069_)
);

NAND3X1 _7427_ (
    .A(_1057__bF$buf1),
    .B(_1065_),
    .C(_1069_),
    .Y(_1070_)
);

INVX1 _7428_ (
    .A(\genblk1[1].u_ce.Xin12b [5]),
    .Y(_1071_)
);

NAND2X1 _7429_ (
    .A(_1026_),
    .B(_1071_),
    .Y(_1072_)
);

INVX1 _7430_ (
    .A(\genblk1[1].u_ce.Xin12b [6]),
    .Y(_1073_)
);

NAND2X1 _7431_ (
    .A(1'h1),
    .B(_1073_),
    .Y(_1074_)
);

NAND3X1 _7432_ (
    .A(_1030__bF$buf3),
    .B(_1074_),
    .C(_1072_),
    .Y(_1075_)
);

INVX1 _7433_ (
    .A(\genblk1[1].u_ce.Xin12b [7]),
    .Y(_1076_)
);

NAND2X1 _7434_ (
    .A(_1026_),
    .B(_1076_),
    .Y(_1077_)
);

INVX1 _7435_ (
    .A(\genblk1[1].u_ce.Xin12b [8]),
    .Y(_1078_)
);

NAND2X1 _7436_ (
    .A(1'h1),
    .B(_1078_),
    .Y(_1079_)
);

NAND3X1 _7437_ (
    .A(1'h0),
    .B(_1079_),
    .C(_1077_),
    .Y(_1080_)
);

NAND3X1 _7438_ (
    .A(1'h0),
    .B(_1075_),
    .C(_1080_),
    .Y(_1081_)
);

INVX1 _7439_ (
    .A(\genblk1[1].u_ce.Xin1 [0]),
    .Y(_1082_)
);

NAND2X1 _7440_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Xin1 [1]),
    .Y(_1083_)
);

OAI21X1 _7441_ (
    .A(1'h1),
    .B(_1082_),
    .C(_1083_),
    .Y(_1084_)
);

NAND2X1 _7442_ (
    .A(1'h0),
    .B(_1084_),
    .Y(_1085_)
);

INVX1 _7443_ (
    .A(\genblk1[1].u_ce.Xin0 [0]),
    .Y(_1086_)
);

NAND2X1 _7444_ (
    .A(\genblk1[1].u_ce.Xin0 [1]),
    .B(1'h1),
    .Y(_1087_)
);

OAI21X1 _7445_ (
    .A(1'h1),
    .B(_1086_),
    .C(_1087_),
    .Y(_1088_)
);

NAND2X1 _7446_ (
    .A(_1030__bF$buf2),
    .B(_1088_),
    .Y(_1089_)
);

NAND3X1 _7447_ (
    .A(_1057__bF$buf0),
    .B(_1085_),
    .C(_1089_),
    .Y(_1090_)
);

NAND2X1 _7448_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Xin12b [5]),
    .Y(_1091_)
);

OAI21X1 _7449_ (
    .A(1'h1),
    .B(_1063_),
    .C(_1091_),
    .Y(_1092_)
);

NAND2X1 _7450_ (
    .A(_1030__bF$buf1),
    .B(_1092_),
    .Y(_1093_)
);

NAND2X1 _7451_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Xin12b [7]),
    .Y(_1094_)
);

OAI21X1 _7452_ (
    .A(1'h1),
    .B(_1073_),
    .C(_1094_),
    .Y(_1095_)
);

NAND2X1 _7453_ (
    .A(1'h0),
    .B(_1095_),
    .Y(_1096_)
);

NAND3X1 _7454_ (
    .A(1'h0),
    .B(_1093_),
    .C(_1096_),
    .Y(_1097_)
);

AOI22X1 _7455_ (
    .A(_1070_),
    .B(_1081_),
    .C(_1090_),
    .D(_1097_),
    .Y(_1098_)
);

NOR2X1 _7456_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1098_),
    .Y(_1099_)
);

OAI21X1 _7457_ (
    .A(_1056_),
    .B(_1060_),
    .C(_1099_),
    .Y(_1100_)
);

AOI21X1 _7458_ (
    .A(1'h0),
    .B(_1055_),
    .C(_1060_),
    .Y(_1101_)
);

OAI21X1 _7459_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1098_),
    .C(_1101_),
    .Y(_1102_)
);

NAND3X1 _7460_ (
    .A(_1053_),
    .B(_1102_),
    .C(_1100_),
    .Y(_1103_)
);

NAND2X1 _7461_ (
    .A(_1101_),
    .B(_1099_),
    .Y(_1104_)
);

OAI22X1 _7462_ (
    .A(_1056_),
    .B(_1060_),
    .C(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .D(_1098_),
    .Y(_1105_)
);

NAND3X1 _7463_ (
    .A(\genblk1[1].u_ce.Yin1 [0]),
    .B(_1105_),
    .C(_1104_),
    .Y(_1106_)
);

NAND3X1 _7464_ (
    .A(_1103_),
    .B(_1106_),
    .C(_1052_),
    .Y(_1107_)
);

INVX1 _7465_ (
    .A(\genblk1[1].u_ce.Yin0 [1]),
    .Y(_1108_)
);

NAND2X1 _7466_ (
    .A(_1038_),
    .B(_1047_),
    .Y(_1109_)
);

OAI21X1 _7467_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf4 ),
    .B(_1045_),
    .C(_1037_),
    .Y(_1110_)
);

AOI21X1 _7468_ (
    .A(_1109_),
    .B(_1110_),
    .C(_1108_),
    .Y(_1111_)
);

INVX1 _7469_ (
    .A(_1050_),
    .Y(_1112_)
);

NAND3X1 _7470_ (
    .A(_1108_),
    .B(_1110_),
    .C(_1109_),
    .Y(_1113_)
);

AOI21X1 _7471_ (
    .A(_1112_),
    .B(_1113_),
    .C(_1111_),
    .Y(_1114_)
);

AOI21X1 _7472_ (
    .A(_1104_),
    .B(_1105_),
    .C(\genblk1[1].u_ce.Yin1 [0]),
    .Y(_1115_)
);

AOI21X1 _7473_ (
    .A(_1100_),
    .B(_1102_),
    .C(_1053_),
    .Y(_1116_)
);

OAI21X1 _7474_ (
    .A(_1115_),
    .B(_1116_),
    .C(_1114_),
    .Y(_1117_)
);

AOI21X1 _7475_ (
    .A(_1107_),
    .B(_1117_),
    .C(_1029_),
    .Y(_1118_)
);

INVX8 _7476_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_1119_)
);

NAND3X1 _7477_ (
    .A(_1057__bF$buf3),
    .B(_1026_),
    .C(_1119__bF$buf5),
    .Y(_1120_)
);

OAI21X1 _7478_ (
    .A(1'h0),
    .B(_1120_),
    .C(\genblk1[1].u_ce.Vld_bF$buf3 ),
    .Y(_1121_)
);

OAI21X1 _7479_ (
    .A(_1121_),
    .B(_1118_),
    .C(_1025_),
    .Y(_868_)
);

INVX1 _7480_ (
    .A(\genblk1[1].u_ce.Ycalc [3]),
    .Y(_1122_)
);

INVX1 _7481_ (
    .A(\genblk1[1].u_ce.Xin12b [9]),
    .Y(_1123_)
);

NAND2X1 _7482_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Xin12b [10]),
    .Y(_1124_)
);

OAI21X1 _7483_ (
    .A(1'h1),
    .B(_1123_),
    .C(_1124_),
    .Y(_1125_)
);

NAND2X1 _7484_ (
    .A(1'h0),
    .B(_1125_),
    .Y(_1126_)
);

OAI21X1 _7485_ (
    .A(1'h0),
    .B(_1034_),
    .C(_1126_),
    .Y(_1127_)
);

OAI22X1 _7486_ (
    .A(_1058_),
    .B(_1031_),
    .C(_1035_),
    .D(_1059_),
    .Y(_1128_)
);

AOI21X1 _7487_ (
    .A(_1127_),
    .B(1'h0),
    .C(_1128_),
    .Y(_1129_)
);

NAND3X1 _7488_ (
    .A(_1101_),
    .B(_1037_),
    .C(_1045_),
    .Y(_1130_)
);

INVX1 _7489_ (
    .A(_1130_),
    .Y(_1131_)
);

NOR2X1 _7490_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1131_),
    .Y(_1132_)
);

NAND2X1 _7491_ (
    .A(_1129_),
    .B(_1132_),
    .Y(_1133_)
);

INVX1 _7492_ (
    .A(_1129_),
    .Y(_1134_)
);

OAI21X1 _7493_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1131_),
    .C(_1134_),
    .Y(_1135_)
);

AOI21X1 _7494_ (
    .A(_1133_),
    .B(_1135_),
    .C(\genblk1[1].u_ce.Yin1 [1]),
    .Y(_1136_)
);

AOI21X1 _7495_ (
    .A(_1052_),
    .B(_1103_),
    .C(_1116_),
    .Y(_1137_)
);

NAND3X1 _7496_ (
    .A(\genblk1[1].u_ce.Yin1 [1]),
    .B(_1135_),
    .C(_1133_),
    .Y(_1138_)
);

NAND2X1 _7497_ (
    .A(_1138_),
    .B(_1137_),
    .Y(_1139_)
);

OAI21X1 _7498_ (
    .A(_1115_),
    .B(_1114_),
    .C(_1106_),
    .Y(_1140_)
);

INVX1 _7499_ (
    .A(\genblk1[1].u_ce.Yin1 [1]),
    .Y(_1141_)
);

NAND2X1 _7500_ (
    .A(_1134_),
    .B(_1132_),
    .Y(_1142_)
);

OAI21X1 _7501_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1131_),
    .C(_1129_),
    .Y(_1143_)
);

AOI21X1 _7502_ (
    .A(_1142_),
    .B(_1143_),
    .C(_1141_),
    .Y(_1144_)
);

OAI21X1 _7503_ (
    .A(_1136_),
    .B(_1144_),
    .C(_1140_),
    .Y(_1145_)
);

OAI21X1 _7504_ (
    .A(_1136_),
    .B(_1139_),
    .C(_1145_),
    .Y(_1146_)
);

OAI21X1 _7505_ (
    .A(_1119__bF$buf4),
    .B(_1028_),
    .C(\genblk1[1].u_ce.Vld_bF$buf2 ),
    .Y(_1147_)
);

INVX1 _7506_ (
    .A(_1147_),
    .Y(_1148_)
);

OAI21X1 _7507_ (
    .A(_1029_),
    .B(_1146_),
    .C(_1148_),
    .Y(_1149_)
);

OAI21X1 _7508_ (
    .A(_1122_),
    .B(\genblk1[1].u_ce.Vld_bF$buf1 ),
    .C(_1149_),
    .Y(_869_)
);

INVX1 _7509_ (
    .A(_1121_),
    .Y(_1150_)
);

INVX1 _7510_ (
    .A(\genblk1[1].u_ce.Yin12b [4]),
    .Y(_1151_)
);

NAND3X1 _7511_ (
    .A(_1101_),
    .B(_1129_),
    .C(_1098_),
    .Y(_1152_)
);

INVX1 _7512_ (
    .A(\genblk1[1].u_ce.Xin12b [10]),
    .Y(_1153_)
);

NAND2X1 _7513_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Xin12b [11]),
    .Y(_1154_)
);

OAI21X1 _7514_ (
    .A(1'h1),
    .B(_1153_),
    .C(_1154_),
    .Y(_1155_)
);

NAND2X1 _7515_ (
    .A(_1030__bF$buf0),
    .B(_1054_),
    .Y(_1156_)
);

OAI21X1 _7516_ (
    .A(_1030__bF$buf4),
    .B(_1155_),
    .C(_1156_),
    .Y(_1157_)
);

NAND2X1 _7517_ (
    .A(_1057__bF$buf2),
    .B(_1044_),
    .Y(_1158_)
);

OAI21X1 _7518_ (
    .A(_1057__bF$buf1),
    .B(_1157_),
    .C(_1158_),
    .Y(_1159_)
);

INVX1 _7519_ (
    .A(_1159_),
    .Y(_1160_)
);

NAND3X1 _7520_ (
    .A(_1119__bF$buf3),
    .B(_1160_),
    .C(_1152_),
    .Y(_1161_)
);

INVX1 _7521_ (
    .A(_1161_),
    .Y(_1162_)
);

AOI21X1 _7522_ (
    .A(_1152_),
    .B(_1119__bF$buf2),
    .C(_1160_),
    .Y(_1163_)
);

OAI21X1 _7523_ (
    .A(_1163_),
    .B(_1162_),
    .C(_1151_),
    .Y(_1164_)
);

OAI21X1 _7524_ (
    .A(_1130_),
    .B(_1134_),
    .C(_1119__bF$buf1),
    .Y(_1165_)
);

NAND2X1 _7525_ (
    .A(_1159_),
    .B(_1165_),
    .Y(_1166_)
);

NAND3X1 _7526_ (
    .A(\genblk1[1].u_ce.Yin12b [4]),
    .B(_1161_),
    .C(_1166_),
    .Y(_1167_)
);

NAND2X1 _7527_ (
    .A(_1167_),
    .B(_1164_),
    .Y(_1168_)
);

INVX1 _7528_ (
    .A(_1136_),
    .Y(_1169_)
);

OAI21X1 _7529_ (
    .A(_1144_),
    .B(_1140_),
    .C(_1169_),
    .Y(_1170_)
);

AOI21X1 _7530_ (
    .A(_1170_),
    .B(_1168_),
    .C(_1029_),
    .Y(_1171_)
);

OAI21X1 _7531_ (
    .A(_1168_),
    .B(_1170_),
    .C(_1171_),
    .Y(_1172_)
);

AOI22X1 _7532_ (
    .A(_987_),
    .B(_1024__bF$buf3),
    .C(_1172_),
    .D(_1150_),
    .Y(_870_)
);

INVX1 _7533_ (
    .A(_1167_),
    .Y(_1173_)
);

AOI21X1 _7534_ (
    .A(_1137_),
    .B(_1138_),
    .C(_1136_),
    .Y(_1174_)
);

AOI21X1 _7535_ (
    .A(_1174_),
    .B(_1164_),
    .C(_1173_),
    .Y(_1175_)
);

INVX1 _7536_ (
    .A(\genblk1[1].u_ce.Yin12b [5]),
    .Y(_1176_)
);

NAND3X1 _7537_ (
    .A(_1129_),
    .B(_1160_),
    .C(_1131_),
    .Y(_1177_)
);

INVX1 _7538_ (
    .A(\genblk1[1].u_ce.Xin12b [11]),
    .Y(_1178_)
);

NOR2X1 _7539_ (
    .A(_1030__bF$buf3),
    .B(_1178_),
    .Y(_1179_)
);

AOI21X1 _7540_ (
    .A(_1030__bF$buf2),
    .B(_1125_),
    .C(_1179_),
    .Y(_1180_)
);

NAND2X1 _7541_ (
    .A(_1057__bF$buf0),
    .B(_1036_),
    .Y(_1181_)
);

OAI21X1 _7542_ (
    .A(_1057__bF$buf3),
    .B(_1180_),
    .C(_1181_),
    .Y(_1182_)
);

NAND3X1 _7543_ (
    .A(_1119__bF$buf0),
    .B(_1182_),
    .C(_1177_),
    .Y(_1183_)
);

INVX1 _7544_ (
    .A(_1182_),
    .Y(_1184_)
);

OAI21X1 _7545_ (
    .A(_1159_),
    .B(_1152_),
    .C(_1119__bF$buf5),
    .Y(_1185_)
);

NAND2X1 _7546_ (
    .A(_1184_),
    .B(_1185_),
    .Y(_1186_)
);

NAND3X1 _7547_ (
    .A(_1176_),
    .B(_1186_),
    .C(_1183_),
    .Y(_1187_)
);

NAND3X1 _7548_ (
    .A(_1119__bF$buf4),
    .B(_1184_),
    .C(_1177_),
    .Y(_1188_)
);

NAND2X1 _7549_ (
    .A(_1182_),
    .B(_1185_),
    .Y(_1189_)
);

NAND3X1 _7550_ (
    .A(\genblk1[1].u_ce.Yin12b [5]),
    .B(_1189_),
    .C(_1188_),
    .Y(_1190_)
);

NAND2X1 _7551_ (
    .A(_1187_),
    .B(_1190_),
    .Y(_1191_)
);

INVX1 _7552_ (
    .A(_1191_),
    .Y(_1192_)
);

NOR2X1 _7553_ (
    .A(_1192_),
    .B(_1175_),
    .Y(_1193_)
);

OAI21X1 _7554_ (
    .A(_1168_),
    .B(_1170_),
    .C(_1167_),
    .Y(_1194_)
);

OAI21X1 _7555_ (
    .A(_1191_),
    .B(_1194_),
    .C(_1028_),
    .Y(_1195_)
);

OAI21X1 _7556_ (
    .A(_1195_),
    .B(_1193_),
    .C(_1150_),
    .Y(_1196_)
);

OAI21X1 _7557_ (
    .A(_995_),
    .B(\genblk1[1].u_ce.Vld_bF$buf0 ),
    .C(_1196_),
    .Y(_871_)
);

NOR2X1 _7558_ (
    .A(_1168_),
    .B(_1191_),
    .Y(_1197_)
);

OAI21X1 _7559_ (
    .A(_1167_),
    .B(_1191_),
    .C(_1190_),
    .Y(_1198_)
);

AOI21X1 _7560_ (
    .A(_1197_),
    .B(_1174_),
    .C(_1198_),
    .Y(_1199_)
);

INVX1 _7561_ (
    .A(\genblk1[1].u_ce.Yin12b [6]),
    .Y(_1200_)
);

NOR2X1 _7562_ (
    .A(_1159_),
    .B(_1152_),
    .Y(_1201_)
);

NAND2X1 _7563_ (
    .A(_1184_),
    .B(_1201_),
    .Y(_1202_)
);

AOI21X1 _7564_ (
    .A(_1030__bF$buf1),
    .B(_1155_),
    .C(_1179_),
    .Y(_1203_)
);

NAND2X1 _7565_ (
    .A(_1057__bF$buf2),
    .B(_1055_),
    .Y(_1204_)
);

OAI21X1 _7566_ (
    .A(_1057__bF$buf1),
    .B(_1203_),
    .C(_1204_),
    .Y(_1205_)
);

NAND3X1 _7567_ (
    .A(_1119__bF$buf3),
    .B(_1205_),
    .C(_1202_),
    .Y(_1206_)
);

NOR3X1 _7568_ (
    .A(_1159_),
    .B(_1182_),
    .C(_1152_),
    .Y(_1207_)
);

INVX1 _7569_ (
    .A(_1205_),
    .Y(_1208_)
);

OAI21X1 _7570_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf4 ),
    .B(_1207_),
    .C(_1208_),
    .Y(_1209_)
);

NAND3X1 _7571_ (
    .A(_1200_),
    .B(_1209_),
    .C(_1206_),
    .Y(_1210_)
);

NAND3X1 _7572_ (
    .A(_1119__bF$buf2),
    .B(_1208_),
    .C(_1202_),
    .Y(_1211_)
);

OAI21X1 _7573_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1207_),
    .C(_1205_),
    .Y(_1212_)
);

NAND3X1 _7574_ (
    .A(\genblk1[1].u_ce.Yin12b [6]),
    .B(_1212_),
    .C(_1211_),
    .Y(_1213_)
);

AND2X2 _7575_ (
    .A(_1210_),
    .B(_1213_),
    .Y(_1214_)
);

INVX1 _7576_ (
    .A(_1214_),
    .Y(_1215_)
);

AOI21X1 _7577_ (
    .A(_1199_),
    .B(_1215_),
    .C(_1029_),
    .Y(_1216_)
);

OAI21X1 _7578_ (
    .A(_1199_),
    .B(_1215_),
    .C(_1216_),
    .Y(_1217_)
);

AOI22X1 _7579_ (
    .A(_986_),
    .B(_1024__bF$buf2),
    .C(_1217_),
    .D(_1150_),
    .Y(_872_)
);

AND2X2 _7580_ (
    .A(_1164_),
    .B(_1167_),
    .Y(_1218_)
);

NAND3X1 _7581_ (
    .A(_1187_),
    .B(_1190_),
    .C(_1218_),
    .Y(_1219_)
);

INVX1 _7582_ (
    .A(_1190_),
    .Y(_1220_)
);

AOI21X1 _7583_ (
    .A(_1173_),
    .B(_1187_),
    .C(_1220_),
    .Y(_1221_)
);

OAI21X1 _7584_ (
    .A(_1170_),
    .B(_1219_),
    .C(_1221_),
    .Y(_1222_)
);

INVX1 _7585_ (
    .A(_1213_),
    .Y(_1223_)
);

AOI21X1 _7586_ (
    .A(_1222_),
    .B(_1210_),
    .C(_1223_),
    .Y(_1224_)
);

INVX1 _7587_ (
    .A(\genblk1[1].u_ce.Yin12b [7]),
    .Y(_1225_)
);

NAND2X1 _7588_ (
    .A(_1208_),
    .B(_1207_),
    .Y(_1226_)
);

NOR2X1 _7589_ (
    .A(_1057__bF$buf0),
    .B(_1178_),
    .Y(_1227_)
);

AOI21X1 _7590_ (
    .A(_1127_),
    .B(_1057__bF$buf3),
    .C(_1227_),
    .Y(_1228_)
);

INVX1 _7591_ (
    .A(_1228_),
    .Y(_1229_)
);

NAND3X1 _7592_ (
    .A(_1119__bF$buf1),
    .B(_1229_),
    .C(_1226_),
    .Y(_1230_)
);

AND2X2 _7593_ (
    .A(_1207_),
    .B(_1208_),
    .Y(_1231_)
);

OAI21X1 _7594_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1231_),
    .C(_1228_),
    .Y(_1232_)
);

NAND3X1 _7595_ (
    .A(_1225_),
    .B(_1230_),
    .C(_1232_),
    .Y(_1233_)
);

NAND3X1 _7596_ (
    .A(_1119__bF$buf0),
    .B(_1228_),
    .C(_1226_),
    .Y(_1234_)
);

OAI21X1 _7597_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1231_),
    .C(_1229_),
    .Y(_1235_)
);

NAND3X1 _7598_ (
    .A(\genblk1[1].u_ce.Yin12b [7]),
    .B(_1234_),
    .C(_1235_),
    .Y(_1236_)
);

AND2X2 _7599_ (
    .A(_1233_),
    .B(_1236_),
    .Y(_1237_)
);

NOR2X1 _7600_ (
    .A(_1237_),
    .B(_1224_),
    .Y(_1238_)
);

NAND2X1 _7601_ (
    .A(_1026_),
    .B(_1030__bF$buf0),
    .Y(_1239_)
);

NAND2X1 _7602_ (
    .A(_1237_),
    .B(_1224_),
    .Y(_1240_)
);

OAI21X1 _7603_ (
    .A(1'h0),
    .B(_1239_),
    .C(_1240_),
    .Y(_1241_)
);

OAI21X1 _7604_ (
    .A(_1238_),
    .B(_1241_),
    .C(_1148_),
    .Y(_1242_)
);

OAI21X1 _7605_ (
    .A(_994_),
    .B(\genblk1[1].u_ce.Vld_bF$buf4 ),
    .C(_1242_),
    .Y(_873_)
);

INVX1 _7606_ (
    .A(\genblk1[1].u_ce.Ycalc [8]),
    .Y(_1243_)
);

AOI21X1 _7607_ (
    .A(_1232_),
    .B(_1230_),
    .C(_1225_),
    .Y(_1244_)
);

OAI21X1 _7608_ (
    .A(_1223_),
    .B(_1244_),
    .C(_1233_),
    .Y(_1245_)
);

NAND3X1 _7609_ (
    .A(_1214_),
    .B(_1237_),
    .C(_1222_),
    .Y(_1246_)
);

INVX1 _7610_ (
    .A(\genblk1[1].u_ce.Yin12b [8]),
    .Y(_1247_)
);

NAND3X1 _7611_ (
    .A(_1208_),
    .B(_1228_),
    .C(_1207_),
    .Y(_1248_)
);

INVX1 _7612_ (
    .A(_1227_),
    .Y(_1249_)
);

OAI21X1 _7613_ (
    .A(1'h0),
    .B(_1157_),
    .C(_1249_),
    .Y(_1250_)
);

NAND3X1 _7614_ (
    .A(_1119__bF$buf5),
    .B(_1250_),
    .C(_1248_),
    .Y(_1251_)
);

INVX1 _7615_ (
    .A(_1250_),
    .Y(_1252_)
);

NAND2X1 _7616_ (
    .A(_1119__bF$buf4),
    .B(_1248_),
    .Y(_1253_)
);

NAND2X1 _7617_ (
    .A(_1252_),
    .B(_1253_),
    .Y(_1254_)
);

NAND3X1 _7618_ (
    .A(_1247_),
    .B(_1251_),
    .C(_1254_),
    .Y(_1255_)
);

NAND3X1 _7619_ (
    .A(_1119__bF$buf3),
    .B(_1252_),
    .C(_1248_),
    .Y(_1256_)
);

NAND2X1 _7620_ (
    .A(_1250_),
    .B(_1253_),
    .Y(_1257_)
);

NAND3X1 _7621_ (
    .A(\genblk1[1].u_ce.Yin12b [8]),
    .B(_1256_),
    .C(_1257_),
    .Y(_1258_)
);

AND2X2 _7622_ (
    .A(_1255_),
    .B(_1258_),
    .Y(_1259_)
);

INVX1 _7623_ (
    .A(_1259_),
    .Y(_1260_)
);

AOI21X1 _7624_ (
    .A(_1246_),
    .B(_1245_),
    .C(_1260_),
    .Y(_1261_)
);

NAND3X1 _7625_ (
    .A(_1233_),
    .B(_1236_),
    .C(_1214_),
    .Y(_1262_)
);

OAI21X1 _7626_ (
    .A(_1262_),
    .B(_1199_),
    .C(_1245_),
    .Y(_1263_)
);

OAI21X1 _7627_ (
    .A(_1259_),
    .B(_1263_),
    .C(_1028_),
    .Y(_1264_)
);

OR2X2 _7628_ (
    .A(_1264_),
    .B(_1261_),
    .Y(_1265_)
);

AOI22X1 _7629_ (
    .A(_1243_),
    .B(_1024__bF$buf1),
    .C(_1265_),
    .D(_1148_),
    .Y(_874_)
);

INVX1 _7630_ (
    .A(\genblk1[1].u_ce.Ycalc [9]),
    .Y(_1266_)
);

INVX1 _7631_ (
    .A(_1258_),
    .Y(_1267_)
);

NOR2X1 _7632_ (
    .A(_1267_),
    .B(_1261_),
    .Y(_1268_)
);

INVX1 _7633_ (
    .A(\genblk1[1].u_ce.Yin12b [9]),
    .Y(_1269_)
);

OAI21X1 _7634_ (
    .A(1'h0),
    .B(_1180_),
    .C(_1249_),
    .Y(_1270_)
);

INVX1 _7635_ (
    .A(_1270_),
    .Y(_1271_)
);

OAI21X1 _7636_ (
    .A(_1250_),
    .B(_1248_),
    .C(_1119__bF$buf2),
    .Y(_1272_)
);

NAND2X1 _7637_ (
    .A(_1271_),
    .B(_1272_),
    .Y(_1273_)
);

NAND3X1 _7638_ (
    .A(_1228_),
    .B(_1252_),
    .C(_1231_),
    .Y(_1274_)
);

NAND3X1 _7639_ (
    .A(_1119__bF$buf1),
    .B(_1270_),
    .C(_1274_),
    .Y(_1275_)
);

NAND3X1 _7640_ (
    .A(_1269_),
    .B(_1273_),
    .C(_1275_),
    .Y(_1276_)
);

AND2X2 _7641_ (
    .A(_1272_),
    .B(_1271_),
    .Y(_1277_)
);

NOR2X1 _7642_ (
    .A(_1271_),
    .B(_1272_),
    .Y(_1278_)
);

OAI21X1 _7643_ (
    .A(_1278_),
    .B(_1277_),
    .C(\genblk1[1].u_ce.Yin12b [9]),
    .Y(_1279_)
);

NAND2X1 _7644_ (
    .A(_1276_),
    .B(_1279_),
    .Y(_1280_)
);

AOI21X1 _7645_ (
    .A(_1268_),
    .B(_1280_),
    .C(_1029_),
    .Y(_1281_)
);

OAI21X1 _7646_ (
    .A(_1268_),
    .B(_1280_),
    .C(_1281_),
    .Y(_1282_)
);

AOI22X1 _7647_ (
    .A(_1266_),
    .B(_1024__bF$buf0),
    .C(_1282_),
    .D(_1148_),
    .Y(_875_)
);

OAI21X1 _7648_ (
    .A(_1258_),
    .B(_1280_),
    .C(_1279_),
    .Y(_1283_)
);

NAND3X1 _7649_ (
    .A(_1276_),
    .B(_1279_),
    .C(_1259_),
    .Y(_1284_)
);

AOI21X1 _7650_ (
    .A(_1245_),
    .B(_1246_),
    .C(_1284_),
    .Y(_1285_)
);

INVX1 _7651_ (
    .A(\genblk1[1].u_ce.Yin12b [10]),
    .Y(_1286_)
);

OAI21X1 _7652_ (
    .A(1'h0),
    .B(_1203_),
    .C(_1249_),
    .Y(_1287_)
);

INVX1 _7653_ (
    .A(_1287_),
    .Y(_1288_)
);

OAI21X1 _7654_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1271_),
    .C(_1272_),
    .Y(_1289_)
);

NAND2X1 _7655_ (
    .A(_1288_),
    .B(_1289_),
    .Y(_1290_)
);

OAI21X1 _7656_ (
    .A(_1270_),
    .B(_1274_),
    .C(_1119__bF$buf0),
    .Y(_1291_)
);

NAND2X1 _7657_ (
    .A(_1287_),
    .B(_1291_),
    .Y(_1292_)
);

NAND2X1 _7658_ (
    .A(_1290_),
    .B(_1292_),
    .Y(_1293_)
);

NAND2X1 _7659_ (
    .A(_1286_),
    .B(_1293_),
    .Y(_1294_)
);

NAND3X1 _7660_ (
    .A(\genblk1[1].u_ce.Yin12b [10]),
    .B(_1290_),
    .C(_1292_),
    .Y(_1295_)
);

AND2X2 _7661_ (
    .A(_1294_),
    .B(_1295_),
    .Y(_1296_)
);

OAI21X1 _7662_ (
    .A(_1283_),
    .B(_1285_),
    .C(_1296_),
    .Y(_1297_)
);

INVX1 _7663_ (
    .A(_1279_),
    .Y(_1298_)
);

AOI21X1 _7664_ (
    .A(_1267_),
    .B(_1276_),
    .C(_1298_),
    .Y(_1299_)
);

AND2X2 _7665_ (
    .A(_1279_),
    .B(_1276_),
    .Y(_1300_)
);

NAND3X1 _7666_ (
    .A(_1259_),
    .B(_1300_),
    .C(_1263_),
    .Y(_1301_)
);

NAND2X1 _7667_ (
    .A(_1295_),
    .B(_1294_),
    .Y(_1302_)
);

NAND3X1 _7668_ (
    .A(_1299_),
    .B(_1302_),
    .C(_1301_),
    .Y(_1303_)
);

NAND3X1 _7669_ (
    .A(_1028_),
    .B(_1303_),
    .C(_1297_),
    .Y(_1304_)
);

AOI22X1 _7670_ (
    .A(_983_),
    .B(_1024__bF$buf4),
    .C(_1304_),
    .D(_1150_),
    .Y(_876_)
);

INVX1 _7671_ (
    .A(_1295_),
    .Y(_1305_)
);

AOI21X1 _7672_ (
    .A(_1301_),
    .B(_1299_),
    .C(_1302_),
    .Y(_1306_)
);

OAI21X1 _7673_ (
    .A(_1287_),
    .B(_1289_),
    .C(_1119__bF$buf5),
    .Y(_1307_)
);

INVX1 _7674_ (
    .A(_1307_),
    .Y(_1308_)
);

NAND2X1 _7675_ (
    .A(\genblk1[1].u_ce.Yin12b [11]),
    .B(_1178_),
    .Y(_1309_)
);

INVX1 _7676_ (
    .A(\genblk1[1].u_ce.Yin12b [11]),
    .Y(_1310_)
);

NAND2X1 _7677_ (
    .A(\genblk1[1].u_ce.Xin12b [11]),
    .B(_1310_),
    .Y(_1311_)
);

NAND2X1 _7678_ (
    .A(_1309_),
    .B(_1311_),
    .Y(_1312_)
);

OR2X2 _7679_ (
    .A(_1308_),
    .B(_1312_),
    .Y(_1313_)
);

NAND2X1 _7680_ (
    .A(_1312_),
    .B(_1308_),
    .Y(_1314_)
);

NAND2X1 _7681_ (
    .A(_1314_),
    .B(_1313_),
    .Y(_1315_)
);

OAI21X1 _7682_ (
    .A(_1305_),
    .B(_1306_),
    .C(_1315_),
    .Y(_1316_)
);

INVX1 _7683_ (
    .A(_1315_),
    .Y(_1317_)
);

NAND3X1 _7684_ (
    .A(_1295_),
    .B(_1317_),
    .C(_1297_),
    .Y(_1318_)
);

NAND3X1 _7685_ (
    .A(_1028_),
    .B(_1318_),
    .C(_1316_),
    .Y(_1319_)
);

AOI22X1 _7686_ (
    .A(_991_),
    .B(_1024__bF$buf3),
    .C(_1319_),
    .D(_1148_),
    .Y(_877_)
);

INVX1 _7687_ (
    .A(\genblk1[1].u_ce.Ycalc [0]),
    .Y(_1320_)
);

OAI21X1 _7688_ (
    .A(1'h0),
    .B(_1239_),
    .C(\genblk1[1].u_ce.Vld_bF$buf3 ),
    .Y(_1321_)
);

INVX2 _7689_ (
    .A(_1321_),
    .Y(_1322_)
);

INVX1 _7690_ (
    .A(\genblk1[1].u_ce.Yin0 [0]),
    .Y(_1323_)
);

AOI21X1 _7691_ (
    .A(_1090_),
    .B(_1097_),
    .C(_1323_),
    .Y(_1324_)
);

OAI21X1 _7692_ (
    .A(_1324_),
    .B(_1050_),
    .C(_1322_),
    .Y(_1325_)
);

OAI21X1 _7693_ (
    .A(_1320_),
    .B(\genblk1[1].u_ce.Vld_bF$buf2 ),
    .C(_1325_),
    .Y(_878_)
);

NAND2X1 _7694_ (
    .A(\genblk1[1].u_ce.Ycalc [1]),
    .B(_1024__bF$buf2),
    .Y(_1326_)
);

NAND3X1 _7695_ (
    .A(_1112_),
    .B(_1049_),
    .C(_1113_),
    .Y(_1327_)
);

OAI21X1 _7696_ (
    .A(_1111_),
    .B(_1051_),
    .C(_1050_),
    .Y(_1328_)
);

AOI21X1 _7697_ (
    .A(_1328_),
    .B(_1327_),
    .C(_1029_),
    .Y(_1329_)
);

OAI21X1 _7698_ (
    .A(_1024__bF$buf1),
    .B(_1329_),
    .C(_1326_),
    .Y(_879_)
);

NAND2X1 _7699_ (
    .A(\genblk1[1].u_ce.Xcalc [0]),
    .B(_1024__bF$buf0),
    .Y(_1330_)
);

MUX2X1 _7700_ (
    .A(\genblk1[1].u_ce.Yin12b [7]),
    .B(\genblk1[1].u_ce.Yin12b [6]),
    .S(1'h1),
    .Y(_1331_)
);

NAND2X1 _7701_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin12b [5]),
    .Y(_1332_)
);

OAI21X1 _7702_ (
    .A(1'h1),
    .B(_1151_),
    .C(_1332_),
    .Y(_1333_)
);

NAND2X1 _7703_ (
    .A(_1030__bF$buf4),
    .B(_1333_),
    .Y(_1334_)
);

OAI21X1 _7704_ (
    .A(_1030__bF$buf3),
    .B(_1331_),
    .C(_1334_),
    .Y(_1335_)
);

NAND2X1 _7705_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin1 [1]),
    .Y(_1336_)
);

OAI21X1 _7706_ (
    .A(1'h1),
    .B(_1053_),
    .C(_1336_),
    .Y(_1337_)
);

NAND2X1 _7707_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin0 [1]),
    .Y(_1338_)
);

OAI21X1 _7708_ (
    .A(1'h1),
    .B(_1323_),
    .C(_1338_),
    .Y(_1339_)
);

MUX2X1 _7709_ (
    .A(_1339_),
    .B(_1337_),
    .S(_1030__bF$buf2),
    .Y(_1340_)
);

NAND2X1 _7710_ (
    .A(_1057__bF$buf2),
    .B(_1340_),
    .Y(_1341_)
);

OAI21X1 _7711_ (
    .A(_1057__bF$buf1),
    .B(_1335_),
    .C(_1341_),
    .Y(_1342_)
);

INVX1 _7712_ (
    .A(_1342_),
    .Y(_1343_)
);

NOR2X1 _7713_ (
    .A(\genblk1[1].u_ce.Xin0 [0]),
    .B(_1343_),
    .Y(_1344_)
);

OAI21X1 _7714_ (
    .A(_1086_),
    .B(_1342_),
    .C(_1322_),
    .Y(_1345_)
);

OAI21X1 _7715_ (
    .A(_1345_),
    .B(_1344_),
    .C(_1330_),
    .Y(_880_)
);

NAND2X1 _7716_ (
    .A(\genblk1[1].u_ce.Xcalc [1]),
    .B(_1024__bF$buf4),
    .Y(_1346_)
);

NOR2X1 _7717_ (
    .A(_1086_),
    .B(_1342_),
    .Y(_1347_)
);

NAND2X1 _7718_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin12b [4]),
    .Y(_1348_)
);

OAI21X1 _7719_ (
    .A(1'h1),
    .B(_1141_),
    .C(_1348_),
    .Y(_1349_)
);

NAND2X1 _7720_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin1 [0]),
    .Y(_1350_)
);

OAI21X1 _7721_ (
    .A(1'h1),
    .B(_1108_),
    .C(_1350_),
    .Y(_1351_)
);

MUX2X1 _7722_ (
    .A(_1351_),
    .B(_1349_),
    .S(_1030__bF$buf1),
    .Y(_1352_)
);

NAND2X1 _7723_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin12b [8]),
    .Y(_1353_)
);

OAI21X1 _7724_ (
    .A(1'h1),
    .B(_1225_),
    .C(_1353_),
    .Y(_1354_)
);

NAND2X1 _7725_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin12b [6]),
    .Y(_1355_)
);

OAI21X1 _7726_ (
    .A(1'h1),
    .B(_1176_),
    .C(_1355_),
    .Y(_1356_)
);

MUX2X1 _7727_ (
    .A(_1356_),
    .B(_1354_),
    .S(_1030__bF$buf0),
    .Y(_1357_)
);

MUX2X1 _7728_ (
    .A(_1357_),
    .B(_1352_),
    .S(1'h0),
    .Y(_1358_)
);

NOR2X1 _7729_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf4 ),
    .B(_1342_),
    .Y(_1359_)
);

NAND2X1 _7730_ (
    .A(_1358_),
    .B(_1359_),
    .Y(_1360_)
);

NAND2X1 _7731_ (
    .A(_1057__bF$buf0),
    .B(_1352_),
    .Y(_1361_)
);

NAND2X1 _7732_ (
    .A(1'h0),
    .B(_1357_),
    .Y(_1362_)
);

NAND2X1 _7733_ (
    .A(_1361_),
    .B(_1362_),
    .Y(_1363_)
);

OAI21X1 _7734_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1342_),
    .C(_1363_),
    .Y(_1364_)
);

NAND3X1 _7735_ (
    .A(\genblk1[1].u_ce.Xin0 [1]),
    .B(_1364_),
    .C(_1360_),
    .Y(_1365_)
);

OAI21X1 _7736_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1342_),
    .C(_1358_),
    .Y(_1366_)
);

NAND2X1 _7737_ (
    .A(_1363_),
    .B(_1359_),
    .Y(_1367_)
);

NAND3X1 _7738_ (
    .A(_1066_),
    .B(_1366_),
    .C(_1367_),
    .Y(_1368_)
);

NAND3X1 _7739_ (
    .A(_1347_),
    .B(_1365_),
    .C(_1368_),
    .Y(_1369_)
);

INVX1 _7740_ (
    .A(_1347_),
    .Y(_1370_)
);

AOI21X1 _7741_ (
    .A(_1367_),
    .B(_1366_),
    .C(_1066_),
    .Y(_1371_)
);

AOI21X1 _7742_ (
    .A(_1360_),
    .B(_1364_),
    .C(\genblk1[1].u_ce.Xin0 [1]),
    .Y(_1372_)
);

OAI21X1 _7743_ (
    .A(_1371_),
    .B(_1372_),
    .C(_1370_),
    .Y(_1373_)
);

AOI21X1 _7744_ (
    .A(_1373_),
    .B(_1369_),
    .C(_1029_),
    .Y(_1374_)
);

OAI21X1 _7745_ (
    .A(_1024__bF$buf3),
    .B(_1374_),
    .C(_1346_),
    .Y(_881_)
);

OAI21X1 _7746_ (
    .A(_1370_),
    .B(_1372_),
    .C(_1365_),
    .Y(_1375_)
);

MUX2X1 _7747_ (
    .A(\genblk1[1].u_ce.Yin12b [9]),
    .B(\genblk1[1].u_ce.Yin12b [8]),
    .S(1'h1),
    .Y(_1376_)
);

MUX2X1 _7748_ (
    .A(_1376_),
    .B(_1331_),
    .S(1'h0),
    .Y(_1377_)
);

NOR2X1 _7749_ (
    .A(1'h0),
    .B(_1030__bF$buf4),
    .Y(_1378_)
);

NAND2X1 _7750_ (
    .A(_1333_),
    .B(_1378_),
    .Y(_1379_)
);

NAND2X1 _7751_ (
    .A(_1027_),
    .B(_1337_),
    .Y(_1380_)
);

NAND2X1 _7752_ (
    .A(_1380_),
    .B(_1379_),
    .Y(_1381_)
);

AOI21X1 _7753_ (
    .A(1'h0),
    .B(_1377_),
    .C(_1381_),
    .Y(_1382_)
);

NAND2X1 _7754_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin12b [7]),
    .Y(_1383_)
);

OAI21X1 _7755_ (
    .A(1'h1),
    .B(_1200_),
    .C(_1383_),
    .Y(_1384_)
);

MUX2X1 _7756_ (
    .A(_1333_),
    .B(_1384_),
    .S(_1030__bF$buf3),
    .Y(_1385_)
);

NAND2X1 _7757_ (
    .A(1'h0),
    .B(_1385_),
    .Y(_1386_)
);

AOI21X1 _7758_ (
    .A(_1341_),
    .B(_1386_),
    .C(_1358_),
    .Y(_1387_)
);

NOR2X1 _7759_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1387_),
    .Y(_1388_)
);

NAND2X1 _7760_ (
    .A(_1382_),
    .B(_1388_),
    .Y(_1389_)
);

INVX1 _7761_ (
    .A(_1382_),
    .Y(_1390_)
);

OAI21X1 _7762_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1387_),
    .C(_1390_),
    .Y(_1391_)
);

AOI21X1 _7763_ (
    .A(_1389_),
    .B(_1391_),
    .C(_1082_),
    .Y(_1392_)
);

NAND3X1 _7764_ (
    .A(_1082_),
    .B(_1391_),
    .C(_1389_),
    .Y(_1393_)
);

INVX1 _7765_ (
    .A(_1393_),
    .Y(_1394_)
);

NOR2X1 _7766_ (
    .A(_1392_),
    .B(_1394_),
    .Y(_1395_)
);

NOR2X1 _7767_ (
    .A(_1375_),
    .B(_1395_),
    .Y(_1396_)
);

AOI21X1 _7768_ (
    .A(_1347_),
    .B(_1368_),
    .C(_1371_),
    .Y(_1397_)
);

INVX1 _7769_ (
    .A(_1395_),
    .Y(_1398_)
);

OAI21X1 _7770_ (
    .A(_1397_),
    .B(_1398_),
    .C(_1322_),
    .Y(_1399_)
);

OAI22X1 _7771_ (
    .A(_999_),
    .B(\genblk1[1].u_ce.Vld_bF$buf1 ),
    .C(_1396_),
    .D(_1399_),
    .Y(_882_)
);

NAND2X1 _7772_ (
    .A(\genblk1[1].u_ce.Xcalc [3]),
    .B(_1024__bF$buf2),
    .Y(_1400_)
);

AOI21X1 _7773_ (
    .A(_1375_),
    .B(_1393_),
    .C(_1392_),
    .Y(_1401_)
);

NAND2X1 _7774_ (
    .A(1'h1),
    .B(_1286_),
    .Y(_1402_)
);

OAI21X1 _7775_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin12b [9]),
    .C(_1402_),
    .Y(_1403_)
);

NAND2X1 _7776_ (
    .A(_1030__bF$buf2),
    .B(_1354_),
    .Y(_1404_)
);

OAI21X1 _7777_ (
    .A(_1030__bF$buf1),
    .B(_1403_),
    .C(_1404_),
    .Y(_1405_)
);

NAND2X1 _7778_ (
    .A(_1356_),
    .B(_1378_),
    .Y(_1406_)
);

NAND2X1 _7779_ (
    .A(_1027_),
    .B(_1349_),
    .Y(_1407_)
);

NAND2X1 _7780_ (
    .A(_1407_),
    .B(_1406_),
    .Y(_1408_)
);

AOI21X1 _7781_ (
    .A(_1405_),
    .B(1'h0),
    .C(_1408_),
    .Y(_1409_)
);

NAND3X1 _7782_ (
    .A(_1382_),
    .B(_1363_),
    .C(_1342_),
    .Y(_1410_)
);

NAND2X1 _7783_ (
    .A(_1119__bF$buf4),
    .B(_1410_),
    .Y(_1411_)
);

OR2X2 _7784_ (
    .A(_1411_),
    .B(_1409_),
    .Y(_1412_)
);

INVX1 _7785_ (
    .A(_1410_),
    .Y(_1413_)
);

OAI21X1 _7786_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf4 ),
    .B(_1413_),
    .C(_1409_),
    .Y(_1414_)
);

NAND3X1 _7787_ (
    .A(\genblk1[1].u_ce.Xin1 [1]),
    .B(_1414_),
    .C(_1412_),
    .Y(_1415_)
);

INVX1 _7788_ (
    .A(_1409_),
    .Y(_1416_)
);

OR2X2 _7789_ (
    .A(_1411_),
    .B(_1416_),
    .Y(_1417_)
);

OAI21X1 _7790_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1413_),
    .C(_1416_),
    .Y(_1418_)
);

NAND3X1 _7791_ (
    .A(_1061_),
    .B(_1418_),
    .C(_1417_),
    .Y(_1419_)
);

NAND2X1 _7792_ (
    .A(_1415_),
    .B(_1419_),
    .Y(_1420_)
);

OR2X2 _7793_ (
    .A(_1401_),
    .B(_1420_),
    .Y(_1421_)
);

NAND2X1 _7794_ (
    .A(_1420_),
    .B(_1401_),
    .Y(_1422_)
);

AOI21X1 _7795_ (
    .A(_1421_),
    .B(_1422_),
    .C(_1029_),
    .Y(_1423_)
);

OAI21X1 _7796_ (
    .A(_1024__bF$buf1),
    .B(_1423_),
    .C(_1400_),
    .Y(_883_)
);

OAI21X1 _7797_ (
    .A(_1420_),
    .B(_1401_),
    .C(_1415_),
    .Y(_1424_)
);

NAND2X1 _7798_ (
    .A(1'h1),
    .B(\genblk1[1].u_ce.Yin12b [11]),
    .Y(_1425_)
);

OAI21X1 _7799_ (
    .A(1'h1),
    .B(_1286_),
    .C(_1425_),
    .Y(_1426_)
);

NAND2X1 _7800_ (
    .A(1'h0),
    .B(_1426_),
    .Y(_1427_)
);

OAI21X1 _7801_ (
    .A(1'h0),
    .B(_1376_),
    .C(_1427_),
    .Y(_1428_)
);

NAND2X1 _7802_ (
    .A(1'h0),
    .B(_1428_),
    .Y(_1429_)
);

OAI21X1 _7803_ (
    .A(1'h0),
    .B(_1385_),
    .C(_1429_),
    .Y(_1430_)
);

INVX1 _7804_ (
    .A(_1430_),
    .Y(_1431_)
);

OAI21X1 _7805_ (
    .A(_1416_),
    .B(_1410_),
    .C(_1119__bF$buf3),
    .Y(_1432_)
);

OR2X2 _7806_ (
    .A(_1432_),
    .B(_1431_),
    .Y(_1433_)
);

NAND2X1 _7807_ (
    .A(_1431_),
    .B(_1432_),
    .Y(_1434_)
);

NAND3X1 _7808_ (
    .A(\genblk1[1].u_ce.Xin12b [4]),
    .B(_1434_),
    .C(_1433_),
    .Y(_1435_)
);

OR2X2 _7809_ (
    .A(_1432_),
    .B(_1430_),
    .Y(_1436_)
);

NAND2X1 _7810_ (
    .A(_1430_),
    .B(_1432_),
    .Y(_1437_)
);

NAND3X1 _7811_ (
    .A(_1063_),
    .B(_1437_),
    .C(_1436_),
    .Y(_1438_)
);

AND2X2 _7812_ (
    .A(_1435_),
    .B(_1438_),
    .Y(_1439_)
);

NAND2X1 _7813_ (
    .A(_1439_),
    .B(_1424_),
    .Y(_1440_)
);

INVX1 _7814_ (
    .A(_1392_),
    .Y(_1441_)
);

OAI21X1 _7815_ (
    .A(_1394_),
    .B(_1397_),
    .C(_1441_),
    .Y(_1442_)
);

INVX1 _7816_ (
    .A(_1415_),
    .Y(_1443_)
);

AOI21X1 _7817_ (
    .A(_1442_),
    .B(_1419_),
    .C(_1443_),
    .Y(_1444_)
);

NAND2X1 _7818_ (
    .A(_1438_),
    .B(_1435_),
    .Y(_1445_)
);

NAND2X1 _7819_ (
    .A(_1445_),
    .B(_1444_),
    .Y(_1446_)
);

NAND2X1 _7820_ (
    .A(_1440_),
    .B(_1446_),
    .Y(_1447_)
);

AOI22X1 _7821_ (
    .A(_1001_),
    .B(_1024__bF$buf0),
    .C(_1447_),
    .D(_1322_),
    .Y(_884_)
);

NAND3X1 _7822_ (
    .A(_1409_),
    .B(_1431_),
    .C(_1413_),
    .Y(_1448_)
);

NOR2X1 _7823_ (
    .A(1'h0),
    .B(_1403_),
    .Y(_1449_)
);

NOR2X1 _7824_ (
    .A(_1030__bF$buf0),
    .B(_1310_),
    .Y(_1450_)
);

OAI21X1 _7825_ (
    .A(_1450_),
    .B(_1449_),
    .C(1'h0),
    .Y(_1451_)
);

OAI21X1 _7826_ (
    .A(1'h0),
    .B(_1357_),
    .C(_1451_),
    .Y(_1452_)
);

NAND3X1 _7827_ (
    .A(_1119__bF$buf2),
    .B(_1452_),
    .C(_1448_),
    .Y(_1453_)
);

INVX1 _7828_ (
    .A(_1452_),
    .Y(_1454_)
);

NAND3X1 _7829_ (
    .A(_1382_),
    .B(_1409_),
    .C(_1387_),
    .Y(_1455_)
);

OAI21X1 _7830_ (
    .A(_1430_),
    .B(_1455_),
    .C(_1119__bF$buf1),
    .Y(_1456_)
);

NAND2X1 _7831_ (
    .A(_1454_),
    .B(_1456_),
    .Y(_1457_)
);

NAND3X1 _7832_ (
    .A(\genblk1[1].u_ce.Xin12b [5]),
    .B(_1457_),
    .C(_1453_),
    .Y(_1458_)
);

NAND3X1 _7833_ (
    .A(_1119__bF$buf0),
    .B(_1454_),
    .C(_1448_),
    .Y(_1459_)
);

NAND2X1 _7834_ (
    .A(_1452_),
    .B(_1456_),
    .Y(_1460_)
);

NAND3X1 _7835_ (
    .A(_1071_),
    .B(_1460_),
    .C(_1459_),
    .Y(_1461_)
);

NAND2X1 _7836_ (
    .A(_1458_),
    .B(_1461_),
    .Y(_1462_)
);

AOI21X1 _7837_ (
    .A(_1440_),
    .B(_1435_),
    .C(_1462_),
    .Y(_1463_)
);

OAI21X1 _7838_ (
    .A(_1445_),
    .B(_1444_),
    .C(_1435_),
    .Y(_1464_)
);

AND2X2 _7839_ (
    .A(_1458_),
    .B(_1461_),
    .Y(_1465_)
);

OAI21X1 _7840_ (
    .A(_1465_),
    .B(_1464_),
    .C(_1322_),
    .Y(_1466_)
);

OAI22X1 _7841_ (
    .A(_1016_),
    .B(\genblk1[1].u_ce.Vld_bF$buf0 ),
    .C(_1463_),
    .D(_1466_),
    .Y(_885_)
);

NOR2X1 _7842_ (
    .A(_1430_),
    .B(_1455_),
    .Y(_1467_)
);

NAND2X1 _7843_ (
    .A(_1454_),
    .B(_1467_),
    .Y(_1468_)
);

AOI21X1 _7844_ (
    .A(_1030__bF$buf4),
    .B(_1426_),
    .C(_1450_),
    .Y(_1469_)
);

NAND2X1 _7845_ (
    .A(_1057__bF$buf3),
    .B(_1377_),
    .Y(_1470_)
);

OAI21X1 _7846_ (
    .A(_1057__bF$buf2),
    .B(_1469_),
    .C(_1470_),
    .Y(_1471_)
);

NAND3X1 _7847_ (
    .A(_1119__bF$buf5),
    .B(_1471_),
    .C(_1468_),
    .Y(_1472_)
);

NOR3X1 _7848_ (
    .A(_1430_),
    .B(_1452_),
    .C(_1455_),
    .Y(_1473_)
);

INVX1 _7849_ (
    .A(_1471_),
    .Y(_1474_)
);

OAI21X1 _7850_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1473_),
    .C(_1474_),
    .Y(_1475_)
);

NAND3X1 _7851_ (
    .A(\genblk1[1].u_ce.Xin12b [6]),
    .B(_1475_),
    .C(_1472_),
    .Y(_1476_)
);

NAND3X1 _7852_ (
    .A(_1119__bF$buf4),
    .B(_1474_),
    .C(_1468_),
    .Y(_1477_)
);

OAI21X1 _7853_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1473_),
    .C(_1471_),
    .Y(_1478_)
);

NAND3X1 _7854_ (
    .A(_1073_),
    .B(_1478_),
    .C(_1477_),
    .Y(_1479_)
);

AND2X2 _7855_ (
    .A(_1476_),
    .B(_1479_),
    .Y(_1480_)
);

NAND2X1 _7856_ (
    .A(_1439_),
    .B(_1465_),
    .Y(_1481_)
);

INVX1 _7857_ (
    .A(_1435_),
    .Y(_1482_)
);

INVX1 _7858_ (
    .A(_1458_),
    .Y(_1483_)
);

AOI21X1 _7859_ (
    .A(_1482_),
    .B(_1461_),
    .C(_1483_),
    .Y(_1484_)
);

OAI21X1 _7860_ (
    .A(_1444_),
    .B(_1481_),
    .C(_1484_),
    .Y(_1485_)
);

AND2X2 _7861_ (
    .A(_1485_),
    .B(_1480_),
    .Y(_1486_)
);

NOR2X1 _7862_ (
    .A(_1480_),
    .B(_1485_),
    .Y(_1487_)
);

OAI21X1 _7863_ (
    .A(_1487_),
    .B(_1486_),
    .C(_1028_),
    .Y(_1488_)
);

NAND2X1 _7864_ (
    .A(\genblk1[1].u_ce.Vld_bF$buf4 ),
    .B(_1488_),
    .Y(_1489_)
);

OAI21X1 _7865_ (
    .A(_1002_),
    .B(\genblk1[1].u_ce.Vld_bF$buf3 ),
    .C(_1489_),
    .Y(_886_)
);

INVX1 _7866_ (
    .A(_1476_),
    .Y(_1490_)
);

NOR2X1 _7867_ (
    .A(_1490_),
    .B(_1486_),
    .Y(_1491_)
);

NAND2X1 _7868_ (
    .A(_1474_),
    .B(_1473_),
    .Y(_1492_)
);

NOR2X1 _7869_ (
    .A(_1057__bF$buf1),
    .B(_1310_),
    .Y(_1493_)
);

AOI21X1 _7870_ (
    .A(_1405_),
    .B(_1057__bF$buf0),
    .C(_1493_),
    .Y(_1494_)
);

NAND3X1 _7871_ (
    .A(_1119__bF$buf3),
    .B(_1494_),
    .C(_1492_),
    .Y(_1495_)
);

INVX1 _7872_ (
    .A(_1495_),
    .Y(_1496_)
);

AOI21X1 _7873_ (
    .A(_1492_),
    .B(_1119__bF$buf2),
    .C(_1494_),
    .Y(_1497_)
);

OAI21X1 _7874_ (
    .A(_1497_),
    .B(_1496_),
    .C(\genblk1[1].u_ce.Xin12b [7]),
    .Y(_1498_)
);

INVX1 _7875_ (
    .A(_1497_),
    .Y(_1499_)
);

NAND3X1 _7876_ (
    .A(_1076_),
    .B(_1495_),
    .C(_1499_),
    .Y(_1500_)
);

AND2X2 _7877_ (
    .A(_1500_),
    .B(_1498_),
    .Y(_1501_)
);

OR2X2 _7878_ (
    .A(_1491_),
    .B(_1501_),
    .Y(_1502_)
);

AOI21X1 _7879_ (
    .A(_1491_),
    .B(_1501_),
    .C(_1321_),
    .Y(_1503_)
);

AOI22X1 _7880_ (
    .A(_1015_),
    .B(_1024__bF$buf4),
    .C(_1502_),
    .D(_1503_),
    .Y(_887_)
);

NOR2X1 _7881_ (
    .A(_1445_),
    .B(_1462_),
    .Y(_1504_)
);

OAI21X1 _7882_ (
    .A(_1435_),
    .B(_1462_),
    .C(_1458_),
    .Y(_1505_)
);

AOI21X1 _7883_ (
    .A(_1504_),
    .B(_1424_),
    .C(_1505_),
    .Y(_1506_)
);

AOI21X1 _7884_ (
    .A(_1499_),
    .B(_1495_),
    .C(_1076_),
    .Y(_1507_)
);

AOI21X1 _7885_ (
    .A(_1490_),
    .B(_1500_),
    .C(_1507_),
    .Y(_1508_)
);

NAND3X1 _7886_ (
    .A(_1480_),
    .B(_1498_),
    .C(_1500_),
    .Y(_1509_)
);

OAI21X1 _7887_ (
    .A(_1509_),
    .B(_1506_),
    .C(_1508_),
    .Y(_1510_)
);

NAND3X1 _7888_ (
    .A(_1474_),
    .B(_1494_),
    .C(_1473_),
    .Y(_1511_)
);

INVX1 _7889_ (
    .A(_1428_),
    .Y(_1512_)
);

INVX1 _7890_ (
    .A(_1493_),
    .Y(_1513_)
);

OAI21X1 _7891_ (
    .A(1'h0),
    .B(_1512_),
    .C(_1513_),
    .Y(_1514_)
);

INVX1 _7892_ (
    .A(_1514_),
    .Y(_1515_)
);

NAND3X1 _7893_ (
    .A(_1119__bF$buf1),
    .B(_1515_),
    .C(_1511_),
    .Y(_1516_)
);

INVX1 _7894_ (
    .A(_1516_),
    .Y(_1517_)
);

AOI21X1 _7895_ (
    .A(_1511_),
    .B(_1119__bF$buf0),
    .C(_1515_),
    .Y(_1518_)
);

OAI21X1 _7896_ (
    .A(_1518_),
    .B(_1517_),
    .C(\genblk1[1].u_ce.Xin12b [8]),
    .Y(_1519_)
);

INVX1 _7897_ (
    .A(_1518_),
    .Y(_1520_)
);

NAND3X1 _7898_ (
    .A(_1078_),
    .B(_1516_),
    .C(_1520_),
    .Y(_1521_)
);

AND2X2 _7899_ (
    .A(_1521_),
    .B(_1519_),
    .Y(_1522_)
);

OR2X2 _7900_ (
    .A(_1510_),
    .B(_1522_),
    .Y(_1523_)
);

INVX1 _7901_ (
    .A(_1523_),
    .Y(_1524_)
);

NAND2X1 _7902_ (
    .A(_1522_),
    .B(_1510_),
    .Y(_1525_)
);

NAND2X1 _7903_ (
    .A(_1322_),
    .B(_1525_),
    .Y(_1526_)
);

OAI22X1 _7904_ (
    .A(_1004_),
    .B(\genblk1[1].u_ce.Vld_bF$buf2 ),
    .C(_1526_),
    .D(_1524_),
    .Y(_888_)
);

NOR3X1 _7905_ (
    .A(_1452_),
    .B(_1471_),
    .C(_1448_),
    .Y(_1527_)
);

NAND3X1 _7906_ (
    .A(_1494_),
    .B(_1515_),
    .C(_1527_),
    .Y(_1528_)
);

OR2X2 _7907_ (
    .A(_1449_),
    .B(_1450_),
    .Y(_1529_)
);

AOI21X1 _7908_ (
    .A(_1529_),
    .B(_1057__bF$buf3),
    .C(_1493_),
    .Y(_1530_)
);

INVX1 _7909_ (
    .A(_1530_),
    .Y(_1531_)
);

NAND3X1 _7910_ (
    .A(_1119__bF$buf5),
    .B(_1531_),
    .C(_1528_),
    .Y(_1532_)
);

OAI21X1 _7911_ (
    .A(_1514_),
    .B(_1511_),
    .C(_1119__bF$buf4),
    .Y(_1533_)
);

NAND2X1 _7912_ (
    .A(_1530_),
    .B(_1533_),
    .Y(_1534_)
);

NAND3X1 _7913_ (
    .A(\genblk1[1].u_ce.Xin12b [9]),
    .B(_1534_),
    .C(_1532_),
    .Y(_1535_)
);

NAND3X1 _7914_ (
    .A(_1119__bF$buf3),
    .B(_1530_),
    .C(_1528_),
    .Y(_1536_)
);

NAND2X1 _7915_ (
    .A(_1531_),
    .B(_1533_),
    .Y(_1537_)
);

NAND3X1 _7916_ (
    .A(_1123_),
    .B(_1537_),
    .C(_1536_),
    .Y(_1538_)
);

NAND2X1 _7917_ (
    .A(_1535_),
    .B(_1538_),
    .Y(_1539_)
);

AOI21X1 _7918_ (
    .A(_1525_),
    .B(_1519_),
    .C(_1539_),
    .Y(_1540_)
);

NAND3X1 _7919_ (
    .A(_1519_),
    .B(_1539_),
    .C(_1525_),
    .Y(_1541_)
);

NAND2X1 _7920_ (
    .A(_1322_),
    .B(_1541_),
    .Y(_1542_)
);

OAI22X1 _7921_ (
    .A(_1012_),
    .B(\genblk1[1].u_ce.Vld_bF$buf1 ),
    .C(_1540_),
    .D(_1542_),
    .Y(_889_)
);

NAND2X1 _7922_ (
    .A(\genblk1[1].u_ce.Xcalc [10]),
    .B(_1024__bF$buf3),
    .Y(_1543_)
);

OAI21X1 _7923_ (
    .A(1'h0),
    .B(_1469_),
    .C(_1513_),
    .Y(_1544_)
);

OAI21X1 _7924_ (
    .A(_1531_),
    .B(_1528_),
    .C(_1119__bF$buf2),
    .Y(_1545_)
);

NOR2X1 _7925_ (
    .A(_1544_),
    .B(_1545_),
    .Y(_1546_)
);

NAND2X1 _7926_ (
    .A(_1544_),
    .B(_1545_),
    .Y(_1547_)
);

INVX1 _7927_ (
    .A(_1547_),
    .Y(_1548_)
);

OAI21X1 _7928_ (
    .A(_1546_),
    .B(_1548_),
    .C(\genblk1[1].u_ce.Xin12b [10]),
    .Y(_1549_)
);

INVX1 _7929_ (
    .A(_1546_),
    .Y(_1550_)
);

NAND3X1 _7930_ (
    .A(_1153_),
    .B(_1547_),
    .C(_1550_),
    .Y(_1551_)
);

AND2X2 _7931_ (
    .A(_1551_),
    .B(_1549_),
    .Y(_1552_)
);

OAI21X1 _7932_ (
    .A(_1519_),
    .B(_1539_),
    .C(_1535_),
    .Y(_1553_)
);

NAND3X1 _7933_ (
    .A(_1480_),
    .B(_1485_),
    .C(_1501_),
    .Y(_1554_)
);

NAND3X1 _7934_ (
    .A(_1535_),
    .B(_1538_),
    .C(_1522_),
    .Y(_1555_)
);

AOI21X1 _7935_ (
    .A(_1554_),
    .B(_1508_),
    .C(_1555_),
    .Y(_1556_)
);

OAI21X1 _7936_ (
    .A(_1553_),
    .B(_1556_),
    .C(_1552_),
    .Y(_1557_)
);

NAND2X1 _7937_ (
    .A(_1549_),
    .B(_1551_),
    .Y(_1558_)
);

NAND2X1 _7938_ (
    .A(_1519_),
    .B(_1521_),
    .Y(_1559_)
);

NOR2X1 _7939_ (
    .A(_1559_),
    .B(_1539_),
    .Y(_1560_)
);

AOI21X1 _7940_ (
    .A(_1510_),
    .B(_1560_),
    .C(_1553_),
    .Y(_1561_)
);

NAND2X1 _7941_ (
    .A(_1558_),
    .B(_1561_),
    .Y(_1562_)
);

AOI21X1 _7942_ (
    .A(_1557_),
    .B(_1562_),
    .C(_1029_),
    .Y(_1563_)
);

OAI21X1 _7943_ (
    .A(_1024__bF$buf2),
    .B(_1563_),
    .C(_1543_),
    .Y(_890_)
);

NAND2X1 _7944_ (
    .A(\genblk1[1].u_ce.Xcalc [11]),
    .B(_1024__bF$buf1),
    .Y(_1564_)
);

OR2X2 _7945_ (
    .A(_1528_),
    .B(_1531_),
    .Y(_1565_)
);

OAI21X1 _7946_ (
    .A(_1544_),
    .B(_1565_),
    .C(_1119__bF$buf1),
    .Y(_1566_)
);

OR2X2 _7947_ (
    .A(_1566_),
    .B(_1312_),
    .Y(_1567_)
);

NAND2X1 _7948_ (
    .A(_1312_),
    .B(_1566_),
    .Y(_1568_)
);

AOI22X1 _7949_ (
    .A(_1567_),
    .B(_1568_),
    .C(_1557_),
    .D(_1549_),
    .Y(_1569_)
);

OAI21X1 _7950_ (
    .A(_1558_),
    .B(_1561_),
    .C(_1549_),
    .Y(_1570_)
);

NAND2X1 _7951_ (
    .A(_1568_),
    .B(_1567_),
    .Y(_1571_)
);

OAI21X1 _7952_ (
    .A(_1571_),
    .B(_1570_),
    .C(_1322_),
    .Y(_1572_)
);

OAI21X1 _7953_ (
    .A(_1569_),
    .B(_1572_),
    .C(_1564_),
    .Y(_891_)
);

NAND2X1 _7954_ (
    .A(1'h1),
    .B(1'h0),
    .Y(_1573_)
);

OAI21X1 _7955_ (
    .A(_1057__bF$buf2),
    .B(_1239_),
    .C(_1573_),
    .Y(_1574_)
);

NOR2X1 _7956_ (
    .A(_1020_),
    .B(_1574_),
    .Y(_1575_)
);

AND2X2 _7957_ (
    .A(_1574_),
    .B(_1020_),
    .Y(_1576_)
);

OR2X2 _7958_ (
    .A(_1576_),
    .B(_1575_),
    .Y(_1577_)
);

NAND2X1 _7959_ (
    .A(\genblk1[1].u_ce.Acalc [0]),
    .B(_1024__bF$buf0),
    .Y(_1578_)
);

OAI21X1 _7960_ (
    .A(_1024__bF$buf4),
    .B(_1577_),
    .C(_1578_),
    .Y(_892_)
);

NAND2X1 _7961_ (
    .A(\genblk1[1].u_ce.Acalc [1]),
    .B(_1024__bF$buf3),
    .Y(_1579_)
);

OAI21X1 _7962_ (
    .A(1'h0),
    .B(_1026_),
    .C(1'h0),
    .Y(_1580_)
);

OAI21X1 _7963_ (
    .A(1'h0),
    .B(_1026_),
    .C(_1580_),
    .Y(_1581_)
);

OAI21X1 _7964_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1574_),
    .C(_1581_),
    .Y(_1582_)
);

OAI21X1 _7965_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf4 ),
    .B(_1581_),
    .C(_1582_),
    .Y(_1583_)
);

OR2X2 _7966_ (
    .A(_1583_),
    .B(\genblk1[1].u_ce.Ain0 [1]),
    .Y(_1584_)
);

NAND2X1 _7967_ (
    .A(\genblk1[1].u_ce.Ain0 [1]),
    .B(_1583_),
    .Y(_1585_)
);

NAND2X1 _7968_ (
    .A(_1585_),
    .B(_1584_),
    .Y(_1586_)
);

NOR2X1 _7969_ (
    .A(_1575_),
    .B(_1586_),
    .Y(_1587_)
);

NAND2X1 _7970_ (
    .A(_1575_),
    .B(_1586_),
    .Y(_1588_)
);

NAND2X1 _7971_ (
    .A(\genblk1[1].u_ce.Vld_bF$buf0 ),
    .B(_1588_),
    .Y(_1589_)
);

OAI21X1 _7972_ (
    .A(_1587_),
    .B(_1589_),
    .C(_1579_),
    .Y(_893_)
);

NAND2X1 _7973_ (
    .A(\genblk1[1].u_ce.Acalc [2]),
    .B(_1024__bF$buf2),
    .Y(_1590_)
);

OAI21X1 _7974_ (
    .A(_1022_),
    .B(_1583_),
    .C(_1588_),
    .Y(_1591_)
);

OAI21X1 _7975_ (
    .A(_1026_),
    .B(_1030__bF$buf3),
    .C(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_1592_)
);

NAND3X1 _7976_ (
    .A(1'h0),
    .B(_1239_),
    .C(_1592_),
    .Y(_1593_)
);

OAI21X1 _7977_ (
    .A(1'h0),
    .B(_1592_),
    .C(_1593_),
    .Y(_1594_)
);

NAND2X1 _7978_ (
    .A(\genblk1[1].u_ce.Ain1 [0]),
    .B(_1594_),
    .Y(_1595_)
);

OR2X2 _7979_ (
    .A(_1594_),
    .B(\genblk1[1].u_ce.Ain1 [0]),
    .Y(_1596_)
);

NAND2X1 _7980_ (
    .A(_1595_),
    .B(_1596_),
    .Y(_1597_)
);

INVX1 _7981_ (
    .A(_1597_),
    .Y(_1598_)
);

NOR2X1 _7982_ (
    .A(_1598_),
    .B(_1591_),
    .Y(_1599_)
);

NAND2X1 _7983_ (
    .A(_1598_),
    .B(_1591_),
    .Y(_1600_)
);

NAND2X1 _7984_ (
    .A(\genblk1[1].u_ce.Vld_bF$buf4 ),
    .B(_1600_),
    .Y(_1601_)
);

OAI21X1 _7985_ (
    .A(_1599_),
    .B(_1601_),
    .C(_1590_),
    .Y(_894_)
);

NAND2X1 _7986_ (
    .A(_1595_),
    .B(_1600_),
    .Y(_1602_)
);

INVX1 _7987_ (
    .A(_1602_),
    .Y(_1603_)
);

INVX1 _7988_ (
    .A(\genblk1[1].u_ce.Ain1 [1]),
    .Y(_1604_)
);

OAI21X1 _7989_ (
    .A(1'h1),
    .B(_1030__bF$buf2),
    .C(1'h0),
    .Y(_1605_)
);

NAND2X1 _7990_ (
    .A(_1119__bF$buf0),
    .B(_1605_),
    .Y(_1606_)
);

OAI21X1 _7991_ (
    .A(1'h0),
    .B(1'h0),
    .C(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .Y(_1607_)
);

OAI21X1 _7992_ (
    .A(_1026_),
    .B(_1607_),
    .C(_1606_),
    .Y(_1608_)
);

NOR2X1 _7993_ (
    .A(_1604_),
    .B(_1608_),
    .Y(_1609_)
);

NAND2X1 _7994_ (
    .A(_1604_),
    .B(_1608_),
    .Y(_1610_)
);

INVX1 _7995_ (
    .A(_1610_),
    .Y(_1611_)
);

OAI21X1 _7996_ (
    .A(_1609_),
    .B(_1611_),
    .C(_1603_),
    .Y(_1612_)
);

INVX1 _7997_ (
    .A(_1609_),
    .Y(_1613_)
);

NAND3X1 _7998_ (
    .A(_1613_),
    .B(_1610_),
    .C(_1602_),
    .Y(_1614_)
);

NAND2X1 _7999_ (
    .A(_1614_),
    .B(_1612_),
    .Y(_1615_)
);

NAND2X1 _8000_ (
    .A(\genblk1[1].u_ce.Acalc [3]),
    .B(_1024__bF$buf1),
    .Y(_1616_)
);

OAI21X1 _8001_ (
    .A(_1024__bF$buf0),
    .B(_1615_),
    .C(_1616_),
    .Y(_895_)
);

NOR2X1 _8002_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1581_),
    .Y(_1617_)
);

NAND3X1 _8003_ (
    .A(1'h1),
    .B(_1057__bF$buf1),
    .C(_1030__bF$buf1),
    .Y(_1618_)
);

AOI21X1 _8004_ (
    .A(_1580_),
    .B(_1618_),
    .C(_1119__bF$buf5),
    .Y(_1619_)
);

NOR2X1 _8005_ (
    .A(_1619_),
    .B(_1617_),
    .Y(_1620_)
);

NAND2X1 _8006_ (
    .A(\genblk1[1].u_ce.Ain12b [4]),
    .B(_1620_),
    .Y(_1621_)
);

INVX1 _8007_ (
    .A(\genblk1[1].u_ce.Ain12b [4]),
    .Y(_1622_)
);

OAI21X1 _8008_ (
    .A(_1619_),
    .B(_1617_),
    .C(_1622_),
    .Y(_1623_)
);

NAND2X1 _8009_ (
    .A(_1623_),
    .B(_1621_),
    .Y(_1624_)
);

AOI21X1 _8010_ (
    .A(_1602_),
    .B(_1610_),
    .C(_1609_),
    .Y(_1625_)
);

AND2X2 _8011_ (
    .A(_1625_),
    .B(_1624_),
    .Y(_1626_)
);

OAI21X1 _8012_ (
    .A(_1624_),
    .B(_1625_),
    .C(\genblk1[1].u_ce.Vld_bF$buf3 ),
    .Y(_1627_)
);

OAI22X1 _8013_ (
    .A(_963_),
    .B(\genblk1[1].u_ce.Vld_bF$buf2 ),
    .C(_1627_),
    .D(_1626_),
    .Y(_896_)
);

NAND2X1 _8014_ (
    .A(\genblk1[1].u_ce.Acalc [5]),
    .B(_1024__bF$buf4),
    .Y(_1628_)
);

OAI21X1 _8015_ (
    .A(_1624_),
    .B(_1625_),
    .C(_1621_),
    .Y(_1629_)
);

OAI21X1 _8016_ (
    .A(1'h1),
    .B(1'h0),
    .C(_1058_),
    .Y(_1630_)
);

NAND2X1 _8017_ (
    .A(_1119__bF$buf4),
    .B(_1630_),
    .Y(_1631_)
);

INVX1 _8018_ (
    .A(_1631_),
    .Y(_1632_)
);

NOR2X1 _8019_ (
    .A(_1119__bF$buf3),
    .B(_1630_),
    .Y(_1633_)
);

NOR2X1 _8020_ (
    .A(_1633_),
    .B(_1632_),
    .Y(_1634_)
);

NAND2X1 _8021_ (
    .A(\genblk1[1].u_ce.Ain12b [5]),
    .B(_1634_),
    .Y(_1635_)
);

INVX1 _8022_ (
    .A(\genblk1[1].u_ce.Ain12b [5]),
    .Y(_1636_)
);

OAI21X1 _8023_ (
    .A(_1633_),
    .B(_1632_),
    .C(_1636_),
    .Y(_1637_)
);

NAND2X1 _8024_ (
    .A(_1637_),
    .B(_1635_),
    .Y(_1638_)
);

INVX1 _8025_ (
    .A(_1638_),
    .Y(_1639_)
);

NOR2X1 _8026_ (
    .A(_1639_),
    .B(_1629_),
    .Y(_1640_)
);

NAND2X1 _8027_ (
    .A(_1639_),
    .B(_1629_),
    .Y(_1641_)
);

NAND2X1 _8028_ (
    .A(\genblk1[1].u_ce.Vld_bF$buf1 ),
    .B(_1641_),
    .Y(_1642_)
);

OAI21X1 _8029_ (
    .A(_1640_),
    .B(_1642_),
    .C(_1628_),
    .Y(_897_)
);

NAND2X1 _8030_ (
    .A(\genblk1[1].u_ce.Acalc [6]),
    .B(_1024__bF$buf3),
    .Y(_1643_)
);

INVX1 _8031_ (
    .A(_1625_),
    .Y(_1644_)
);

NOR2X1 _8032_ (
    .A(_1624_),
    .B(_1638_),
    .Y(_1645_)
);

OAI21X1 _8033_ (
    .A(_1621_),
    .B(_1638_),
    .C(_1635_),
    .Y(_1646_)
);

AOI21X1 _8034_ (
    .A(_1644_),
    .B(_1645_),
    .C(_1646_),
    .Y(_1647_)
);

OAI21X1 _8035_ (
    .A(1'h0),
    .B(_1573_),
    .C(_1028_),
    .Y(_1648_)
);

NOR2X1 _8036_ (
    .A(_1119__bF$buf2),
    .B(_1648_),
    .Y(_1649_)
);

NAND2X1 _8037_ (
    .A(_1119__bF$buf1),
    .B(_1648_),
    .Y(_1650_)
);

INVX1 _8038_ (
    .A(_1650_),
    .Y(_1651_)
);

NOR2X1 _8039_ (
    .A(_1649_),
    .B(_1651_),
    .Y(_1652_)
);

NAND2X1 _8040_ (
    .A(\genblk1[1].u_ce.Ain12b [6]),
    .B(_1652_),
    .Y(_1653_)
);

OR2X2 _8041_ (
    .A(_1652_),
    .B(\genblk1[1].u_ce.Ain12b [6]),
    .Y(_1654_)
);

AND2X2 _8042_ (
    .A(_1654_),
    .B(_1653_),
    .Y(_1655_)
);

INVX1 _8043_ (
    .A(_1655_),
    .Y(_1656_)
);

AND2X2 _8044_ (
    .A(_1647_),
    .B(_1656_),
    .Y(_1657_)
);

OAI21X1 _8045_ (
    .A(_1656_),
    .B(_1647_),
    .C(\genblk1[1].u_ce.Vld_bF$buf0 ),
    .Y(_1658_)
);

OAI21X1 _8046_ (
    .A(_1658_),
    .B(_1657_),
    .C(_1643_),
    .Y(_898_)
);

OAI21X1 _8047_ (
    .A(_1656_),
    .B(_1647_),
    .C(_1653_),
    .Y(_1659_)
);

OAI21X1 _8048_ (
    .A(1'h0),
    .B(1'h1),
    .C(\genblk1[1].u_ce.Ain12b_11_bF$buf0 ),
    .Y(_1660_)
);

NAND2X1 _8049_ (
    .A(_1660_),
    .B(_1120_),
    .Y(_1661_)
);

INVX1 _8050_ (
    .A(_1661_),
    .Y(_1662_)
);

NAND2X1 _8051_ (
    .A(\genblk1[1].u_ce.Ain12b [7]),
    .B(_1662_),
    .Y(_1663_)
);

INVX1 _8052_ (
    .A(_1663_),
    .Y(_1664_)
);

NOR2X1 _8053_ (
    .A(\genblk1[1].u_ce.Ain12b [7]),
    .B(_1662_),
    .Y(_1665_)
);

NOR2X1 _8054_ (
    .A(_1665_),
    .B(_1664_),
    .Y(_1666_)
);

INVX1 _8055_ (
    .A(_1666_),
    .Y(_1667_)
);

OR2X2 _8056_ (
    .A(_1659_),
    .B(_1667_),
    .Y(_1668_)
);

AOI21X1 _8057_ (
    .A(_1659_),
    .B(_1667_),
    .C(_1024__bF$buf2),
    .Y(_1669_)
);

AOI22X1 _8058_ (
    .A(_977_),
    .B(_1024__bF$buf1),
    .C(_1668_),
    .D(_1669_),
    .Y(_899_)
);

NAND2X1 _8059_ (
    .A(\genblk1[1].u_ce.Acalc [8]),
    .B(_1024__bF$buf0),
    .Y(_1670_)
);

OAI21X1 _8060_ (
    .A(_1665_),
    .B(_1653_),
    .C(_1663_),
    .Y(_1671_)
);

NAND2X1 _8061_ (
    .A(_1666_),
    .B(_1655_),
    .Y(_1672_)
);

INVX1 _8062_ (
    .A(_1672_),
    .Y(_1673_)
);

AOI21X1 _8063_ (
    .A(_1673_),
    .B(_1646_),
    .C(_1671_),
    .Y(_1674_)
);

NAND2X1 _8064_ (
    .A(_1645_),
    .B(_1673_),
    .Y(_1675_)
);

OAI21X1 _8065_ (
    .A(_1675_),
    .B(_1625_),
    .C(_1674_),
    .Y(_1676_)
);

INVX1 _8066_ (
    .A(\genblk1[1].u_ce.Ain12b [8]),
    .Y(_1677_)
);

NAND2X1 _8067_ (
    .A(_1119__bF$buf0),
    .B(_1027_),
    .Y(_1678_)
);

NAND2X1 _8068_ (
    .A(_1607_),
    .B(_1678_),
    .Y(_1679_)
);

OR2X2 _8069_ (
    .A(_1679_),
    .B(_1677_),
    .Y(_1680_)
);

NAND2X1 _8070_ (
    .A(_1677_),
    .B(_1679_),
    .Y(_1681_)
);

AND2X2 _8071_ (
    .A(_1680_),
    .B(_1681_),
    .Y(_1682_)
);

NOR2X1 _8072_ (
    .A(_1682_),
    .B(_1676_),
    .Y(_1683_)
);

NAND2X1 _8073_ (
    .A(_1682_),
    .B(_1676_),
    .Y(_1684_)
);

NAND2X1 _8074_ (
    .A(\genblk1[1].u_ce.Vld_bF$buf4 ),
    .B(_1684_),
    .Y(_1685_)
);

OAI21X1 _8075_ (
    .A(_1683_),
    .B(_1685_),
    .C(_1670_),
    .Y(_900_)
);

NAND2X1 _8076_ (
    .A(\genblk1[1].u_ce.Acalc [9]),
    .B(_1024__bF$buf4),
    .Y(_1686_)
);

OAI21X1 _8077_ (
    .A(_1677_),
    .B(_1679_),
    .C(_1684_),
    .Y(_1687_)
);

INVX1 _8078_ (
    .A(\genblk1[1].u_ce.Ain12b [9]),
    .Y(_1688_)
);

NAND2X1 _8079_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf4 ),
    .B(_1688_),
    .Y(_1689_)
);

NOR2X1 _8080_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1688_),
    .Y(_1690_)
);

INVX1 _8081_ (
    .A(_1690_),
    .Y(_1691_)
);

NAND2X1 _8082_ (
    .A(_1689_),
    .B(_1691_),
    .Y(_1692_)
);

INVX1 _8083_ (
    .A(_1692_),
    .Y(_1693_)
);

NOR2X1 _8084_ (
    .A(_1693_),
    .B(_1687_),
    .Y(_1694_)
);

NAND2X1 _8085_ (
    .A(_1693_),
    .B(_1687_),
    .Y(_1695_)
);

NAND2X1 _8086_ (
    .A(\genblk1[1].u_ce.Vld_bF$buf3 ),
    .B(_1695_),
    .Y(_1696_)
);

OAI21X1 _8087_ (
    .A(_1694_),
    .B(_1696_),
    .C(_1686_),
    .Y(_901_)
);

AOI21X1 _8088_ (
    .A(_1687_),
    .B(_1689_),
    .C(_1690_),
    .Y(_1697_)
);

INVX1 _8089_ (
    .A(\genblk1[1].u_ce.Ain12b [10]),
    .Y(_1698_)
);

NAND2X1 _8090_ (
    .A(\genblk1[1].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1698_),
    .Y(_1699_)
);

NAND2X1 _8091_ (
    .A(\genblk1[1].u_ce.Ain12b [10]),
    .B(_1119__bF$buf5),
    .Y(_1700_)
);

NAND2X1 _8092_ (
    .A(_1699_),
    .B(_1700_),
    .Y(_1701_)
);

AND2X2 _8093_ (
    .A(_1697_),
    .B(_1701_),
    .Y(_1702_)
);

OAI21X1 _8094_ (
    .A(_1701_),
    .B(_1697_),
    .C(\genblk1[1].u_ce.Vld_bF$buf2 ),
    .Y(_1703_)
);

OAI22X1 _8095_ (
    .A(_959_),
    .B(\genblk1[1].u_ce.Vld_bF$buf1 ),
    .C(_1703_),
    .D(_1702_),
    .Y(_902_)
);

NAND2X1 _8096_ (
    .A(\genblk1[1].u_ce.Acalc [11]),
    .B(_1024__bF$buf3),
    .Y(_1704_)
);

OAI21X1 _8097_ (
    .A(_1701_),
    .B(_1697_),
    .C(_1700_),
    .Y(_1705_)
);

OAI21X1 _8098_ (
    .A(_1024__bF$buf2),
    .B(_1705_),
    .C(_1704_),
    .Y(_903_)
);

INVX1 _8099_ (
    .A(_958_),
    .Y(_1706_)
);

NAND3X1 _8100_ (
    .A(_1011_),
    .B(\genblk1[1].u_ce.LoadCtl [5]),
    .C(_969_),
    .Y(_1707_)
);

NOR2X1 _8101_ (
    .A(_1706_),
    .B(_1707_),
    .Y(_1708_)
);

NAND2X1 _8102_ (
    .A(\genblk1[0].u_ce.X_ [0]),
    .B(_1708_),
    .Y(_1709_)
);

OAI21X1 _8103_ (
    .A(_1153_),
    .B(_1708_),
    .C(_1709_),
    .Y(_904_)
);

NAND2X1 _8104_ (
    .A(\genblk1[0].u_ce.X_ [1]),
    .B(_1708_),
    .Y(_1710_)
);

OAI21X1 _8105_ (
    .A(_1178_),
    .B(_1708_),
    .C(_1710_),
    .Y(_905_)
);

INVX1 _8106_ (
    .A(\genblk1[0].u_ce.X_ [0]),
    .Y(_1711_)
);

NAND3X1 _8107_ (
    .A(\genblk1[1].u_ce.LoadCtl [4]),
    .B(_958_),
    .C(_969_),
    .Y(_1712_)
);

NAND2X1 _8108_ (
    .A(\genblk1[1].u_ce.Xin12b [8]),
    .B(_1712_),
    .Y(_1713_)
);

OAI21X1 _8109_ (
    .A(_1711_),
    .B(_1712_),
    .C(_1713_),
    .Y(_906_)
);

INVX1 _8110_ (
    .A(\genblk1[0].u_ce.X_ [1]),
    .Y(_1714_)
);

NAND2X1 _8111_ (
    .A(\genblk1[1].u_ce.Xin12b [9]),
    .B(_1712_),
    .Y(_1715_)
);

OAI21X1 _8112_ (
    .A(_1714_),
    .B(_1712_),
    .C(_1715_),
    .Y(_907_)
);

NAND2X1 _8113_ (
    .A(_969_),
    .B(_965_),
    .Y(_1716_)
);

OAI21X1 _8114_ (
    .A(_970_),
    .B(_978_),
    .C(\genblk1[1].u_ce.Xin12b [6]),
    .Y(_1717_)
);

OAI21X1 _8115_ (
    .A(_1711_),
    .B(_1716_),
    .C(_1717_),
    .Y(_908_)
);

OAI21X1 _8116_ (
    .A(_970_),
    .B(_978_),
    .C(\genblk1[1].u_ce.Xin12b [7]),
    .Y(_1718_)
);

OAI21X1 _8117_ (
    .A(_1714_),
    .B(_1716_),
    .C(_1718_),
    .Y(_909_)
);

NOR2X1 _8118_ (
    .A(_962_),
    .B(_970_),
    .Y(_1719_)
);

NAND2X1 _8119_ (
    .A(\genblk1[0].u_ce.X_ [0]),
    .B(_1719_),
    .Y(_1720_)
);

OAI21X1 _8120_ (
    .A(_1063_),
    .B(_1719_),
    .C(_1720_),
    .Y(_910_)
);

NAND2X1 _8121_ (
    .A(\genblk1[0].u_ce.X_ [1]),
    .B(_1719_),
    .Y(_1721_)
);

OAI21X1 _8122_ (
    .A(_1071_),
    .B(_1719_),
    .C(_1721_),
    .Y(_911_)
);

OAI21X1 _8123_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_971_),
    .C(\genblk1[1].u_ce.Xin1 [0]),
    .Y(_1722_)
);

OAI21X1 _8124_ (
    .A(_1711_),
    .B(_1000_),
    .C(_1722_),
    .Y(_912_)
);

OAI21X1 _8125_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_971_),
    .C(\genblk1[1].u_ce.Xin1 [1]),
    .Y(_1723_)
);

OAI21X1 _8126_ (
    .A(_1714_),
    .B(_1000_),
    .C(_1723_),
    .Y(_913_)
);

NAND2X1 _8127_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[0].u_ce.X_ [0]),
    .Y(_1724_)
);

OAI21X1 _8128_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_1086_),
    .C(_1724_),
    .Y(_914_)
);

NAND2X1 _8129_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[0].u_ce.X_ [1]),
    .Y(_1725_)
);

OAI21X1 _8130_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_1066_),
    .C(_1725_),
    .Y(_915_)
);

NAND2X1 _8131_ (
    .A(\genblk1[0].u_ce.Y_ [0]),
    .B(_1708_),
    .Y(_1726_)
);

OAI21X1 _8132_ (
    .A(_1286_),
    .B(_1708_),
    .C(_1726_),
    .Y(_916_)
);

NAND2X1 _8133_ (
    .A(\genblk1[0].u_ce.Y_ [1]),
    .B(_1708_),
    .Y(_1727_)
);

OAI21X1 _8134_ (
    .A(_1310_),
    .B(_1708_),
    .C(_1727_),
    .Y(_917_)
);

INVX1 _8135_ (
    .A(\genblk1[0].u_ce.Y_ [0]),
    .Y(_1728_)
);

NAND2X1 _8136_ (
    .A(\genblk1[1].u_ce.Yin12b [8]),
    .B(_1712_),
    .Y(_1729_)
);

OAI21X1 _8137_ (
    .A(_1728_),
    .B(_1712_),
    .C(_1729_),
    .Y(_918_)
);

INVX1 _8138_ (
    .A(\genblk1[0].u_ce.Y_ [1]),
    .Y(_1730_)
);

NAND2X1 _8139_ (
    .A(\genblk1[1].u_ce.Yin12b [9]),
    .B(_1712_),
    .Y(_1731_)
);

OAI21X1 _8140_ (
    .A(_1730_),
    .B(_1712_),
    .C(_1731_),
    .Y(_919_)
);

OAI21X1 _8141_ (
    .A(_970_),
    .B(_978_),
    .C(\genblk1[1].u_ce.Yin12b [6]),
    .Y(_938_)
);

OAI21X1 _8142_ (
    .A(_1728_),
    .B(_1716_),
    .C(_938_),
    .Y(_920_)
);

OAI21X1 _8143_ (
    .A(_970_),
    .B(_978_),
    .C(\genblk1[1].u_ce.Yin12b [7]),
    .Y(_939_)
);

OAI21X1 _8144_ (
    .A(_1730_),
    .B(_1716_),
    .C(_939_),
    .Y(_921_)
);

NAND2X1 _8145_ (
    .A(\genblk1[0].u_ce.Y_ [0]),
    .B(_1719_),
    .Y(_940_)
);

OAI21X1 _8146_ (
    .A(_1151_),
    .B(_1719_),
    .C(_940_),
    .Y(_922_)
);

NAND2X1 _8147_ (
    .A(\genblk1[0].u_ce.Y_ [1]),
    .B(_1719_),
    .Y(_941_)
);

OAI21X1 _8148_ (
    .A(_1176_),
    .B(_1719_),
    .C(_941_),
    .Y(_923_)
);

OAI21X1 _8149_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_971_),
    .C(\genblk1[1].u_ce.Yin1 [0]),
    .Y(_942_)
);

OAI21X1 _8150_ (
    .A(_1728_),
    .B(_1000_),
    .C(_942_),
    .Y(_924_)
);

OAI21X1 _8151_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_971_),
    .C(\genblk1[1].u_ce.Yin1 [1]),
    .Y(_943_)
);

OAI21X1 _8152_ (
    .A(_1730_),
    .B(_1000_),
    .C(_943_),
    .Y(_925_)
);

NAND2X1 _8153_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[0].u_ce.Y_ [0]),
    .Y(_944_)
);

OAI21X1 _8154_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_1323_),
    .C(_944_),
    .Y(_926_)
);

NAND2X1 _8155_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[0].u_ce.Y_ [1]),
    .Y(_945_)
);

OAI21X1 _8156_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_1108_),
    .C(_945_),
    .Y(_927_)
);

NAND2X1 _8157_ (
    .A(\a[1] [0]),
    .B(_1708_),
    .Y(_946_)
);

OAI21X1 _8158_ (
    .A(_1698_),
    .B(_1708_),
    .C(_946_),
    .Y(_928_)
);

NAND2X1 _8159_ (
    .A(\a[1] [1]),
    .B(_1708_),
    .Y(_947_)
);

OAI21X1 _8160_ (
    .A(_1119__bF$buf4),
    .B(_1708_),
    .C(_947_),
    .Y(_929_)
);

INVX1 _8161_ (
    .A(\a[1] [0]),
    .Y(_948_)
);

NAND2X1 _8162_ (
    .A(\genblk1[1].u_ce.Ain12b [8]),
    .B(_1712_),
    .Y(_949_)
);

OAI21X1 _8163_ (
    .A(_948_),
    .B(_1712_),
    .C(_949_),
    .Y(_930_)
);

INVX1 _8164_ (
    .A(\a[1] [1]),
    .Y(_950_)
);

NAND2X1 _8165_ (
    .A(\genblk1[1].u_ce.Ain12b [9]),
    .B(_1712_),
    .Y(_951_)
);

OAI21X1 _8166_ (
    .A(_950_),
    .B(_1712_),
    .C(_951_),
    .Y(_931_)
);

OAI21X1 _8167_ (
    .A(_970_),
    .B(_978_),
    .C(\genblk1[1].u_ce.Ain12b [6]),
    .Y(_952_)
);

OAI21X1 _8168_ (
    .A(_948_),
    .B(_1716_),
    .C(_952_),
    .Y(_932_)
);

OAI21X1 _8169_ (
    .A(_970_),
    .B(_978_),
    .C(\genblk1[1].u_ce.Ain12b [7]),
    .Y(_953_)
);

OAI21X1 _8170_ (
    .A(_950_),
    .B(_1716_),
    .C(_953_),
    .Y(_933_)
);

NAND2X1 _8171_ (
    .A(\a[1] [0]),
    .B(_1719_),
    .Y(_954_)
);

OAI21X1 _8172_ (
    .A(_1622_),
    .B(_1719_),
    .C(_954_),
    .Y(_934_)
);

NAND2X1 _8173_ (
    .A(\a[1] [1]),
    .B(_1719_),
    .Y(_955_)
);

OAI21X1 _8174_ (
    .A(_1636_),
    .B(_1719_),
    .C(_955_),
    .Y(_935_)
);

OAI21X1 _8175_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_971_),
    .C(\genblk1[1].u_ce.Ain1 [0]),
    .Y(_956_)
);

OAI21X1 _8176_ (
    .A(_948_),
    .B(_1000_),
    .C(_956_),
    .Y(_936_)
);

OAI21X1 _8177_ (
    .A(\genblk1[1].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_971_),
    .C(\genblk1[1].u_ce.Ain1 [1]),
    .Y(_957_)
);

OAI21X1 _8178_ (
    .A(_950_),
    .B(_1000_),
    .C(_957_),
    .Y(_937_)
);

DFFPOSX1 _8179_ (
    .CLK(clk_bF$buf29),
    .D(_866_),
    .Q(\genblk1[1].u_ce.Ain0 [0])
);

DFFPOSX1 _8180_ (
    .CLK(clk_bF$buf28),
    .D(_867_),
    .Q(\genblk1[1].u_ce.Ain0 [1])
);

DFFPOSX1 _8181_ (
    .CLK(clk_bF$buf27),
    .D(_868_),
    .Q(\genblk1[1].u_ce.Ycalc [2])
);

DFFPOSX1 _8182_ (
    .CLK(clk_bF$buf26),
    .D(_869_),
    .Q(\genblk1[1].u_ce.Ycalc [3])
);

DFFPOSX1 _8183_ (
    .CLK(clk_bF$buf25),
    .D(_870_),
    .Q(\genblk1[1].u_ce.Ycalc [4])
);

DFFPOSX1 _8184_ (
    .CLK(clk_bF$buf24),
    .D(_871_),
    .Q(\genblk1[1].u_ce.Ycalc [5])
);

DFFPOSX1 _8185_ (
    .CLK(clk_bF$buf23),
    .D(_872_),
    .Q(\genblk1[1].u_ce.Ycalc [6])
);

DFFPOSX1 _8186_ (
    .CLK(clk_bF$buf22),
    .D(_873_),
    .Q(\genblk1[1].u_ce.Ycalc [7])
);

DFFPOSX1 _8187_ (
    .CLK(clk_bF$buf21),
    .D(_874_),
    .Q(\genblk1[1].u_ce.Ycalc [8])
);

DFFPOSX1 _8188_ (
    .CLK(clk_bF$buf20),
    .D(_875_),
    .Q(\genblk1[1].u_ce.Ycalc [9])
);

DFFPOSX1 _8189_ (
    .CLK(clk_bF$buf19),
    .D(_876_),
    .Q(\genblk1[1].u_ce.Ycalc [10])
);

DFFPOSX1 _8190_ (
    .CLK(clk_bF$buf18),
    .D(_877_),
    .Q(\genblk1[1].u_ce.Ycalc [11])
);

DFFPOSX1 _8191_ (
    .CLK(clk_bF$buf17),
    .D(_878_),
    .Q(\genblk1[1].u_ce.Ycalc [0])
);

DFFPOSX1 _8192_ (
    .CLK(clk_bF$buf16),
    .D(_879_),
    .Q(\genblk1[1].u_ce.Ycalc [1])
);

DFFPOSX1 _8193_ (
    .CLK(clk_bF$buf15),
    .D(_880_),
    .Q(\genblk1[1].u_ce.Xcalc [0])
);

DFFPOSX1 _8194_ (
    .CLK(clk_bF$buf14),
    .D(_881_),
    .Q(\genblk1[1].u_ce.Xcalc [1])
);

DFFPOSX1 _8195_ (
    .CLK(clk_bF$buf13),
    .D(_882_),
    .Q(\genblk1[1].u_ce.Xcalc [2])
);

DFFPOSX1 _8196_ (
    .CLK(clk_bF$buf12),
    .D(_883_),
    .Q(\genblk1[1].u_ce.Xcalc [3])
);

DFFPOSX1 _8197_ (
    .CLK(clk_bF$buf11),
    .D(_884_),
    .Q(\genblk1[1].u_ce.Xcalc [4])
);

DFFPOSX1 _8198_ (
    .CLK(clk_bF$buf10),
    .D(_885_),
    .Q(\genblk1[1].u_ce.Xcalc [5])
);

DFFPOSX1 _8199_ (
    .CLK(clk_bF$buf9),
    .D(_886_),
    .Q(\genblk1[1].u_ce.Xcalc [6])
);

DFFPOSX1 _8200_ (
    .CLK(clk_bF$buf8),
    .D(_887_),
    .Q(\genblk1[1].u_ce.Xcalc [7])
);

DFFPOSX1 _8201_ (
    .CLK(clk_bF$buf7),
    .D(_888_),
    .Q(\genblk1[1].u_ce.Xcalc [8])
);

DFFPOSX1 _8202_ (
    .CLK(clk_bF$buf6),
    .D(_889_),
    .Q(\genblk1[1].u_ce.Xcalc [9])
);

DFFPOSX1 _8203_ (
    .CLK(clk_bF$buf5),
    .D(_890_),
    .Q(\genblk1[1].u_ce.Xcalc [10])
);

DFFPOSX1 _8204_ (
    .CLK(clk_bF$buf4),
    .D(_891_),
    .Q(\genblk1[1].u_ce.Xcalc [11])
);

DFFPOSX1 _8205_ (
    .CLK(clk_bF$buf3),
    .D(_892_),
    .Q(\genblk1[1].u_ce.Acalc [0])
);

DFFPOSX1 _8206_ (
    .CLK(clk_bF$buf2),
    .D(_893_),
    .Q(\genblk1[1].u_ce.Acalc [1])
);

DFFPOSX1 _8207_ (
    .CLK(clk_bF$buf1),
    .D(_894_),
    .Q(\genblk1[1].u_ce.Acalc [2])
);

DFFPOSX1 _8208_ (
    .CLK(clk_bF$buf0),
    .D(_895_),
    .Q(\genblk1[1].u_ce.Acalc [3])
);

DFFPOSX1 _8209_ (
    .CLK(clk_bF$buf75),
    .D(_896_),
    .Q(\genblk1[1].u_ce.Acalc [4])
);

DFFPOSX1 _8210_ (
    .CLK(clk_bF$buf74),
    .D(_897_),
    .Q(\genblk1[1].u_ce.Acalc [5])
);

DFFPOSX1 _8211_ (
    .CLK(clk_bF$buf73),
    .D(_898_),
    .Q(\genblk1[1].u_ce.Acalc [6])
);

DFFPOSX1 _8212_ (
    .CLK(clk_bF$buf72),
    .D(_899_),
    .Q(\genblk1[1].u_ce.Acalc [7])
);

DFFPOSX1 _8213_ (
    .CLK(clk_bF$buf71),
    .D(_900_),
    .Q(\genblk1[1].u_ce.Acalc [8])
);

DFFPOSX1 _8214_ (
    .CLK(clk_bF$buf70),
    .D(_901_),
    .Q(\genblk1[1].u_ce.Acalc [9])
);

DFFPOSX1 _8215_ (
    .CLK(clk_bF$buf69),
    .D(_902_),
    .Q(\genblk1[1].u_ce.Acalc [10])
);

DFFPOSX1 _8216_ (
    .CLK(clk_bF$buf68),
    .D(_903_),
    .Q(\genblk1[1].u_ce.Acalc [11])
);

DFFPOSX1 _8217_ (
    .CLK(clk_bF$buf67),
    .D(_904_),
    .Q(\genblk1[1].u_ce.Xin12b [10])
);

DFFPOSX1 _8218_ (
    .CLK(clk_bF$buf66),
    .D(_905_),
    .Q(\genblk1[1].u_ce.Xin12b [11])
);

DFFPOSX1 _8219_ (
    .CLK(clk_bF$buf65),
    .D(_906_),
    .Q(\genblk1[1].u_ce.Xin12b [8])
);

DFFPOSX1 _8220_ (
    .CLK(clk_bF$buf64),
    .D(_907_),
    .Q(\genblk1[1].u_ce.Xin12b [9])
);

DFFPOSX1 _8221_ (
    .CLK(clk_bF$buf63),
    .D(_908_),
    .Q(\genblk1[1].u_ce.Xin12b [6])
);

DFFPOSX1 _8222_ (
    .CLK(clk_bF$buf62),
    .D(_909_),
    .Q(\genblk1[1].u_ce.Xin12b [7])
);

DFFPOSX1 _8223_ (
    .CLK(clk_bF$buf61),
    .D(_910_),
    .Q(\genblk1[1].u_ce.Xin12b [4])
);

DFFPOSX1 _8224_ (
    .CLK(clk_bF$buf60),
    .D(_911_),
    .Q(\genblk1[1].u_ce.Xin12b [5])
);

DFFPOSX1 _8225_ (
    .CLK(clk_bF$buf59),
    .D(_912_),
    .Q(\genblk1[1].u_ce.Xin1 [0])
);

DFFPOSX1 _8226_ (
    .CLK(clk_bF$buf58),
    .D(_913_),
    .Q(\genblk1[1].u_ce.Xin1 [1])
);

DFFPOSX1 _8227_ (
    .CLK(clk_bF$buf57),
    .D(_914_),
    .Q(\genblk1[1].u_ce.Xin0 [0])
);

DFFPOSX1 _8228_ (
    .CLK(clk_bF$buf56),
    .D(_915_),
    .Q(\genblk1[1].u_ce.Xin0 [1])
);

DFFPOSX1 _8229_ (
    .CLK(clk_bF$buf55),
    .D(_916_),
    .Q(\genblk1[1].u_ce.Yin12b [10])
);

DFFPOSX1 _8230_ (
    .CLK(clk_bF$buf54),
    .D(_917_),
    .Q(\genblk1[1].u_ce.Yin12b [11])
);

DFFPOSX1 _8231_ (
    .CLK(clk_bF$buf53),
    .D(_918_),
    .Q(\genblk1[1].u_ce.Yin12b [8])
);

DFFPOSX1 _8232_ (
    .CLK(clk_bF$buf52),
    .D(_919_),
    .Q(\genblk1[1].u_ce.Yin12b [9])
);

DFFPOSX1 _8233_ (
    .CLK(clk_bF$buf51),
    .D(_920_),
    .Q(\genblk1[1].u_ce.Yin12b [6])
);

DFFPOSX1 _8234_ (
    .CLK(clk_bF$buf50),
    .D(_921_),
    .Q(\genblk1[1].u_ce.Yin12b [7])
);

DFFPOSX1 _8235_ (
    .CLK(clk_bF$buf49),
    .D(_922_),
    .Q(\genblk1[1].u_ce.Yin12b [4])
);

DFFPOSX1 _8236_ (
    .CLK(clk_bF$buf48),
    .D(_923_),
    .Q(\genblk1[1].u_ce.Yin12b [5])
);

DFFPOSX1 _8237_ (
    .CLK(clk_bF$buf47),
    .D(_924_),
    .Q(\genblk1[1].u_ce.Yin1 [0])
);

DFFPOSX1 _8238_ (
    .CLK(clk_bF$buf46),
    .D(_925_),
    .Q(\genblk1[1].u_ce.Yin1 [1])
);

DFFPOSX1 _8239_ (
    .CLK(clk_bF$buf45),
    .D(_926_),
    .Q(\genblk1[1].u_ce.Yin0 [0])
);

DFFPOSX1 _8240_ (
    .CLK(clk_bF$buf44),
    .D(_927_),
    .Q(\genblk1[1].u_ce.Yin0 [1])
);

DFFPOSX1 _8241_ (
    .CLK(clk_bF$buf43),
    .D(_928_),
    .Q(\genblk1[1].u_ce.Ain12b [10])
);

DFFPOSX1 _8242_ (
    .CLK(clk_bF$buf42),
    .D(_929_),
    .Q(\genblk1[1].u_ce.Ain12b [11])
);

DFFPOSX1 _8243_ (
    .CLK(clk_bF$buf41),
    .D(_930_),
    .Q(\genblk1[1].u_ce.Ain12b [8])
);

DFFPOSX1 _8244_ (
    .CLK(clk_bF$buf40),
    .D(_931_),
    .Q(\genblk1[1].u_ce.Ain12b [9])
);

DFFPOSX1 _8245_ (
    .CLK(clk_bF$buf39),
    .D(_932_),
    .Q(\genblk1[1].u_ce.Ain12b [6])
);

DFFPOSX1 _8246_ (
    .CLK(clk_bF$buf38),
    .D(_933_),
    .Q(\genblk1[1].u_ce.Ain12b [7])
);

DFFPOSX1 _8247_ (
    .CLK(clk_bF$buf37),
    .D(_934_),
    .Q(\genblk1[1].u_ce.Ain12b [4])
);

DFFPOSX1 _8248_ (
    .CLK(clk_bF$buf36),
    .D(_935_),
    .Q(\genblk1[1].u_ce.Ain12b [5])
);

DFFPOSX1 _8249_ (
    .CLK(clk_bF$buf35),
    .D(_936_),
    .Q(\genblk1[1].u_ce.Ain1 [0])
);

DFFPOSX1 _8250_ (
    .CLK(clk_bF$buf34),
    .D(_937_),
    .Q(\genblk1[1].u_ce.Ain1 [1])
);

DFFPOSX1 _8251_ (
    .CLK(clk_bF$buf33),
    .D(\genblk1[0].u_ce.ISout ),
    .Q(\genblk1[1].u_ce.ISpipe [0])
);

DFFPOSX1 _8252_ (
    .CLK(clk_bF$buf32),
    .D(\genblk1[1].u_ce.ISpipe [0]),
    .Q(\genblk1[1].u_ce.ISpipe [1])
);

DFFPOSX1 _8253_ (
    .CLK(clk_bF$buf31),
    .D(\genblk1[1].u_ce.ISpipe [1]),
    .Q(\genblk1[1].u_ce.ISpipe [2])
);

DFFPOSX1 _8254_ (
    .CLK(clk_bF$buf30),
    .D(\genblk1[1].u_ce.ISpipe [2]),
    .Q(\genblk1[1].u_ce.ISpipe [3])
);

DFFPOSX1 _8255_ (
    .CLK(clk_bF$buf29),
    .D(\genblk1[1].u_ce.ISpipe [3]),
    .Q(\genblk1[1].u_ce.ISpipe [4])
);

DFFPOSX1 _8256_ (
    .CLK(clk_bF$buf28),
    .D(\genblk1[1].u_ce.ISpipe [4]),
    .Q(\genblk1[1].u_ce.ISpipe [5])
);

DFFPOSX1 _8257_ (
    .CLK(clk_bF$buf27),
    .D(\genblk1[1].u_ce.ISpipe [5]),
    .Q(\genblk1[1].u_ce.ISout )
);

DFFPOSX1 _8258_ (
    .CLK(clk_bF$buf26),
    .D(\genblk1[0].u_ce.Vld_bF$buf0 ),
    .Q(\genblk1[1].u_ce.LoadCtl [0])
);

DFFPOSX1 _8259_ (
    .CLK(clk_bF$buf25),
    .D(\genblk1[1].u_ce.LoadCtl_0_bF$buf3 ),
    .Q(\genblk1[1].u_ce.LoadCtl [1])
);

DFFPOSX1 _8260_ (
    .CLK(clk_bF$buf24),
    .D(\genblk1[1].u_ce.LoadCtl [1]),
    .Q(\genblk1[1].u_ce.LoadCtl [2])
);

DFFPOSX1 _8261_ (
    .CLK(clk_bF$buf23),
    .D(\genblk1[1].u_ce.LoadCtl [2]),
    .Q(\genblk1[1].u_ce.LoadCtl [3])
);

DFFPOSX1 _8262_ (
    .CLK(clk_bF$buf22),
    .D(\genblk1[1].u_ce.LoadCtl [3]),
    .Q(\genblk1[1].u_ce.LoadCtl [4])
);

DFFPOSX1 _8263_ (
    .CLK(clk_bF$buf21),
    .D(\genblk1[1].u_ce.LoadCtl [4]),
    .Q(\genblk1[1].u_ce.LoadCtl [5])
);

DFFPOSX1 _8264_ (
    .CLK(clk_bF$buf20),
    .D(\genblk1[1].u_ce.LoadCtl [5]),
    .Q(\genblk1[1].u_ce.Vld )
);

NOR2X1 _8265_ (
    .A(\genblk1[2].u_ce.LoadCtl [3]),
    .B(\genblk1[2].u_ce.LoadCtl [2]),
    .Y(_1824_)
);

INVX1 _8266_ (
    .A(\genblk1[2].u_ce.Acalc [10]),
    .Y(_1825_)
);

NAND2X1 _8267_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(\genblk1[2].u_ce.Acalc [8]),
    .Y(_1826_)
);

OAI21X1 _8268_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(_1825_),
    .C(_1826_),
    .Y(_1827_)
);

INVX2 _8269_ (
    .A(\genblk1[2].u_ce.LoadCtl [2]),
    .Y(_1828_)
);

INVX1 _8270_ (
    .A(\genblk1[2].u_ce.Acalc [4]),
    .Y(_1829_)
);

INVX1 _8271_ (
    .A(\genblk1[2].u_ce.LoadCtl [3]),
    .Y(_1830_)
);

NOR2X1 _8272_ (
    .A(\genblk1[2].u_ce.LoadCtl [2]),
    .B(_1830_),
    .Y(_1831_)
);

NAND2X1 _8273_ (
    .A(\genblk1[2].u_ce.Acalc [6]),
    .B(_1831_),
    .Y(_1832_)
);

OAI21X1 _8274_ (
    .A(_1828_),
    .B(_1829_),
    .C(_1832_),
    .Y(_1833_)
);

AOI21X1 _8275_ (
    .A(_1824_),
    .B(_1827_),
    .C(_1833_),
    .Y(_1834_)
);

NOR2X1 _8276_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[2].u_ce.LoadCtl [1]),
    .Y(_1835_)
);

INVX4 _8277_ (
    .A(_1835_),
    .Y(_1836_)
);

INVX2 _8278_ (
    .A(\genblk1[2].u_ce.LoadCtl [1]),
    .Y(_1837_)
);

NOR2X1 _8279_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_1837_),
    .Y(_1838_)
);

AOI22X1 _8280_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[2].u_ce.Acalc [0]),
    .C(_1838_),
    .D(\genblk1[2].u_ce.Acalc [2]),
    .Y(_1839_)
);

OAI21X1 _8281_ (
    .A(_1836_),
    .B(_1834_),
    .C(_1839_),
    .Y(\a[3] [0])
);

INVX1 _8282_ (
    .A(\genblk1[2].u_ce.Acalc [11]),
    .Y(_1840_)
);

NAND2X1 _8283_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(\genblk1[2].u_ce.Acalc [9]),
    .Y(_1841_)
);

OAI21X1 _8284_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(_1840_),
    .C(_1841_),
    .Y(_1842_)
);

INVX1 _8285_ (
    .A(\genblk1[2].u_ce.Acalc [7]),
    .Y(_1843_)
);

INVX4 _8286_ (
    .A(_1831_),
    .Y(_1844_)
);

NAND2X1 _8287_ (
    .A(\genblk1[2].u_ce.LoadCtl [2]),
    .B(\genblk1[2].u_ce.Acalc [5]),
    .Y(_1845_)
);

OAI21X1 _8288_ (
    .A(_1843_),
    .B(_1844_),
    .C(_1845_),
    .Y(_1846_)
);

AOI21X1 _8289_ (
    .A(_1824_),
    .B(_1842_),
    .C(_1846_),
    .Y(_1847_)
);

AOI22X1 _8290_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[2].u_ce.Acalc [1]),
    .C(_1838_),
    .D(\genblk1[2].u_ce.Acalc [3]),
    .Y(_1848_)
);

OAI21X1 _8291_ (
    .A(_1836_),
    .B(_1847_),
    .C(_1848_),
    .Y(\a[3] [1])
);

INVX1 _8292_ (
    .A(\genblk1[2].u_ce.Ycalc [10]),
    .Y(_1849_)
);

NAND2X1 _8293_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(\genblk1[2].u_ce.Ycalc [8]),
    .Y(_1850_)
);

OAI21X1 _8294_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(_1849_),
    .C(_1850_),
    .Y(_1851_)
);

INVX1 _8295_ (
    .A(\genblk1[2].u_ce.Ycalc [6]),
    .Y(_1852_)
);

INVX1 _8296_ (
    .A(\genblk1[2].u_ce.Ycalc [4]),
    .Y(_1853_)
);

OAI22X1 _8297_ (
    .A(_1828_),
    .B(_1853_),
    .C(_1852_),
    .D(_1844_),
    .Y(_1854_)
);

AOI21X1 _8298_ (
    .A(_1824_),
    .B(_1851_),
    .C(_1854_),
    .Y(_1855_)
);

AOI22X1 _8299_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[2].u_ce.Ycalc [0]),
    .C(_1838_),
    .D(\genblk1[2].u_ce.Ycalc [2]),
    .Y(_1856_)
);

OAI21X1 _8300_ (
    .A(_1836_),
    .B(_1855_),
    .C(_1856_),
    .Y(\genblk1[2].u_ce.Y_ [0])
);

INVX1 _8301_ (
    .A(\genblk1[2].u_ce.Ycalc [11]),
    .Y(_1857_)
);

NAND2X1 _8302_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(\genblk1[2].u_ce.Ycalc [9]),
    .Y(_1858_)
);

OAI21X1 _8303_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(_1857_),
    .C(_1858_),
    .Y(_1859_)
);

INVX1 _8304_ (
    .A(\genblk1[2].u_ce.Ycalc [7]),
    .Y(_1860_)
);

INVX1 _8305_ (
    .A(\genblk1[2].u_ce.Ycalc [5]),
    .Y(_1861_)
);

OAI22X1 _8306_ (
    .A(_1828_),
    .B(_1861_),
    .C(_1860_),
    .D(_1844_),
    .Y(_1862_)
);

AOI21X1 _8307_ (
    .A(_1824_),
    .B(_1859_),
    .C(_1862_),
    .Y(_1863_)
);

AOI22X1 _8308_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[2].u_ce.Ycalc [1]),
    .C(_1838_),
    .D(\genblk1[2].u_ce.Ycalc [3]),
    .Y(_1864_)
);

OAI21X1 _8309_ (
    .A(_1836_),
    .B(_1863_),
    .C(_1864_),
    .Y(\genblk1[2].u_ce.Y_ [1])
);

INVX1 _8310_ (
    .A(\genblk1[2].u_ce.Xcalc [2]),
    .Y(_1865_)
);

INVX2 _8311_ (
    .A(_1838_),
    .Y(_1866_)
);

INVX1 _8312_ (
    .A(\genblk1[2].u_ce.Xcalc [4]),
    .Y(_1867_)
);

INVX1 _8313_ (
    .A(\genblk1[2].u_ce.Xcalc [6]),
    .Y(_1868_)
);

NOR2X1 _8314_ (
    .A(_1830_),
    .B(_1868_),
    .Y(_1869_)
);

INVX1 _8315_ (
    .A(\genblk1[2].u_ce.Xcalc [8]),
    .Y(_1870_)
);

NAND2X1 _8316_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(_1870_),
    .Y(_1871_)
);

OAI21X1 _8317_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(\genblk1[2].u_ce.Xcalc [10]),
    .C(_1871_),
    .Y(_1872_)
);

NOR2X1 _8318_ (
    .A(\genblk1[2].u_ce.LoadCtl [3]),
    .B(_1872_),
    .Y(_1873_)
);

OAI21X1 _8319_ (
    .A(_1869_),
    .B(_1873_),
    .C(_1828_),
    .Y(_1874_)
);

OAI21X1 _8320_ (
    .A(_1828_),
    .B(_1867_),
    .C(_1874_),
    .Y(_1875_)
);

AOI22X1 _8321_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[2].u_ce.Xcalc [0]),
    .C(_1875_),
    .D(_1835_),
    .Y(_1876_)
);

OAI21X1 _8322_ (
    .A(_1865_),
    .B(_1866_),
    .C(_1876_),
    .Y(\genblk1[2].u_ce.X_ [0])
);

INVX1 _8323_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .Y(_1877_)
);

INVX1 _8324_ (
    .A(\genblk1[2].u_ce.Xcalc [9]),
    .Y(_1878_)
);

NAND2X1 _8325_ (
    .A(\genblk1[2].u_ce.Xcalc [11]),
    .B(_1877_),
    .Y(_1879_)
);

OAI21X1 _8326_ (
    .A(_1877_),
    .B(_1878_),
    .C(_1879_),
    .Y(_1880_)
);

INVX1 _8327_ (
    .A(\genblk1[2].u_ce.Xcalc [7]),
    .Y(_1881_)
);

INVX1 _8328_ (
    .A(\genblk1[2].u_ce.Xcalc [5]),
    .Y(_1882_)
);

OAI22X1 _8329_ (
    .A(_1828_),
    .B(_1882_),
    .C(_1881_),
    .D(_1844_),
    .Y(_1883_)
);

AOI21X1 _8330_ (
    .A(_1824_),
    .B(_1880_),
    .C(_1883_),
    .Y(_1884_)
);

AOI22X1 _8331_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[2].u_ce.Xcalc [1]),
    .C(_1838_),
    .D(\genblk1[2].u_ce.Xcalc [3]),
    .Y(_1885_)
);

OAI21X1 _8332_ (
    .A(_1836_),
    .B(_1884_),
    .C(_1885_),
    .Y(\genblk1[2].u_ce.X_ [1])
);

INVX1 _8333_ (
    .A(\genblk1[2].u_ce.Ain0 [0]),
    .Y(_1886_)
);

NAND2X1 _8334_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\a[2] [0]),
    .Y(_1887_)
);

OAI21X1 _8335_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_1886_),
    .C(_1887_),
    .Y(_1732_)
);

INVX1 _8336_ (
    .A(\genblk1[2].u_ce.Ain0 [1]),
    .Y(_1888_)
);

NAND2X1 _8337_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\a[2] [1]),
    .Y(_1889_)
);

OAI21X1 _8338_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_1888_),
    .C(_1889_),
    .Y(_1733_)
);

INVX8 _8339_ (
    .A(\genblk1[2].u_ce.Vld_bF$buf3 ),
    .Y(_1890_)
);

NAND2X1 _8340_ (
    .A(\genblk1[2].u_ce.Ycalc [2]),
    .B(_1890__bF$buf4),
    .Y(_1891_)
);

INVX2 _8341_ (
    .A(1'h0),
    .Y(_1892_)
);

NOR2X1 _8342_ (
    .A(1'h0),
    .B(1'h1),
    .Y(_1893_)
);

NAND2X1 _8343_ (
    .A(_1892_),
    .B(_1893_),
    .Y(_1894_)
);

INVX2 _8344_ (
    .A(_1894_),
    .Y(_1895_)
);

INVX8 _8345_ (
    .A(1'h1),
    .Y(_1896_)
);

MUX2X1 _8346_ (
    .A(\genblk1[2].u_ce.Xin12b [4]),
    .B(\genblk1[2].u_ce.Xin1 [1]),
    .S(1'h0),
    .Y(_1897_)
);

MUX2X1 _8347_ (
    .A(\genblk1[2].u_ce.Xin1 [0]),
    .B(\genblk1[2].u_ce.Xin0 [1]),
    .S(1'h0),
    .Y(_1898_)
);

MUX2X1 _8348_ (
    .A(_1898_),
    .B(_1897_),
    .S(_1896__bF$buf4),
    .Y(_1899_)
);

MUX2X1 _8349_ (
    .A(\genblk1[2].u_ce.Xin12b [8]),
    .B(\genblk1[2].u_ce.Xin12b [7]),
    .S(1'h0),
    .Y(_1900_)
);

MUX2X1 _8350_ (
    .A(\genblk1[2].u_ce.Xin12b [6]),
    .B(\genblk1[2].u_ce.Xin12b [5]),
    .S(1'h0),
    .Y(_1901_)
);

MUX2X1 _8351_ (
    .A(_1901_),
    .B(_1900_),
    .S(_1896__bF$buf3),
    .Y(_1902_)
);

MUX2X1 _8352_ (
    .A(_1902_),
    .B(_1899_),
    .S(1'h0),
    .Y(_1903_)
);

INVX1 _8353_ (
    .A(_1903_),
    .Y(_1904_)
);

MUX2X1 _8354_ (
    .A(\genblk1[2].u_ce.Xin1 [1]),
    .B(\genblk1[2].u_ce.Xin1 [0]),
    .S(1'h0),
    .Y(_1905_)
);

MUX2X1 _8355_ (
    .A(\genblk1[2].u_ce.Xin0 [1]),
    .B(\genblk1[2].u_ce.Xin0 [0]),
    .S(1'h0),
    .Y(_1906_)
);

MUX2X1 _8356_ (
    .A(_1906_),
    .B(_1905_),
    .S(_1896__bF$buf2),
    .Y(_1907_)
);

MUX2X1 _8357_ (
    .A(\genblk1[2].u_ce.Xin12b [7]),
    .B(\genblk1[2].u_ce.Xin12b [6]),
    .S(1'h0),
    .Y(_1908_)
);

MUX2X1 _8358_ (
    .A(\genblk1[2].u_ce.Xin12b [5]),
    .B(\genblk1[2].u_ce.Xin12b [4]),
    .S(1'h0),
    .Y(_1909_)
);

MUX2X1 _8359_ (
    .A(_1909_),
    .B(_1908_),
    .S(_1896__bF$buf1),
    .Y(_1910_)
);

MUX2X1 _8360_ (
    .A(_1910_),
    .B(_1907_),
    .S(1'h0),
    .Y(_1911_)
);

OAI21X1 _8361_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf4 ),
    .B(_1911_),
    .C(_1904_),
    .Y(_1912_)
);

NOR2X1 _8362_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .B(_1911_),
    .Y(_1913_)
);

NAND2X1 _8363_ (
    .A(_1903_),
    .B(_1913_),
    .Y(_1914_)
);

NAND3X1 _8364_ (
    .A(\genblk1[2].u_ce.Yin0 [1]),
    .B(_1912_),
    .C(_1914_),
    .Y(_1915_)
);

NOR2X1 _8365_ (
    .A(\genblk1[2].u_ce.Yin0 [0]),
    .B(_1911_),
    .Y(_1916_)
);

AOI21X1 _8366_ (
    .A(_1914_),
    .B(_1912_),
    .C(\genblk1[2].u_ce.Yin0 [1]),
    .Y(_1917_)
);

OAI21X1 _8367_ (
    .A(_1916_),
    .B(_1917_),
    .C(_1915_),
    .Y(_1918_)
);

INVX1 _8368_ (
    .A(\genblk1[2].u_ce.Yin1 [0]),
    .Y(_1919_)
);

MUX2X1 _8369_ (
    .A(\genblk1[2].u_ce.Xin12b [9]),
    .B(\genblk1[2].u_ce.Xin12b [8]),
    .S(1'h0),
    .Y(_1920_)
);

MUX2X1 _8370_ (
    .A(_1920_),
    .B(_1908_),
    .S(1'h1),
    .Y(_1921_)
);

AND2X2 _8371_ (
    .A(_1921_),
    .B(1'h0),
    .Y(_1922_)
);

INVX4 _8372_ (
    .A(1'h0),
    .Y(_1923_)
);

NAND2X1 _8373_ (
    .A(_1923__bF$buf3),
    .B(_1896__bF$buf0),
    .Y(_1924_)
);

NAND2X1 _8374_ (
    .A(1'h1),
    .B(_1923__bF$buf2),
    .Y(_1925_)
);

OAI22X1 _8375_ (
    .A(_1924_),
    .B(_1905_),
    .C(_1909_),
    .D(_1925_),
    .Y(_1926_)
);

INVX1 _8376_ (
    .A(\genblk1[2].u_ce.Xin1 [1]),
    .Y(_1927_)
);

NAND2X1 _8377_ (
    .A(_1892_),
    .B(_1927_),
    .Y(_1928_)
);

INVX1 _8378_ (
    .A(\genblk1[2].u_ce.Xin12b [4]),
    .Y(_1929_)
);

NAND2X1 _8379_ (
    .A(1'h0),
    .B(_1929_),
    .Y(_1930_)
);

NAND3X1 _8380_ (
    .A(1'h1),
    .B(_1930_),
    .C(_1928_),
    .Y(_1931_)
);

INVX1 _8381_ (
    .A(\genblk1[2].u_ce.Xin0 [1]),
    .Y(_1932_)
);

NAND2X1 _8382_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Xin1 [0]),
    .Y(_1933_)
);

OAI21X1 _8383_ (
    .A(1'h0),
    .B(_1932_),
    .C(_1933_),
    .Y(_1934_)
);

NAND2X1 _8384_ (
    .A(_1896__bF$buf4),
    .B(_1934_),
    .Y(_1935_)
);

NAND3X1 _8385_ (
    .A(_1923__bF$buf1),
    .B(_1931_),
    .C(_1935_),
    .Y(_1936_)
);

INVX1 _8386_ (
    .A(\genblk1[2].u_ce.Xin12b [5]),
    .Y(_1937_)
);

NAND2X1 _8387_ (
    .A(_1892_),
    .B(_1937_),
    .Y(_1938_)
);

INVX1 _8388_ (
    .A(\genblk1[2].u_ce.Xin12b [6]),
    .Y(_1939_)
);

NAND2X1 _8389_ (
    .A(1'h0),
    .B(_1939_),
    .Y(_1940_)
);

NAND3X1 _8390_ (
    .A(_1896__bF$buf3),
    .B(_1940_),
    .C(_1938_),
    .Y(_1941_)
);

INVX1 _8391_ (
    .A(\genblk1[2].u_ce.Xin12b [7]),
    .Y(_1942_)
);

NAND2X1 _8392_ (
    .A(_1892_),
    .B(_1942_),
    .Y(_1943_)
);

INVX1 _8393_ (
    .A(\genblk1[2].u_ce.Xin12b [8]),
    .Y(_1944_)
);

NAND2X1 _8394_ (
    .A(1'h0),
    .B(_1944_),
    .Y(_1945_)
);

NAND3X1 _8395_ (
    .A(1'h1),
    .B(_1945_),
    .C(_1943_),
    .Y(_1946_)
);

NAND3X1 _8396_ (
    .A(1'h0),
    .B(_1941_),
    .C(_1946_),
    .Y(_1947_)
);

INVX1 _8397_ (
    .A(\genblk1[2].u_ce.Xin1 [0]),
    .Y(_1948_)
);

NAND2X1 _8398_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Xin1 [1]),
    .Y(_1949_)
);

OAI21X1 _8399_ (
    .A(1'h0),
    .B(_1948_),
    .C(_1949_),
    .Y(_1950_)
);

NAND2X1 _8400_ (
    .A(1'h1),
    .B(_1950_),
    .Y(_1951_)
);

INVX1 _8401_ (
    .A(\genblk1[2].u_ce.Xin0 [0]),
    .Y(_1952_)
);

NAND2X1 _8402_ (
    .A(\genblk1[2].u_ce.Xin0 [1]),
    .B(1'h0),
    .Y(_1953_)
);

OAI21X1 _8403_ (
    .A(1'h0),
    .B(_1952_),
    .C(_1953_),
    .Y(_1954_)
);

NAND2X1 _8404_ (
    .A(_1896__bF$buf2),
    .B(_1954_),
    .Y(_1955_)
);

NAND3X1 _8405_ (
    .A(_1923__bF$buf0),
    .B(_1951_),
    .C(_1955_),
    .Y(_1956_)
);

NAND2X1 _8406_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Xin12b [5]),
    .Y(_1957_)
);

OAI21X1 _8407_ (
    .A(1'h0),
    .B(_1929_),
    .C(_1957_),
    .Y(_1958_)
);

NAND2X1 _8408_ (
    .A(_1896__bF$buf1),
    .B(_1958_),
    .Y(_1959_)
);

NAND2X1 _8409_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Xin12b [7]),
    .Y(_1960_)
);

OAI21X1 _8410_ (
    .A(1'h0),
    .B(_1939_),
    .C(_1960_),
    .Y(_1961_)
);

NAND2X1 _8411_ (
    .A(1'h1),
    .B(_1961_),
    .Y(_1962_)
);

NAND3X1 _8412_ (
    .A(1'h0),
    .B(_1959_),
    .C(_1962_),
    .Y(_1963_)
);

AOI22X1 _8413_ (
    .A(_1936_),
    .B(_1947_),
    .C(_1956_),
    .D(_1963_),
    .Y(_1964_)
);

NOR2X1 _8414_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1964_),
    .Y(_1965_)
);

OAI21X1 _8415_ (
    .A(_1922_),
    .B(_1926_),
    .C(_1965_),
    .Y(_1966_)
);

AOI21X1 _8416_ (
    .A(1'h0),
    .B(_1921_),
    .C(_1926_),
    .Y(_1967_)
);

OAI21X1 _8417_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1964_),
    .C(_1967_),
    .Y(_1968_)
);

NAND3X1 _8418_ (
    .A(_1919_),
    .B(_1968_),
    .C(_1966_),
    .Y(_1969_)
);

NAND2X1 _8419_ (
    .A(_1967_),
    .B(_1965_),
    .Y(_1970_)
);

OAI22X1 _8420_ (
    .A(_1922_),
    .B(_1926_),
    .C(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .D(_1964_),
    .Y(_1971_)
);

NAND3X1 _8421_ (
    .A(\genblk1[2].u_ce.Yin1 [0]),
    .B(_1971_),
    .C(_1970_),
    .Y(_1972_)
);

NAND3X1 _8422_ (
    .A(_1969_),
    .B(_1972_),
    .C(_1918_),
    .Y(_1973_)
);

INVX1 _8423_ (
    .A(\genblk1[2].u_ce.Yin0 [1]),
    .Y(_1974_)
);

NAND2X1 _8424_ (
    .A(_1904_),
    .B(_1913_),
    .Y(_1975_)
);

OAI21X1 _8425_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf4 ),
    .B(_1911_),
    .C(_1903_),
    .Y(_1976_)
);

AOI21X1 _8426_ (
    .A(_1975_),
    .B(_1976_),
    .C(_1974_),
    .Y(_1977_)
);

INVX1 _8427_ (
    .A(_1916_),
    .Y(_1978_)
);

NAND3X1 _8428_ (
    .A(_1974_),
    .B(_1976_),
    .C(_1975_),
    .Y(_1979_)
);

AOI21X1 _8429_ (
    .A(_1978_),
    .B(_1979_),
    .C(_1977_),
    .Y(_1980_)
);

AOI21X1 _8430_ (
    .A(_1970_),
    .B(_1971_),
    .C(\genblk1[2].u_ce.Yin1 [0]),
    .Y(_1981_)
);

AOI21X1 _8431_ (
    .A(_1966_),
    .B(_1968_),
    .C(_1919_),
    .Y(_1982_)
);

OAI21X1 _8432_ (
    .A(_1981_),
    .B(_1982_),
    .C(_1980_),
    .Y(_1983_)
);

AOI21X1 _8433_ (
    .A(_1973_),
    .B(_1983_),
    .C(_1895_),
    .Y(_1984_)
);

INVX8 _8434_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_1985_)
);

NAND3X1 _8435_ (
    .A(_1923__bF$buf3),
    .B(_1892_),
    .C(_1985__bF$buf5),
    .Y(_1986_)
);

OAI21X1 _8436_ (
    .A(1'h1),
    .B(_1986_),
    .C(\genblk1[2].u_ce.Vld_bF$buf2 ),
    .Y(_1987_)
);

OAI21X1 _8437_ (
    .A(_1987_),
    .B(_1984_),
    .C(_1891_),
    .Y(_1734_)
);

INVX1 _8438_ (
    .A(\genblk1[2].u_ce.Ycalc [3]),
    .Y(_1988_)
);

INVX1 _8439_ (
    .A(\genblk1[2].u_ce.Xin12b [9]),
    .Y(_1989_)
);

NAND2X1 _8440_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Xin12b [10]),
    .Y(_1990_)
);

OAI21X1 _8441_ (
    .A(1'h0),
    .B(_1989_),
    .C(_1990_),
    .Y(_1991_)
);

NAND2X1 _8442_ (
    .A(1'h1),
    .B(_1991_),
    .Y(_1992_)
);

OAI21X1 _8443_ (
    .A(1'h1),
    .B(_1900_),
    .C(_1992_),
    .Y(_1993_)
);

OAI22X1 _8444_ (
    .A(_1924_),
    .B(_1897_),
    .C(_1901_),
    .D(_1925_),
    .Y(_1994_)
);

AOI21X1 _8445_ (
    .A(_1993_),
    .B(1'h0),
    .C(_1994_),
    .Y(_1995_)
);

NAND3X1 _8446_ (
    .A(_1967_),
    .B(_1903_),
    .C(_1911_),
    .Y(_1996_)
);

INVX1 _8447_ (
    .A(_1996_),
    .Y(_1997_)
);

NOR2X1 _8448_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_1997_),
    .Y(_1998_)
);

NAND2X1 _8449_ (
    .A(_1995_),
    .B(_1998_),
    .Y(_1999_)
);

INVX1 _8450_ (
    .A(_1995_),
    .Y(_2000_)
);

OAI21X1 _8451_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .B(_1997_),
    .C(_2000_),
    .Y(_2001_)
);

AOI21X1 _8452_ (
    .A(_1999_),
    .B(_2001_),
    .C(\genblk1[2].u_ce.Yin1 [1]),
    .Y(_2002_)
);

AOI21X1 _8453_ (
    .A(_1918_),
    .B(_1969_),
    .C(_1982_),
    .Y(_2003_)
);

NAND3X1 _8454_ (
    .A(\genblk1[2].u_ce.Yin1 [1]),
    .B(_2001_),
    .C(_1999_),
    .Y(_2004_)
);

NAND2X1 _8455_ (
    .A(_2004_),
    .B(_2003_),
    .Y(_2005_)
);

OAI21X1 _8456_ (
    .A(_1981_),
    .B(_1980_),
    .C(_1972_),
    .Y(_2006_)
);

INVX1 _8457_ (
    .A(\genblk1[2].u_ce.Yin1 [1]),
    .Y(_2007_)
);

NAND2X1 _8458_ (
    .A(_2000_),
    .B(_1998_),
    .Y(_2008_)
);

OAI21X1 _8459_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .B(_1997_),
    .C(_1995_),
    .Y(_2009_)
);

AOI21X1 _8460_ (
    .A(_2008_),
    .B(_2009_),
    .C(_2007_),
    .Y(_2010_)
);

OAI21X1 _8461_ (
    .A(_2002_),
    .B(_2010_),
    .C(_2006_),
    .Y(_2011_)
);

OAI21X1 _8462_ (
    .A(_2002_),
    .B(_2005_),
    .C(_2011_),
    .Y(_2012_)
);

OAI21X1 _8463_ (
    .A(_1985__bF$buf4),
    .B(_1894_),
    .C(\genblk1[2].u_ce.Vld_bF$buf1 ),
    .Y(_2013_)
);

INVX1 _8464_ (
    .A(_2013_),
    .Y(_2014_)
);

OAI21X1 _8465_ (
    .A(_1895_),
    .B(_2012_),
    .C(_2014_),
    .Y(_2015_)
);

OAI21X1 _8466_ (
    .A(_1988_),
    .B(\genblk1[2].u_ce.Vld_bF$buf0 ),
    .C(_2015_),
    .Y(_1735_)
);

INVX1 _8467_ (
    .A(_1987_),
    .Y(_2016_)
);

INVX1 _8468_ (
    .A(\genblk1[2].u_ce.Yin12b [4]),
    .Y(_2017_)
);

NAND3X1 _8469_ (
    .A(_1967_),
    .B(_1995_),
    .C(_1964_),
    .Y(_2018_)
);

INVX1 _8470_ (
    .A(\genblk1[2].u_ce.Xin12b [10]),
    .Y(_2019_)
);

NAND2X1 _8471_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Xin12b [11]),
    .Y(_2020_)
);

OAI21X1 _8472_ (
    .A(1'h0),
    .B(_2019_),
    .C(_2020_),
    .Y(_2021_)
);

NAND2X1 _8473_ (
    .A(_1896__bF$buf0),
    .B(_1920_),
    .Y(_2022_)
);

OAI21X1 _8474_ (
    .A(_1896__bF$buf4),
    .B(_2021_),
    .C(_2022_),
    .Y(_2023_)
);

NAND2X1 _8475_ (
    .A(_1923__bF$buf2),
    .B(_1910_),
    .Y(_2024_)
);

OAI21X1 _8476_ (
    .A(_1923__bF$buf1),
    .B(_2023_),
    .C(_2024_),
    .Y(_2025_)
);

INVX1 _8477_ (
    .A(_2025_),
    .Y(_2026_)
);

NAND3X1 _8478_ (
    .A(_1985__bF$buf3),
    .B(_2026_),
    .C(_2018_),
    .Y(_2027_)
);

INVX1 _8479_ (
    .A(_2027_),
    .Y(_2028_)
);

AOI21X1 _8480_ (
    .A(_2018_),
    .B(_1985__bF$buf2),
    .C(_2026_),
    .Y(_2029_)
);

OAI21X1 _8481_ (
    .A(_2029_),
    .B(_2028_),
    .C(_2017_),
    .Y(_2030_)
);

OAI21X1 _8482_ (
    .A(_1996_),
    .B(_2000_),
    .C(_1985__bF$buf1),
    .Y(_2031_)
);

NAND2X1 _8483_ (
    .A(_2025_),
    .B(_2031_),
    .Y(_2032_)
);

NAND3X1 _8484_ (
    .A(\genblk1[2].u_ce.Yin12b [4]),
    .B(_2027_),
    .C(_2032_),
    .Y(_2033_)
);

NAND2X1 _8485_ (
    .A(_2033_),
    .B(_2030_),
    .Y(_2034_)
);

INVX1 _8486_ (
    .A(_2002_),
    .Y(_2035_)
);

OAI21X1 _8487_ (
    .A(_2010_),
    .B(_2006_),
    .C(_2035_),
    .Y(_2036_)
);

AOI21X1 _8488_ (
    .A(_2036_),
    .B(_2034_),
    .C(_1895_),
    .Y(_2037_)
);

OAI21X1 _8489_ (
    .A(_2034_),
    .B(_2036_),
    .C(_2037_),
    .Y(_2038_)
);

AOI22X1 _8490_ (
    .A(_1853_),
    .B(_1890__bF$buf3),
    .C(_2038_),
    .D(_2016_),
    .Y(_1736_)
);

INVX1 _8491_ (
    .A(_2033_),
    .Y(_2039_)
);

AOI21X1 _8492_ (
    .A(_2003_),
    .B(_2004_),
    .C(_2002_),
    .Y(_2040_)
);

AOI21X1 _8493_ (
    .A(_2040_),
    .B(_2030_),
    .C(_2039_),
    .Y(_2041_)
);

INVX1 _8494_ (
    .A(\genblk1[2].u_ce.Yin12b [5]),
    .Y(_2042_)
);

NAND3X1 _8495_ (
    .A(_1995_),
    .B(_2026_),
    .C(_1997_),
    .Y(_2043_)
);

INVX1 _8496_ (
    .A(\genblk1[2].u_ce.Xin12b [11]),
    .Y(_2044_)
);

NOR2X1 _8497_ (
    .A(_1896__bF$buf3),
    .B(_2044_),
    .Y(_2045_)
);

AOI21X1 _8498_ (
    .A(_1896__bF$buf2),
    .B(_1991_),
    .C(_2045_),
    .Y(_2046_)
);

NAND2X1 _8499_ (
    .A(_1923__bF$buf0),
    .B(_1902_),
    .Y(_2047_)
);

OAI21X1 _8500_ (
    .A(_1923__bF$buf3),
    .B(_2046_),
    .C(_2047_),
    .Y(_2048_)
);

NAND3X1 _8501_ (
    .A(_1985__bF$buf0),
    .B(_2048_),
    .C(_2043_),
    .Y(_2049_)
);

INVX1 _8502_ (
    .A(_2048_),
    .Y(_2050_)
);

OAI21X1 _8503_ (
    .A(_2025_),
    .B(_2018_),
    .C(_1985__bF$buf5),
    .Y(_2051_)
);

NAND2X1 _8504_ (
    .A(_2050_),
    .B(_2051_),
    .Y(_2052_)
);

NAND3X1 _8505_ (
    .A(_2042_),
    .B(_2052_),
    .C(_2049_),
    .Y(_2053_)
);

NAND3X1 _8506_ (
    .A(_1985__bF$buf4),
    .B(_2050_),
    .C(_2043_),
    .Y(_2054_)
);

NAND2X1 _8507_ (
    .A(_2048_),
    .B(_2051_),
    .Y(_2055_)
);

NAND3X1 _8508_ (
    .A(\genblk1[2].u_ce.Yin12b [5]),
    .B(_2055_),
    .C(_2054_),
    .Y(_2056_)
);

NAND2X1 _8509_ (
    .A(_2053_),
    .B(_2056_),
    .Y(_2057_)
);

INVX1 _8510_ (
    .A(_2057_),
    .Y(_2058_)
);

NOR2X1 _8511_ (
    .A(_2058_),
    .B(_2041_),
    .Y(_2059_)
);

OAI21X1 _8512_ (
    .A(_2034_),
    .B(_2036_),
    .C(_2033_),
    .Y(_2060_)
);

OAI21X1 _8513_ (
    .A(_2057_),
    .B(_2060_),
    .C(_1894_),
    .Y(_2061_)
);

OAI21X1 _8514_ (
    .A(_2061_),
    .B(_2059_),
    .C(_2016_),
    .Y(_2062_)
);

OAI21X1 _8515_ (
    .A(_1861_),
    .B(\genblk1[2].u_ce.Vld_bF$buf4 ),
    .C(_2062_),
    .Y(_1737_)
);

NOR2X1 _8516_ (
    .A(_2034_),
    .B(_2057_),
    .Y(_2063_)
);

OAI21X1 _8517_ (
    .A(_2033_),
    .B(_2057_),
    .C(_2056_),
    .Y(_2064_)
);

AOI21X1 _8518_ (
    .A(_2063_),
    .B(_2040_),
    .C(_2064_),
    .Y(_2065_)
);

INVX1 _8519_ (
    .A(\genblk1[2].u_ce.Yin12b [6]),
    .Y(_2066_)
);

NOR2X1 _8520_ (
    .A(_2025_),
    .B(_2018_),
    .Y(_2067_)
);

NAND2X1 _8521_ (
    .A(_2050_),
    .B(_2067_),
    .Y(_2068_)
);

AOI21X1 _8522_ (
    .A(_1896__bF$buf1),
    .B(_2021_),
    .C(_2045_),
    .Y(_2069_)
);

NAND2X1 _8523_ (
    .A(_1923__bF$buf2),
    .B(_1921_),
    .Y(_2070_)
);

OAI21X1 _8524_ (
    .A(_1923__bF$buf1),
    .B(_2069_),
    .C(_2070_),
    .Y(_2071_)
);

NAND3X1 _8525_ (
    .A(_1985__bF$buf3),
    .B(_2071_),
    .C(_2068_),
    .Y(_2072_)
);

NOR3X1 _8526_ (
    .A(_2025_),
    .B(_2048_),
    .C(_2018_),
    .Y(_2073_)
);

INVX1 _8527_ (
    .A(_2071_),
    .Y(_2074_)
);

OAI21X1 _8528_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf4 ),
    .B(_2073_),
    .C(_2074_),
    .Y(_2075_)
);

NAND3X1 _8529_ (
    .A(_2066_),
    .B(_2075_),
    .C(_2072_),
    .Y(_2076_)
);

NAND3X1 _8530_ (
    .A(_1985__bF$buf2),
    .B(_2074_),
    .C(_2068_),
    .Y(_2077_)
);

OAI21X1 _8531_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2073_),
    .C(_2071_),
    .Y(_2078_)
);

NAND3X1 _8532_ (
    .A(\genblk1[2].u_ce.Yin12b [6]),
    .B(_2078_),
    .C(_2077_),
    .Y(_2079_)
);

AND2X2 _8533_ (
    .A(_2076_),
    .B(_2079_),
    .Y(_2080_)
);

INVX1 _8534_ (
    .A(_2080_),
    .Y(_2081_)
);

AOI21X1 _8535_ (
    .A(_2065_),
    .B(_2081_),
    .C(_1895_),
    .Y(_2082_)
);

OAI21X1 _8536_ (
    .A(_2065_),
    .B(_2081_),
    .C(_2082_),
    .Y(_2083_)
);

AOI22X1 _8537_ (
    .A(_1852_),
    .B(_1890__bF$buf2),
    .C(_2083_),
    .D(_2016_),
    .Y(_1738_)
);

AND2X2 _8538_ (
    .A(_2030_),
    .B(_2033_),
    .Y(_2084_)
);

NAND3X1 _8539_ (
    .A(_2053_),
    .B(_2056_),
    .C(_2084_),
    .Y(_2085_)
);

INVX1 _8540_ (
    .A(_2056_),
    .Y(_2086_)
);

AOI21X1 _8541_ (
    .A(_2039_),
    .B(_2053_),
    .C(_2086_),
    .Y(_2087_)
);

OAI21X1 _8542_ (
    .A(_2036_),
    .B(_2085_),
    .C(_2087_),
    .Y(_2088_)
);

INVX1 _8543_ (
    .A(_2079_),
    .Y(_2089_)
);

AOI21X1 _8544_ (
    .A(_2088_),
    .B(_2076_),
    .C(_2089_),
    .Y(_2090_)
);

INVX1 _8545_ (
    .A(\genblk1[2].u_ce.Yin12b [7]),
    .Y(_2091_)
);

NAND2X1 _8546_ (
    .A(_2074_),
    .B(_2073_),
    .Y(_2092_)
);

NOR2X1 _8547_ (
    .A(_1923__bF$buf0),
    .B(_2044_),
    .Y(_2093_)
);

AOI21X1 _8548_ (
    .A(_1993_),
    .B(_1923__bF$buf3),
    .C(_2093_),
    .Y(_2094_)
);

INVX1 _8549_ (
    .A(_2094_),
    .Y(_2095_)
);

NAND3X1 _8550_ (
    .A(_1985__bF$buf1),
    .B(_2095_),
    .C(_2092_),
    .Y(_2096_)
);

AND2X2 _8551_ (
    .A(_2073_),
    .B(_2074_),
    .Y(_2097_)
);

OAI21X1 _8552_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2097_),
    .C(_2094_),
    .Y(_2098_)
);

NAND3X1 _8553_ (
    .A(_2091_),
    .B(_2096_),
    .C(_2098_),
    .Y(_2099_)
);

NAND3X1 _8554_ (
    .A(_1985__bF$buf0),
    .B(_2094_),
    .C(_2092_),
    .Y(_2100_)
);

OAI21X1 _8555_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .B(_2097_),
    .C(_2095_),
    .Y(_2101_)
);

NAND3X1 _8556_ (
    .A(\genblk1[2].u_ce.Yin12b [7]),
    .B(_2100_),
    .C(_2101_),
    .Y(_2102_)
);

AND2X2 _8557_ (
    .A(_2099_),
    .B(_2102_),
    .Y(_2103_)
);

NOR2X1 _8558_ (
    .A(_2103_),
    .B(_2090_),
    .Y(_2104_)
);

NAND2X1 _8559_ (
    .A(_1892_),
    .B(_1896__bF$buf0),
    .Y(_2105_)
);

NAND2X1 _8560_ (
    .A(_2103_),
    .B(_2090_),
    .Y(_2106_)
);

OAI21X1 _8561_ (
    .A(1'h0),
    .B(_2105_),
    .C(_2106_),
    .Y(_2107_)
);

OAI21X1 _8562_ (
    .A(_2104_),
    .B(_2107_),
    .C(_2014_),
    .Y(_2108_)
);

OAI21X1 _8563_ (
    .A(_1860_),
    .B(\genblk1[2].u_ce.Vld_bF$buf3 ),
    .C(_2108_),
    .Y(_1739_)
);

INVX1 _8564_ (
    .A(\genblk1[2].u_ce.Ycalc [8]),
    .Y(_2109_)
);

AOI21X1 _8565_ (
    .A(_2098_),
    .B(_2096_),
    .C(_2091_),
    .Y(_2110_)
);

OAI21X1 _8566_ (
    .A(_2089_),
    .B(_2110_),
    .C(_2099_),
    .Y(_2111_)
);

NAND3X1 _8567_ (
    .A(_2080_),
    .B(_2103_),
    .C(_2088_),
    .Y(_2112_)
);

INVX1 _8568_ (
    .A(\genblk1[2].u_ce.Yin12b [8]),
    .Y(_2113_)
);

NAND3X1 _8569_ (
    .A(_2074_),
    .B(_2094_),
    .C(_2073_),
    .Y(_2114_)
);

INVX1 _8570_ (
    .A(_2093_),
    .Y(_2115_)
);

OAI21X1 _8571_ (
    .A(1'h0),
    .B(_2023_),
    .C(_2115_),
    .Y(_2116_)
);

NAND3X1 _8572_ (
    .A(_1985__bF$buf5),
    .B(_2116_),
    .C(_2114_),
    .Y(_2117_)
);

INVX1 _8573_ (
    .A(_2116_),
    .Y(_2118_)
);

NAND2X1 _8574_ (
    .A(_1985__bF$buf4),
    .B(_2114_),
    .Y(_2119_)
);

NAND2X1 _8575_ (
    .A(_2118_),
    .B(_2119_),
    .Y(_2120_)
);

NAND3X1 _8576_ (
    .A(_2113_),
    .B(_2117_),
    .C(_2120_),
    .Y(_2121_)
);

NAND3X1 _8577_ (
    .A(_1985__bF$buf3),
    .B(_2118_),
    .C(_2114_),
    .Y(_2122_)
);

NAND2X1 _8578_ (
    .A(_2116_),
    .B(_2119_),
    .Y(_2123_)
);

NAND3X1 _8579_ (
    .A(\genblk1[2].u_ce.Yin12b [8]),
    .B(_2122_),
    .C(_2123_),
    .Y(_2124_)
);

AND2X2 _8580_ (
    .A(_2121_),
    .B(_2124_),
    .Y(_2125_)
);

INVX1 _8581_ (
    .A(_2125_),
    .Y(_2126_)
);

AOI21X1 _8582_ (
    .A(_2112_),
    .B(_2111_),
    .C(_2126_),
    .Y(_2127_)
);

NAND3X1 _8583_ (
    .A(_2099_),
    .B(_2102_),
    .C(_2080_),
    .Y(_2128_)
);

OAI21X1 _8584_ (
    .A(_2128_),
    .B(_2065_),
    .C(_2111_),
    .Y(_2129_)
);

OAI21X1 _8585_ (
    .A(_2125_),
    .B(_2129_),
    .C(_1894_),
    .Y(_2130_)
);

OR2X2 _8586_ (
    .A(_2130_),
    .B(_2127_),
    .Y(_2131_)
);

AOI22X1 _8587_ (
    .A(_2109_),
    .B(_1890__bF$buf1),
    .C(_2131_),
    .D(_2014_),
    .Y(_1740_)
);

INVX1 _8588_ (
    .A(\genblk1[2].u_ce.Ycalc [9]),
    .Y(_2132_)
);

INVX1 _8589_ (
    .A(_2124_),
    .Y(_2133_)
);

NOR2X1 _8590_ (
    .A(_2133_),
    .B(_2127_),
    .Y(_2134_)
);

INVX1 _8591_ (
    .A(\genblk1[2].u_ce.Yin12b [9]),
    .Y(_2135_)
);

OAI21X1 _8592_ (
    .A(1'h0),
    .B(_2046_),
    .C(_2115_),
    .Y(_2136_)
);

INVX1 _8593_ (
    .A(_2136_),
    .Y(_2137_)
);

OAI21X1 _8594_ (
    .A(_2116_),
    .B(_2114_),
    .C(_1985__bF$buf2),
    .Y(_2138_)
);

NAND2X1 _8595_ (
    .A(_2137_),
    .B(_2138_),
    .Y(_2139_)
);

NAND3X1 _8596_ (
    .A(_2094_),
    .B(_2118_),
    .C(_2097_),
    .Y(_2140_)
);

NAND3X1 _8597_ (
    .A(_1985__bF$buf1),
    .B(_2136_),
    .C(_2140_),
    .Y(_2141_)
);

NAND3X1 _8598_ (
    .A(_2135_),
    .B(_2139_),
    .C(_2141_),
    .Y(_2142_)
);

AND2X2 _8599_ (
    .A(_2138_),
    .B(_2137_),
    .Y(_2143_)
);

NOR2X1 _8600_ (
    .A(_2137_),
    .B(_2138_),
    .Y(_2144_)
);

OAI21X1 _8601_ (
    .A(_2144_),
    .B(_2143_),
    .C(\genblk1[2].u_ce.Yin12b [9]),
    .Y(_2145_)
);

NAND2X1 _8602_ (
    .A(_2142_),
    .B(_2145_),
    .Y(_2146_)
);

AOI21X1 _8603_ (
    .A(_2134_),
    .B(_2146_),
    .C(_1895_),
    .Y(_2147_)
);

OAI21X1 _8604_ (
    .A(_2134_),
    .B(_2146_),
    .C(_2147_),
    .Y(_2148_)
);

AOI22X1 _8605_ (
    .A(_2132_),
    .B(_1890__bF$buf0),
    .C(_2148_),
    .D(_2014_),
    .Y(_1741_)
);

OAI21X1 _8606_ (
    .A(_2124_),
    .B(_2146_),
    .C(_2145_),
    .Y(_2149_)
);

NAND3X1 _8607_ (
    .A(_2142_),
    .B(_2145_),
    .C(_2125_),
    .Y(_2150_)
);

AOI21X1 _8608_ (
    .A(_2111_),
    .B(_2112_),
    .C(_2150_),
    .Y(_2151_)
);

INVX1 _8609_ (
    .A(\genblk1[2].u_ce.Yin12b [10]),
    .Y(_2152_)
);

OAI21X1 _8610_ (
    .A(1'h0),
    .B(_2069_),
    .C(_2115_),
    .Y(_2153_)
);

INVX1 _8611_ (
    .A(_2153_),
    .Y(_2154_)
);

OAI21X1 _8612_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2137_),
    .C(_2138_),
    .Y(_2155_)
);

NAND2X1 _8613_ (
    .A(_2154_),
    .B(_2155_),
    .Y(_2156_)
);

OAI21X1 _8614_ (
    .A(_2136_),
    .B(_2140_),
    .C(_1985__bF$buf0),
    .Y(_2157_)
);

NAND2X1 _8615_ (
    .A(_2153_),
    .B(_2157_),
    .Y(_2158_)
);

NAND2X1 _8616_ (
    .A(_2156_),
    .B(_2158_),
    .Y(_2159_)
);

NAND2X1 _8617_ (
    .A(_2152_),
    .B(_2159_),
    .Y(_2160_)
);

NAND3X1 _8618_ (
    .A(\genblk1[2].u_ce.Yin12b [10]),
    .B(_2156_),
    .C(_2158_),
    .Y(_2161_)
);

AND2X2 _8619_ (
    .A(_2160_),
    .B(_2161_),
    .Y(_2162_)
);

OAI21X1 _8620_ (
    .A(_2149_),
    .B(_2151_),
    .C(_2162_),
    .Y(_2163_)
);

INVX1 _8621_ (
    .A(_2145_),
    .Y(_2164_)
);

AOI21X1 _8622_ (
    .A(_2133_),
    .B(_2142_),
    .C(_2164_),
    .Y(_2165_)
);

AND2X2 _8623_ (
    .A(_2145_),
    .B(_2142_),
    .Y(_2166_)
);

NAND3X1 _8624_ (
    .A(_2125_),
    .B(_2166_),
    .C(_2129_),
    .Y(_2167_)
);

NAND2X1 _8625_ (
    .A(_2161_),
    .B(_2160_),
    .Y(_2168_)
);

NAND3X1 _8626_ (
    .A(_2165_),
    .B(_2168_),
    .C(_2167_),
    .Y(_2169_)
);

NAND3X1 _8627_ (
    .A(_1894_),
    .B(_2169_),
    .C(_2163_),
    .Y(_2170_)
);

AOI22X1 _8628_ (
    .A(_1849_),
    .B(_1890__bF$buf4),
    .C(_2170_),
    .D(_2016_),
    .Y(_1742_)
);

INVX1 _8629_ (
    .A(_2161_),
    .Y(_2171_)
);

AOI21X1 _8630_ (
    .A(_2167_),
    .B(_2165_),
    .C(_2168_),
    .Y(_2172_)
);

OAI21X1 _8631_ (
    .A(_2153_),
    .B(_2155_),
    .C(_1985__bF$buf5),
    .Y(_2173_)
);

INVX1 _8632_ (
    .A(_2173_),
    .Y(_2174_)
);

NAND2X1 _8633_ (
    .A(\genblk1[2].u_ce.Yin12b [11]),
    .B(_2044_),
    .Y(_2175_)
);

INVX1 _8634_ (
    .A(\genblk1[2].u_ce.Yin12b [11]),
    .Y(_2176_)
);

NAND2X1 _8635_ (
    .A(\genblk1[2].u_ce.Xin12b [11]),
    .B(_2176_),
    .Y(_2177_)
);

NAND2X1 _8636_ (
    .A(_2175_),
    .B(_2177_),
    .Y(_2178_)
);

OR2X2 _8637_ (
    .A(_2174_),
    .B(_2178_),
    .Y(_2179_)
);

NAND2X1 _8638_ (
    .A(_2178_),
    .B(_2174_),
    .Y(_2180_)
);

NAND2X1 _8639_ (
    .A(_2180_),
    .B(_2179_),
    .Y(_2181_)
);

OAI21X1 _8640_ (
    .A(_2171_),
    .B(_2172_),
    .C(_2181_),
    .Y(_2182_)
);

INVX1 _8641_ (
    .A(_2181_),
    .Y(_2183_)
);

NAND3X1 _8642_ (
    .A(_2161_),
    .B(_2183_),
    .C(_2163_),
    .Y(_2184_)
);

NAND3X1 _8643_ (
    .A(_1894_),
    .B(_2184_),
    .C(_2182_),
    .Y(_2185_)
);

AOI22X1 _8644_ (
    .A(_1857_),
    .B(_1890__bF$buf3),
    .C(_2185_),
    .D(_2014_),
    .Y(_1743_)
);

INVX1 _8645_ (
    .A(\genblk1[2].u_ce.Ycalc [0]),
    .Y(_2186_)
);

OAI21X1 _8646_ (
    .A(1'h0),
    .B(_2105_),
    .C(\genblk1[2].u_ce.Vld_bF$buf2 ),
    .Y(_2187_)
);

INVX2 _8647_ (
    .A(_2187_),
    .Y(_2188_)
);

INVX1 _8648_ (
    .A(\genblk1[2].u_ce.Yin0 [0]),
    .Y(_2189_)
);

AOI21X1 _8649_ (
    .A(_1956_),
    .B(_1963_),
    .C(_2189_),
    .Y(_2190_)
);

OAI21X1 _8650_ (
    .A(_2190_),
    .B(_1916_),
    .C(_2188_),
    .Y(_2191_)
);

OAI21X1 _8651_ (
    .A(_2186_),
    .B(\genblk1[2].u_ce.Vld_bF$buf1 ),
    .C(_2191_),
    .Y(_1744_)
);

NAND2X1 _8652_ (
    .A(\genblk1[2].u_ce.Ycalc [1]),
    .B(_1890__bF$buf2),
    .Y(_2192_)
);

NAND3X1 _8653_ (
    .A(_1978_),
    .B(_1915_),
    .C(_1979_),
    .Y(_2193_)
);

OAI21X1 _8654_ (
    .A(_1977_),
    .B(_1917_),
    .C(_1916_),
    .Y(_2194_)
);

AOI21X1 _8655_ (
    .A(_2194_),
    .B(_2193_),
    .C(_1895_),
    .Y(_2195_)
);

OAI21X1 _8656_ (
    .A(_1890__bF$buf1),
    .B(_2195_),
    .C(_2192_),
    .Y(_1745_)
);

NAND2X1 _8657_ (
    .A(\genblk1[2].u_ce.Xcalc [0]),
    .B(_1890__bF$buf0),
    .Y(_2196_)
);

MUX2X1 _8658_ (
    .A(\genblk1[2].u_ce.Yin12b [7]),
    .B(\genblk1[2].u_ce.Yin12b [6]),
    .S(1'h0),
    .Y(_2197_)
);

NAND2X1 _8659_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin12b [5]),
    .Y(_2198_)
);

OAI21X1 _8660_ (
    .A(1'h0),
    .B(_2017_),
    .C(_2198_),
    .Y(_2199_)
);

NAND2X1 _8661_ (
    .A(_1896__bF$buf4),
    .B(_2199_),
    .Y(_2200_)
);

OAI21X1 _8662_ (
    .A(_1896__bF$buf3),
    .B(_2197_),
    .C(_2200_),
    .Y(_2201_)
);

NAND2X1 _8663_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin1 [1]),
    .Y(_2202_)
);

OAI21X1 _8664_ (
    .A(1'h0),
    .B(_1919_),
    .C(_2202_),
    .Y(_2203_)
);

NAND2X1 _8665_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin0 [1]),
    .Y(_2204_)
);

OAI21X1 _8666_ (
    .A(1'h0),
    .B(_2189_),
    .C(_2204_),
    .Y(_2205_)
);

MUX2X1 _8667_ (
    .A(_2205_),
    .B(_2203_),
    .S(_1896__bF$buf2),
    .Y(_2206_)
);

NAND2X1 _8668_ (
    .A(_1923__bF$buf2),
    .B(_2206_),
    .Y(_2207_)
);

OAI21X1 _8669_ (
    .A(_1923__bF$buf1),
    .B(_2201_),
    .C(_2207_),
    .Y(_2208_)
);

INVX1 _8670_ (
    .A(_2208_),
    .Y(_2209_)
);

NOR2X1 _8671_ (
    .A(\genblk1[2].u_ce.Xin0 [0]),
    .B(_2209_),
    .Y(_2210_)
);

OAI21X1 _8672_ (
    .A(_1952_),
    .B(_2208_),
    .C(_2188_),
    .Y(_2211_)
);

OAI21X1 _8673_ (
    .A(_2211_),
    .B(_2210_),
    .C(_2196_),
    .Y(_1746_)
);

NAND2X1 _8674_ (
    .A(\genblk1[2].u_ce.Xcalc [1]),
    .B(_1890__bF$buf4),
    .Y(_2212_)
);

NOR2X1 _8675_ (
    .A(_1952_),
    .B(_2208_),
    .Y(_2213_)
);

NAND2X1 _8676_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin12b [4]),
    .Y(_2214_)
);

OAI21X1 _8677_ (
    .A(1'h0),
    .B(_2007_),
    .C(_2214_),
    .Y(_2215_)
);

NAND2X1 _8678_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin1 [0]),
    .Y(_2216_)
);

OAI21X1 _8679_ (
    .A(1'h0),
    .B(_1974_),
    .C(_2216_),
    .Y(_2217_)
);

MUX2X1 _8680_ (
    .A(_2217_),
    .B(_2215_),
    .S(_1896__bF$buf1),
    .Y(_2218_)
);

NAND2X1 _8681_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin12b [8]),
    .Y(_2219_)
);

OAI21X1 _8682_ (
    .A(1'h0),
    .B(_2091_),
    .C(_2219_),
    .Y(_2220_)
);

NAND2X1 _8683_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin12b [6]),
    .Y(_2221_)
);

OAI21X1 _8684_ (
    .A(1'h0),
    .B(_2042_),
    .C(_2221_),
    .Y(_2222_)
);

MUX2X1 _8685_ (
    .A(_2222_),
    .B(_2220_),
    .S(_1896__bF$buf0),
    .Y(_2223_)
);

MUX2X1 _8686_ (
    .A(_2223_),
    .B(_2218_),
    .S(1'h0),
    .Y(_2224_)
);

NOR2X1 _8687_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf4 ),
    .B(_2208_),
    .Y(_2225_)
);

NAND2X1 _8688_ (
    .A(_2224_),
    .B(_2225_),
    .Y(_2226_)
);

NAND2X1 _8689_ (
    .A(_1923__bF$buf0),
    .B(_2218_),
    .Y(_2227_)
);

NAND2X1 _8690_ (
    .A(1'h0),
    .B(_2223_),
    .Y(_2228_)
);

NAND2X1 _8691_ (
    .A(_2227_),
    .B(_2228_),
    .Y(_2229_)
);

OAI21X1 _8692_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2208_),
    .C(_2229_),
    .Y(_2230_)
);

NAND3X1 _8693_ (
    .A(\genblk1[2].u_ce.Xin0 [1]),
    .B(_2230_),
    .C(_2226_),
    .Y(_2231_)
);

OAI21X1 _8694_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2208_),
    .C(_2224_),
    .Y(_2232_)
);

NAND2X1 _8695_ (
    .A(_2229_),
    .B(_2225_),
    .Y(_2233_)
);

NAND3X1 _8696_ (
    .A(_1932_),
    .B(_2232_),
    .C(_2233_),
    .Y(_2234_)
);

NAND3X1 _8697_ (
    .A(_2213_),
    .B(_2231_),
    .C(_2234_),
    .Y(_2235_)
);

INVX1 _8698_ (
    .A(_2213_),
    .Y(_2236_)
);

AOI21X1 _8699_ (
    .A(_2233_),
    .B(_2232_),
    .C(_1932_),
    .Y(_2237_)
);

AOI21X1 _8700_ (
    .A(_2226_),
    .B(_2230_),
    .C(\genblk1[2].u_ce.Xin0 [1]),
    .Y(_2238_)
);

OAI21X1 _8701_ (
    .A(_2237_),
    .B(_2238_),
    .C(_2236_),
    .Y(_2239_)
);

AOI21X1 _8702_ (
    .A(_2239_),
    .B(_2235_),
    .C(_1895_),
    .Y(_2240_)
);

OAI21X1 _8703_ (
    .A(_1890__bF$buf3),
    .B(_2240_),
    .C(_2212_),
    .Y(_1747_)
);

OAI21X1 _8704_ (
    .A(_2236_),
    .B(_2238_),
    .C(_2231_),
    .Y(_2241_)
);

MUX2X1 _8705_ (
    .A(\genblk1[2].u_ce.Yin12b [9]),
    .B(\genblk1[2].u_ce.Yin12b [8]),
    .S(1'h0),
    .Y(_2242_)
);

MUX2X1 _8706_ (
    .A(_2242_),
    .B(_2197_),
    .S(1'h1),
    .Y(_2243_)
);

NOR2X1 _8707_ (
    .A(1'h0),
    .B(_1896__bF$buf4),
    .Y(_2244_)
);

NAND2X1 _8708_ (
    .A(_2199_),
    .B(_2244_),
    .Y(_2245_)
);

NAND2X1 _8709_ (
    .A(_1893_),
    .B(_2203_),
    .Y(_2246_)
);

NAND2X1 _8710_ (
    .A(_2246_),
    .B(_2245_),
    .Y(_2247_)
);

AOI21X1 _8711_ (
    .A(1'h0),
    .B(_2243_),
    .C(_2247_),
    .Y(_2248_)
);

NAND2X1 _8712_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin12b [7]),
    .Y(_2249_)
);

OAI21X1 _8713_ (
    .A(1'h0),
    .B(_2066_),
    .C(_2249_),
    .Y(_2250_)
);

MUX2X1 _8714_ (
    .A(_2199_),
    .B(_2250_),
    .S(_1896__bF$buf3),
    .Y(_2251_)
);

NAND2X1 _8715_ (
    .A(1'h0),
    .B(_2251_),
    .Y(_2252_)
);

AOI21X1 _8716_ (
    .A(_2207_),
    .B(_2252_),
    .C(_2224_),
    .Y(_2253_)
);

NOR2X1 _8717_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .B(_2253_),
    .Y(_2254_)
);

NAND2X1 _8718_ (
    .A(_2248_),
    .B(_2254_),
    .Y(_2255_)
);

INVX1 _8719_ (
    .A(_2248_),
    .Y(_2256_)
);

OAI21X1 _8720_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2253_),
    .C(_2256_),
    .Y(_2257_)
);

AOI21X1 _8721_ (
    .A(_2255_),
    .B(_2257_),
    .C(_1948_),
    .Y(_2258_)
);

NAND3X1 _8722_ (
    .A(_1948_),
    .B(_2257_),
    .C(_2255_),
    .Y(_2259_)
);

INVX1 _8723_ (
    .A(_2259_),
    .Y(_2260_)
);

NOR2X1 _8724_ (
    .A(_2258_),
    .B(_2260_),
    .Y(_2261_)
);

NOR2X1 _8725_ (
    .A(_2241_),
    .B(_2261_),
    .Y(_2262_)
);

AOI21X1 _8726_ (
    .A(_2213_),
    .B(_2234_),
    .C(_2237_),
    .Y(_2263_)
);

INVX1 _8727_ (
    .A(_2261_),
    .Y(_2264_)
);

OAI21X1 _8728_ (
    .A(_2263_),
    .B(_2264_),
    .C(_2188_),
    .Y(_2265_)
);

OAI22X1 _8729_ (
    .A(_1865_),
    .B(\genblk1[2].u_ce.Vld_bF$buf0 ),
    .C(_2262_),
    .D(_2265_),
    .Y(_1748_)
);

NAND2X1 _8730_ (
    .A(\genblk1[2].u_ce.Xcalc [3]),
    .B(_1890__bF$buf2),
    .Y(_2266_)
);

AOI21X1 _8731_ (
    .A(_2241_),
    .B(_2259_),
    .C(_2258_),
    .Y(_2267_)
);

NAND2X1 _8732_ (
    .A(1'h0),
    .B(_2152_),
    .Y(_2268_)
);

OAI21X1 _8733_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin12b [9]),
    .C(_2268_),
    .Y(_2269_)
);

NAND2X1 _8734_ (
    .A(_1896__bF$buf2),
    .B(_2220_),
    .Y(_2270_)
);

OAI21X1 _8735_ (
    .A(_1896__bF$buf1),
    .B(_2269_),
    .C(_2270_),
    .Y(_2271_)
);

NAND2X1 _8736_ (
    .A(_2222_),
    .B(_2244_),
    .Y(_2272_)
);

NAND2X1 _8737_ (
    .A(_1893_),
    .B(_2215_),
    .Y(_2273_)
);

NAND2X1 _8738_ (
    .A(_2273_),
    .B(_2272_),
    .Y(_2274_)
);

AOI21X1 _8739_ (
    .A(_2271_),
    .B(1'h0),
    .C(_2274_),
    .Y(_2275_)
);

NAND3X1 _8740_ (
    .A(_2248_),
    .B(_2229_),
    .C(_2208_),
    .Y(_2276_)
);

NAND2X1 _8741_ (
    .A(_1985__bF$buf4),
    .B(_2276_),
    .Y(_2277_)
);

OR2X2 _8742_ (
    .A(_2277_),
    .B(_2275_),
    .Y(_2278_)
);

INVX1 _8743_ (
    .A(_2276_),
    .Y(_2279_)
);

OAI21X1 _8744_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf4 ),
    .B(_2279_),
    .C(_2275_),
    .Y(_2280_)
);

NAND3X1 _8745_ (
    .A(\genblk1[2].u_ce.Xin1 [1]),
    .B(_2280_),
    .C(_2278_),
    .Y(_2281_)
);

INVX1 _8746_ (
    .A(_2275_),
    .Y(_2282_)
);

OR2X2 _8747_ (
    .A(_2277_),
    .B(_2282_),
    .Y(_2283_)
);

OAI21X1 _8748_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2279_),
    .C(_2282_),
    .Y(_2284_)
);

NAND3X1 _8749_ (
    .A(_1927_),
    .B(_2284_),
    .C(_2283_),
    .Y(_2285_)
);

NAND2X1 _8750_ (
    .A(_2281_),
    .B(_2285_),
    .Y(_2286_)
);

OR2X2 _8751_ (
    .A(_2267_),
    .B(_2286_),
    .Y(_2287_)
);

NAND2X1 _8752_ (
    .A(_2286_),
    .B(_2267_),
    .Y(_2288_)
);

AOI21X1 _8753_ (
    .A(_2287_),
    .B(_2288_),
    .C(_1895_),
    .Y(_2289_)
);

OAI21X1 _8754_ (
    .A(_1890__bF$buf1),
    .B(_2289_),
    .C(_2266_),
    .Y(_1749_)
);

OAI21X1 _8755_ (
    .A(_2286_),
    .B(_2267_),
    .C(_2281_),
    .Y(_2290_)
);

NAND2X1 _8756_ (
    .A(1'h0),
    .B(\genblk1[2].u_ce.Yin12b [11]),
    .Y(_2291_)
);

OAI21X1 _8757_ (
    .A(1'h0),
    .B(_2152_),
    .C(_2291_),
    .Y(_2292_)
);

NAND2X1 _8758_ (
    .A(1'h1),
    .B(_2292_),
    .Y(_2293_)
);

OAI21X1 _8759_ (
    .A(1'h1),
    .B(_2242_),
    .C(_2293_),
    .Y(_2294_)
);

NAND2X1 _8760_ (
    .A(1'h0),
    .B(_2294_),
    .Y(_2295_)
);

OAI21X1 _8761_ (
    .A(1'h0),
    .B(_2251_),
    .C(_2295_),
    .Y(_2296_)
);

INVX1 _8762_ (
    .A(_2296_),
    .Y(_2297_)
);

OAI21X1 _8763_ (
    .A(_2282_),
    .B(_2276_),
    .C(_1985__bF$buf3),
    .Y(_2298_)
);

OR2X2 _8764_ (
    .A(_2298_),
    .B(_2297_),
    .Y(_2299_)
);

NAND2X1 _8765_ (
    .A(_2297_),
    .B(_2298_),
    .Y(_2300_)
);

NAND3X1 _8766_ (
    .A(\genblk1[2].u_ce.Xin12b [4]),
    .B(_2300_),
    .C(_2299_),
    .Y(_2301_)
);

OR2X2 _8767_ (
    .A(_2298_),
    .B(_2296_),
    .Y(_2302_)
);

NAND2X1 _8768_ (
    .A(_2296_),
    .B(_2298_),
    .Y(_2303_)
);

NAND3X1 _8769_ (
    .A(_1929_),
    .B(_2303_),
    .C(_2302_),
    .Y(_2304_)
);

AND2X2 _8770_ (
    .A(_2301_),
    .B(_2304_),
    .Y(_2305_)
);

NAND2X1 _8771_ (
    .A(_2305_),
    .B(_2290_),
    .Y(_2306_)
);

INVX1 _8772_ (
    .A(_2258_),
    .Y(_2307_)
);

OAI21X1 _8773_ (
    .A(_2260_),
    .B(_2263_),
    .C(_2307_),
    .Y(_2308_)
);

INVX1 _8774_ (
    .A(_2281_),
    .Y(_2309_)
);

AOI21X1 _8775_ (
    .A(_2308_),
    .B(_2285_),
    .C(_2309_),
    .Y(_2310_)
);

NAND2X1 _8776_ (
    .A(_2304_),
    .B(_2301_),
    .Y(_2311_)
);

NAND2X1 _8777_ (
    .A(_2311_),
    .B(_2310_),
    .Y(_2312_)
);

NAND2X1 _8778_ (
    .A(_2306_),
    .B(_2312_),
    .Y(_2313_)
);

AOI22X1 _8779_ (
    .A(_1867_),
    .B(_1890__bF$buf0),
    .C(_2313_),
    .D(_2188_),
    .Y(_1750_)
);

NAND3X1 _8780_ (
    .A(_2275_),
    .B(_2297_),
    .C(_2279_),
    .Y(_2314_)
);

NOR2X1 _8781_ (
    .A(1'h1),
    .B(_2269_),
    .Y(_2315_)
);

NOR2X1 _8782_ (
    .A(_1896__bF$buf0),
    .B(_2176_),
    .Y(_2316_)
);

OAI21X1 _8783_ (
    .A(_2316_),
    .B(_2315_),
    .C(1'h0),
    .Y(_2317_)
);

OAI21X1 _8784_ (
    .A(1'h0),
    .B(_2223_),
    .C(_2317_),
    .Y(_2318_)
);

NAND3X1 _8785_ (
    .A(_1985__bF$buf2),
    .B(_2318_),
    .C(_2314_),
    .Y(_2319_)
);

INVX1 _8786_ (
    .A(_2318_),
    .Y(_2320_)
);

NAND3X1 _8787_ (
    .A(_2248_),
    .B(_2275_),
    .C(_2253_),
    .Y(_2321_)
);

OAI21X1 _8788_ (
    .A(_2296_),
    .B(_2321_),
    .C(_1985__bF$buf1),
    .Y(_2322_)
);

NAND2X1 _8789_ (
    .A(_2320_),
    .B(_2322_),
    .Y(_2323_)
);

NAND3X1 _8790_ (
    .A(\genblk1[2].u_ce.Xin12b [5]),
    .B(_2323_),
    .C(_2319_),
    .Y(_2324_)
);

NAND3X1 _8791_ (
    .A(_1985__bF$buf0),
    .B(_2320_),
    .C(_2314_),
    .Y(_2325_)
);

NAND2X1 _8792_ (
    .A(_2318_),
    .B(_2322_),
    .Y(_2326_)
);

NAND3X1 _8793_ (
    .A(_1937_),
    .B(_2326_),
    .C(_2325_),
    .Y(_2327_)
);

NAND2X1 _8794_ (
    .A(_2324_),
    .B(_2327_),
    .Y(_2328_)
);

AOI21X1 _8795_ (
    .A(_2306_),
    .B(_2301_),
    .C(_2328_),
    .Y(_2329_)
);

OAI21X1 _8796_ (
    .A(_2311_),
    .B(_2310_),
    .C(_2301_),
    .Y(_2330_)
);

AND2X2 _8797_ (
    .A(_2324_),
    .B(_2327_),
    .Y(_2331_)
);

OAI21X1 _8798_ (
    .A(_2331_),
    .B(_2330_),
    .C(_2188_),
    .Y(_2332_)
);

OAI22X1 _8799_ (
    .A(_1882_),
    .B(\genblk1[2].u_ce.Vld_bF$buf4 ),
    .C(_2329_),
    .D(_2332_),
    .Y(_1751_)
);

NOR2X1 _8800_ (
    .A(_2296_),
    .B(_2321_),
    .Y(_2333_)
);

NAND2X1 _8801_ (
    .A(_2320_),
    .B(_2333_),
    .Y(_2334_)
);

AOI21X1 _8802_ (
    .A(_1896__bF$buf4),
    .B(_2292_),
    .C(_2316_),
    .Y(_2335_)
);

NAND2X1 _8803_ (
    .A(_1923__bF$buf3),
    .B(_2243_),
    .Y(_2336_)
);

OAI21X1 _8804_ (
    .A(_1923__bF$buf2),
    .B(_2335_),
    .C(_2336_),
    .Y(_2337_)
);

NAND3X1 _8805_ (
    .A(_1985__bF$buf5),
    .B(_2337_),
    .C(_2334_),
    .Y(_2338_)
);

NOR3X1 _8806_ (
    .A(_2296_),
    .B(_2318_),
    .C(_2321_),
    .Y(_2339_)
);

INVX1 _8807_ (
    .A(_2337_),
    .Y(_2340_)
);

OAI21X1 _8808_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2339_),
    .C(_2340_),
    .Y(_2341_)
);

NAND3X1 _8809_ (
    .A(\genblk1[2].u_ce.Xin12b [6]),
    .B(_2341_),
    .C(_2338_),
    .Y(_2342_)
);

NAND3X1 _8810_ (
    .A(_1985__bF$buf4),
    .B(_2340_),
    .C(_2334_),
    .Y(_2343_)
);

OAI21X1 _8811_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .B(_2339_),
    .C(_2337_),
    .Y(_2344_)
);

NAND3X1 _8812_ (
    .A(_1939_),
    .B(_2344_),
    .C(_2343_),
    .Y(_2345_)
);

AND2X2 _8813_ (
    .A(_2342_),
    .B(_2345_),
    .Y(_2346_)
);

NAND2X1 _8814_ (
    .A(_2305_),
    .B(_2331_),
    .Y(_2347_)
);

INVX1 _8815_ (
    .A(_2301_),
    .Y(_2348_)
);

INVX1 _8816_ (
    .A(_2324_),
    .Y(_2349_)
);

AOI21X1 _8817_ (
    .A(_2348_),
    .B(_2327_),
    .C(_2349_),
    .Y(_2350_)
);

OAI21X1 _8818_ (
    .A(_2310_),
    .B(_2347_),
    .C(_2350_),
    .Y(_2351_)
);

AND2X2 _8819_ (
    .A(_2351_),
    .B(_2346_),
    .Y(_2352_)
);

NOR2X1 _8820_ (
    .A(_2346_),
    .B(_2351_),
    .Y(_2353_)
);

OAI21X1 _8821_ (
    .A(_2353_),
    .B(_2352_),
    .C(_1894_),
    .Y(_2354_)
);

NAND2X1 _8822_ (
    .A(\genblk1[2].u_ce.Vld_bF$buf3 ),
    .B(_2354_),
    .Y(_2355_)
);

OAI21X1 _8823_ (
    .A(_1868_),
    .B(\genblk1[2].u_ce.Vld_bF$buf2 ),
    .C(_2355_),
    .Y(_1752_)
);

INVX1 _8824_ (
    .A(_2342_),
    .Y(_2356_)
);

NOR2X1 _8825_ (
    .A(_2356_),
    .B(_2352_),
    .Y(_2357_)
);

NAND2X1 _8826_ (
    .A(_2340_),
    .B(_2339_),
    .Y(_2358_)
);

NOR2X1 _8827_ (
    .A(_1923__bF$buf1),
    .B(_2176_),
    .Y(_2359_)
);

AOI21X1 _8828_ (
    .A(_2271_),
    .B(_1923__bF$buf0),
    .C(_2359_),
    .Y(_2360_)
);

NAND3X1 _8829_ (
    .A(_1985__bF$buf3),
    .B(_2360_),
    .C(_2358_),
    .Y(_2361_)
);

INVX1 _8830_ (
    .A(_2361_),
    .Y(_2362_)
);

AOI21X1 _8831_ (
    .A(_2358_),
    .B(_1985__bF$buf2),
    .C(_2360_),
    .Y(_2363_)
);

OAI21X1 _8832_ (
    .A(_2363_),
    .B(_2362_),
    .C(\genblk1[2].u_ce.Xin12b [7]),
    .Y(_2364_)
);

INVX1 _8833_ (
    .A(_2363_),
    .Y(_2365_)
);

NAND3X1 _8834_ (
    .A(_1942_),
    .B(_2361_),
    .C(_2365_),
    .Y(_2366_)
);

AND2X2 _8835_ (
    .A(_2366_),
    .B(_2364_),
    .Y(_2367_)
);

OR2X2 _8836_ (
    .A(_2357_),
    .B(_2367_),
    .Y(_2368_)
);

AOI21X1 _8837_ (
    .A(_2357_),
    .B(_2367_),
    .C(_2187_),
    .Y(_2369_)
);

AOI22X1 _8838_ (
    .A(_1881_),
    .B(_1890__bF$buf4),
    .C(_2368_),
    .D(_2369_),
    .Y(_1753_)
);

NOR2X1 _8839_ (
    .A(_2311_),
    .B(_2328_),
    .Y(_2370_)
);

OAI21X1 _8840_ (
    .A(_2301_),
    .B(_2328_),
    .C(_2324_),
    .Y(_2371_)
);

AOI21X1 _8841_ (
    .A(_2370_),
    .B(_2290_),
    .C(_2371_),
    .Y(_2372_)
);

AOI21X1 _8842_ (
    .A(_2365_),
    .B(_2361_),
    .C(_1942_),
    .Y(_2373_)
);

AOI21X1 _8843_ (
    .A(_2356_),
    .B(_2366_),
    .C(_2373_),
    .Y(_2374_)
);

NAND3X1 _8844_ (
    .A(_2346_),
    .B(_2364_),
    .C(_2366_),
    .Y(_2375_)
);

OAI21X1 _8845_ (
    .A(_2375_),
    .B(_2372_),
    .C(_2374_),
    .Y(_2376_)
);

NAND3X1 _8846_ (
    .A(_2340_),
    .B(_2360_),
    .C(_2339_),
    .Y(_2377_)
);

INVX1 _8847_ (
    .A(_2294_),
    .Y(_2378_)
);

INVX1 _8848_ (
    .A(_2359_),
    .Y(_2379_)
);

OAI21X1 _8849_ (
    .A(1'h0),
    .B(_2378_),
    .C(_2379_),
    .Y(_2380_)
);

INVX1 _8850_ (
    .A(_2380_),
    .Y(_2381_)
);

NAND3X1 _8851_ (
    .A(_1985__bF$buf1),
    .B(_2381_),
    .C(_2377_),
    .Y(_2382_)
);

INVX1 _8852_ (
    .A(_2382_),
    .Y(_2383_)
);

AOI21X1 _8853_ (
    .A(_2377_),
    .B(_1985__bF$buf0),
    .C(_2381_),
    .Y(_2384_)
);

OAI21X1 _8854_ (
    .A(_2384_),
    .B(_2383_),
    .C(\genblk1[2].u_ce.Xin12b [8]),
    .Y(_2385_)
);

INVX1 _8855_ (
    .A(_2384_),
    .Y(_2386_)
);

NAND3X1 _8856_ (
    .A(_1944_),
    .B(_2382_),
    .C(_2386_),
    .Y(_2387_)
);

AND2X2 _8857_ (
    .A(_2387_),
    .B(_2385_),
    .Y(_2388_)
);

OR2X2 _8858_ (
    .A(_2376_),
    .B(_2388_),
    .Y(_2389_)
);

INVX1 _8859_ (
    .A(_2389_),
    .Y(_2390_)
);

NAND2X1 _8860_ (
    .A(_2388_),
    .B(_2376_),
    .Y(_2391_)
);

NAND2X1 _8861_ (
    .A(_2188_),
    .B(_2391_),
    .Y(_2392_)
);

OAI22X1 _8862_ (
    .A(_1870_),
    .B(\genblk1[2].u_ce.Vld_bF$buf1 ),
    .C(_2392_),
    .D(_2390_),
    .Y(_1754_)
);

NOR3X1 _8863_ (
    .A(_2318_),
    .B(_2337_),
    .C(_2314_),
    .Y(_2393_)
);

NAND3X1 _8864_ (
    .A(_2360_),
    .B(_2381_),
    .C(_2393_),
    .Y(_2394_)
);

OR2X2 _8865_ (
    .A(_2315_),
    .B(_2316_),
    .Y(_2395_)
);

AOI21X1 _8866_ (
    .A(_2395_),
    .B(_1923__bF$buf3),
    .C(_2359_),
    .Y(_2396_)
);

INVX1 _8867_ (
    .A(_2396_),
    .Y(_2397_)
);

NAND3X1 _8868_ (
    .A(_1985__bF$buf5),
    .B(_2397_),
    .C(_2394_),
    .Y(_2398_)
);

OAI21X1 _8869_ (
    .A(_2380_),
    .B(_2377_),
    .C(_1985__bF$buf4),
    .Y(_2399_)
);

NAND2X1 _8870_ (
    .A(_2396_),
    .B(_2399_),
    .Y(_2400_)
);

NAND3X1 _8871_ (
    .A(\genblk1[2].u_ce.Xin12b [9]),
    .B(_2400_),
    .C(_2398_),
    .Y(_2401_)
);

NAND3X1 _8872_ (
    .A(_1985__bF$buf3),
    .B(_2396_),
    .C(_2394_),
    .Y(_2402_)
);

NAND2X1 _8873_ (
    .A(_2397_),
    .B(_2399_),
    .Y(_2403_)
);

NAND3X1 _8874_ (
    .A(_1989_),
    .B(_2403_),
    .C(_2402_),
    .Y(_2404_)
);

NAND2X1 _8875_ (
    .A(_2401_),
    .B(_2404_),
    .Y(_2405_)
);

AOI21X1 _8876_ (
    .A(_2391_),
    .B(_2385_),
    .C(_2405_),
    .Y(_2406_)
);

NAND3X1 _8877_ (
    .A(_2385_),
    .B(_2405_),
    .C(_2391_),
    .Y(_2407_)
);

NAND2X1 _8878_ (
    .A(_2188_),
    .B(_2407_),
    .Y(_2408_)
);

OAI22X1 _8879_ (
    .A(_1878_),
    .B(\genblk1[2].u_ce.Vld_bF$buf0 ),
    .C(_2406_),
    .D(_2408_),
    .Y(_1755_)
);

NAND2X1 _8880_ (
    .A(\genblk1[2].u_ce.Xcalc [10]),
    .B(_1890__bF$buf3),
    .Y(_2409_)
);

OAI21X1 _8881_ (
    .A(1'h0),
    .B(_2335_),
    .C(_2379_),
    .Y(_2410_)
);

OAI21X1 _8882_ (
    .A(_2397_),
    .B(_2394_),
    .C(_1985__bF$buf2),
    .Y(_2411_)
);

NOR2X1 _8883_ (
    .A(_2410_),
    .B(_2411_),
    .Y(_2412_)
);

NAND2X1 _8884_ (
    .A(_2410_),
    .B(_2411_),
    .Y(_2413_)
);

INVX1 _8885_ (
    .A(_2413_),
    .Y(_2414_)
);

OAI21X1 _8886_ (
    .A(_2412_),
    .B(_2414_),
    .C(\genblk1[2].u_ce.Xin12b [10]),
    .Y(_2415_)
);

INVX1 _8887_ (
    .A(_2412_),
    .Y(_2416_)
);

NAND3X1 _8888_ (
    .A(_2019_),
    .B(_2413_),
    .C(_2416_),
    .Y(_2417_)
);

AND2X2 _8889_ (
    .A(_2417_),
    .B(_2415_),
    .Y(_2418_)
);

OAI21X1 _8890_ (
    .A(_2385_),
    .B(_2405_),
    .C(_2401_),
    .Y(_2419_)
);

NAND3X1 _8891_ (
    .A(_2346_),
    .B(_2351_),
    .C(_2367_),
    .Y(_2420_)
);

NAND3X1 _8892_ (
    .A(_2401_),
    .B(_2404_),
    .C(_2388_),
    .Y(_2421_)
);

AOI21X1 _8893_ (
    .A(_2420_),
    .B(_2374_),
    .C(_2421_),
    .Y(_2422_)
);

OAI21X1 _8894_ (
    .A(_2419_),
    .B(_2422_),
    .C(_2418_),
    .Y(_2423_)
);

NAND2X1 _8895_ (
    .A(_2415_),
    .B(_2417_),
    .Y(_2424_)
);

NAND2X1 _8896_ (
    .A(_2385_),
    .B(_2387_),
    .Y(_2425_)
);

NOR2X1 _8897_ (
    .A(_2425_),
    .B(_2405_),
    .Y(_2426_)
);

AOI21X1 _8898_ (
    .A(_2376_),
    .B(_2426_),
    .C(_2419_),
    .Y(_2427_)
);

NAND2X1 _8899_ (
    .A(_2424_),
    .B(_2427_),
    .Y(_2428_)
);

AOI21X1 _8900_ (
    .A(_2423_),
    .B(_2428_),
    .C(_1895_),
    .Y(_2429_)
);

OAI21X1 _8901_ (
    .A(_1890__bF$buf2),
    .B(_2429_),
    .C(_2409_),
    .Y(_1756_)
);

NAND2X1 _8902_ (
    .A(\genblk1[2].u_ce.Xcalc [11]),
    .B(_1890__bF$buf1),
    .Y(_2430_)
);

OR2X2 _8903_ (
    .A(_2394_),
    .B(_2397_),
    .Y(_2431_)
);

OAI21X1 _8904_ (
    .A(_2410_),
    .B(_2431_),
    .C(_1985__bF$buf1),
    .Y(_2432_)
);

OR2X2 _8905_ (
    .A(_2432_),
    .B(_2178_),
    .Y(_2433_)
);

NAND2X1 _8906_ (
    .A(_2178_),
    .B(_2432_),
    .Y(_2434_)
);

AOI22X1 _8907_ (
    .A(_2433_),
    .B(_2434_),
    .C(_2423_),
    .D(_2415_),
    .Y(_2435_)
);

OAI21X1 _8908_ (
    .A(_2424_),
    .B(_2427_),
    .C(_2415_),
    .Y(_2436_)
);

NAND2X1 _8909_ (
    .A(_2434_),
    .B(_2433_),
    .Y(_2437_)
);

OAI21X1 _8910_ (
    .A(_2437_),
    .B(_2436_),
    .C(_2188_),
    .Y(_2438_)
);

OAI21X1 _8911_ (
    .A(_2435_),
    .B(_2438_),
    .C(_2430_),
    .Y(_1757_)
);

NAND2X1 _8912_ (
    .A(1'h0),
    .B(1'h1),
    .Y(_2439_)
);

OAI21X1 _8913_ (
    .A(_1923__bF$buf2),
    .B(_2105_),
    .C(_2439_),
    .Y(_2440_)
);

NOR2X1 _8914_ (
    .A(_1886_),
    .B(_2440_),
    .Y(_2441_)
);

AND2X2 _8915_ (
    .A(_2440_),
    .B(_1886_),
    .Y(_2442_)
);

OR2X2 _8916_ (
    .A(_2442_),
    .B(_2441_),
    .Y(_2443_)
);

NAND2X1 _8917_ (
    .A(\genblk1[2].u_ce.Acalc [0]),
    .B(_1890__bF$buf0),
    .Y(_2444_)
);

OAI21X1 _8918_ (
    .A(_1890__bF$buf4),
    .B(_2443_),
    .C(_2444_),
    .Y(_1758_)
);

NAND2X1 _8919_ (
    .A(\genblk1[2].u_ce.Acalc [1]),
    .B(_1890__bF$buf3),
    .Y(_2445_)
);

OAI21X1 _8920_ (
    .A(1'h1),
    .B(_1892_),
    .C(1'h0),
    .Y(_2446_)
);

OAI21X1 _8921_ (
    .A(1'h0),
    .B(_1892_),
    .C(_2446_),
    .Y(_2447_)
);

OAI21X1 _8922_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2440_),
    .C(_2447_),
    .Y(_2448_)
);

OAI21X1 _8923_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf4 ),
    .B(_2447_),
    .C(_2448_),
    .Y(_2449_)
);

OR2X2 _8924_ (
    .A(_2449_),
    .B(\genblk1[2].u_ce.Ain0 [1]),
    .Y(_2450_)
);

NAND2X1 _8925_ (
    .A(\genblk1[2].u_ce.Ain0 [1]),
    .B(_2449_),
    .Y(_2451_)
);

NAND2X1 _8926_ (
    .A(_2451_),
    .B(_2450_),
    .Y(_2452_)
);

NOR2X1 _8927_ (
    .A(_2441_),
    .B(_2452_),
    .Y(_2453_)
);

NAND2X1 _8928_ (
    .A(_2441_),
    .B(_2452_),
    .Y(_2454_)
);

NAND2X1 _8929_ (
    .A(\genblk1[2].u_ce.Vld_bF$buf4 ),
    .B(_2454_),
    .Y(_2455_)
);

OAI21X1 _8930_ (
    .A(_2453_),
    .B(_2455_),
    .C(_2445_),
    .Y(_1759_)
);

NAND2X1 _8931_ (
    .A(\genblk1[2].u_ce.Acalc [2]),
    .B(_1890__bF$buf2),
    .Y(_2456_)
);

OAI21X1 _8932_ (
    .A(_1888_),
    .B(_2449_),
    .C(_2454_),
    .Y(_2457_)
);

OAI21X1 _8933_ (
    .A(_1892_),
    .B(_1896__bF$buf3),
    .C(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .Y(_2458_)
);

NAND3X1 _8934_ (
    .A(1'h0),
    .B(_2105_),
    .C(_2458_),
    .Y(_2459_)
);

OAI21X1 _8935_ (
    .A(1'h0),
    .B(_2458_),
    .C(_2459_),
    .Y(_2460_)
);

NAND2X1 _8936_ (
    .A(\genblk1[2].u_ce.Ain1 [0]),
    .B(_2460_),
    .Y(_2461_)
);

OR2X2 _8937_ (
    .A(_2460_),
    .B(\genblk1[2].u_ce.Ain1 [0]),
    .Y(_2462_)
);

NAND2X1 _8938_ (
    .A(_2461_),
    .B(_2462_),
    .Y(_2463_)
);

INVX1 _8939_ (
    .A(_2463_),
    .Y(_2464_)
);

NOR2X1 _8940_ (
    .A(_2464_),
    .B(_2457_),
    .Y(_2465_)
);

NAND2X1 _8941_ (
    .A(_2464_),
    .B(_2457_),
    .Y(_2466_)
);

NAND2X1 _8942_ (
    .A(\genblk1[2].u_ce.Vld_bF$buf3 ),
    .B(_2466_),
    .Y(_2467_)
);

OAI21X1 _8943_ (
    .A(_2465_),
    .B(_2467_),
    .C(_2456_),
    .Y(_1760_)
);

NAND2X1 _8944_ (
    .A(_2461_),
    .B(_2466_),
    .Y(_2468_)
);

INVX1 _8945_ (
    .A(_2468_),
    .Y(_2469_)
);

INVX1 _8946_ (
    .A(\genblk1[2].u_ce.Ain1 [1]),
    .Y(_2470_)
);

OAI21X1 _8947_ (
    .A(1'h0),
    .B(_1896__bF$buf2),
    .C(1'h0),
    .Y(_2471_)
);

NAND2X1 _8948_ (
    .A(_1985__bF$buf0),
    .B(_2471_),
    .Y(_2472_)
);

OAI21X1 _8949_ (
    .A(1'h0),
    .B(1'h1),
    .C(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .Y(_2473_)
);

OAI21X1 _8950_ (
    .A(_1892_),
    .B(_2473_),
    .C(_2472_),
    .Y(_2474_)
);

NOR2X1 _8951_ (
    .A(_2470_),
    .B(_2474_),
    .Y(_2475_)
);

NAND2X1 _8952_ (
    .A(_2470_),
    .B(_2474_),
    .Y(_2476_)
);

INVX1 _8953_ (
    .A(_2476_),
    .Y(_2477_)
);

OAI21X1 _8954_ (
    .A(_2475_),
    .B(_2477_),
    .C(_2469_),
    .Y(_2478_)
);

INVX1 _8955_ (
    .A(_2475_),
    .Y(_2479_)
);

NAND3X1 _8956_ (
    .A(_2479_),
    .B(_2476_),
    .C(_2468_),
    .Y(_2480_)
);

NAND2X1 _8957_ (
    .A(_2480_),
    .B(_2478_),
    .Y(_2481_)
);

NAND2X1 _8958_ (
    .A(\genblk1[2].u_ce.Acalc [3]),
    .B(_1890__bF$buf1),
    .Y(_2482_)
);

OAI21X1 _8959_ (
    .A(_1890__bF$buf0),
    .B(_2481_),
    .C(_2482_),
    .Y(_1761_)
);

NOR2X1 _8960_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf1 ),
    .B(_2447_),
    .Y(_2483_)
);

NAND3X1 _8961_ (
    .A(1'h0),
    .B(_1923__bF$buf1),
    .C(_1896__bF$buf1),
    .Y(_2484_)
);

AOI21X1 _8962_ (
    .A(_2446_),
    .B(_2484_),
    .C(_1985__bF$buf5),
    .Y(_2485_)
);

NOR2X1 _8963_ (
    .A(_2485_),
    .B(_2483_),
    .Y(_2486_)
);

NAND2X1 _8964_ (
    .A(\genblk1[2].u_ce.Ain12b [4]),
    .B(_2486_),
    .Y(_2487_)
);

INVX1 _8965_ (
    .A(\genblk1[2].u_ce.Ain12b [4]),
    .Y(_2488_)
);

OAI21X1 _8966_ (
    .A(_2485_),
    .B(_2483_),
    .C(_2488_),
    .Y(_2489_)
);

NAND2X1 _8967_ (
    .A(_2489_),
    .B(_2487_),
    .Y(_2490_)
);

AOI21X1 _8968_ (
    .A(_2468_),
    .B(_2476_),
    .C(_2475_),
    .Y(_2491_)
);

AND2X2 _8969_ (
    .A(_2491_),
    .B(_2490_),
    .Y(_2492_)
);

OAI21X1 _8970_ (
    .A(_2490_),
    .B(_2491_),
    .C(\genblk1[2].u_ce.Vld_bF$buf2 ),
    .Y(_2493_)
);

OAI22X1 _8971_ (
    .A(_1829_),
    .B(\genblk1[2].u_ce.Vld_bF$buf1 ),
    .C(_2493_),
    .D(_2492_),
    .Y(_1762_)
);

NAND2X1 _8972_ (
    .A(\genblk1[2].u_ce.Acalc [5]),
    .B(_1890__bF$buf4),
    .Y(_2494_)
);

OAI21X1 _8973_ (
    .A(_2490_),
    .B(_2491_),
    .C(_2487_),
    .Y(_2495_)
);

OAI21X1 _8974_ (
    .A(1'h0),
    .B(1'h1),
    .C(_1924_),
    .Y(_2496_)
);

NAND2X1 _8975_ (
    .A(_1985__bF$buf4),
    .B(_2496_),
    .Y(_2497_)
);

INVX1 _8976_ (
    .A(_2497_),
    .Y(_2498_)
);

NOR2X1 _8977_ (
    .A(_1985__bF$buf3),
    .B(_2496_),
    .Y(_2499_)
);

NOR2X1 _8978_ (
    .A(_2499_),
    .B(_2498_),
    .Y(_2500_)
);

NAND2X1 _8979_ (
    .A(\genblk1[2].u_ce.Ain12b [5]),
    .B(_2500_),
    .Y(_2501_)
);

INVX1 _8980_ (
    .A(\genblk1[2].u_ce.Ain12b [5]),
    .Y(_2502_)
);

OAI21X1 _8981_ (
    .A(_2499_),
    .B(_2498_),
    .C(_2502_),
    .Y(_2503_)
);

NAND2X1 _8982_ (
    .A(_2503_),
    .B(_2501_),
    .Y(_2504_)
);

INVX1 _8983_ (
    .A(_2504_),
    .Y(_2505_)
);

NOR2X1 _8984_ (
    .A(_2505_),
    .B(_2495_),
    .Y(_2506_)
);

NAND2X1 _8985_ (
    .A(_2505_),
    .B(_2495_),
    .Y(_2507_)
);

NAND2X1 _8986_ (
    .A(\genblk1[2].u_ce.Vld_bF$buf0 ),
    .B(_2507_),
    .Y(_2508_)
);

OAI21X1 _8987_ (
    .A(_2506_),
    .B(_2508_),
    .C(_2494_),
    .Y(_1763_)
);

NAND2X1 _8988_ (
    .A(\genblk1[2].u_ce.Acalc [6]),
    .B(_1890__bF$buf3),
    .Y(_2509_)
);

INVX1 _8989_ (
    .A(_2491_),
    .Y(_2510_)
);

NOR2X1 _8990_ (
    .A(_2490_),
    .B(_2504_),
    .Y(_2511_)
);

OAI21X1 _8991_ (
    .A(_2487_),
    .B(_2504_),
    .C(_2501_),
    .Y(_2512_)
);

AOI21X1 _8992_ (
    .A(_2510_),
    .B(_2511_),
    .C(_2512_),
    .Y(_2513_)
);

OAI21X1 _8993_ (
    .A(1'h0),
    .B(_2439_),
    .C(_1894_),
    .Y(_2514_)
);

NOR2X1 _8994_ (
    .A(_1985__bF$buf2),
    .B(_2514_),
    .Y(_2515_)
);

NAND2X1 _8995_ (
    .A(_1985__bF$buf1),
    .B(_2514_),
    .Y(_2516_)
);

INVX1 _8996_ (
    .A(_2516_),
    .Y(_2517_)
);

NOR2X1 _8997_ (
    .A(_2515_),
    .B(_2517_),
    .Y(_2518_)
);

NAND2X1 _8998_ (
    .A(\genblk1[2].u_ce.Ain12b [6]),
    .B(_2518_),
    .Y(_2519_)
);

OR2X2 _8999_ (
    .A(_2518_),
    .B(\genblk1[2].u_ce.Ain12b [6]),
    .Y(_2520_)
);

AND2X2 _9000_ (
    .A(_2520_),
    .B(_2519_),
    .Y(_2521_)
);

INVX1 _9001_ (
    .A(_2521_),
    .Y(_2522_)
);

AND2X2 _9002_ (
    .A(_2513_),
    .B(_2522_),
    .Y(_2523_)
);

OAI21X1 _9003_ (
    .A(_2522_),
    .B(_2513_),
    .C(\genblk1[2].u_ce.Vld_bF$buf4 ),
    .Y(_2524_)
);

OAI21X1 _9004_ (
    .A(_2524_),
    .B(_2523_),
    .C(_2509_),
    .Y(_1764_)
);

OAI21X1 _9005_ (
    .A(_2522_),
    .B(_2513_),
    .C(_2519_),
    .Y(_2525_)
);

OAI21X1 _9006_ (
    .A(1'h0),
    .B(1'h0),
    .C(\genblk1[2].u_ce.Ain12b_11_bF$buf0 ),
    .Y(_2526_)
);

NAND2X1 _9007_ (
    .A(_2526_),
    .B(_1986_),
    .Y(_2527_)
);

INVX1 _9008_ (
    .A(_2527_),
    .Y(_2528_)
);

NAND2X1 _9009_ (
    .A(\genblk1[2].u_ce.Ain12b [7]),
    .B(_2528_),
    .Y(_2529_)
);

INVX1 _9010_ (
    .A(_2529_),
    .Y(_2530_)
);

NOR2X1 _9011_ (
    .A(\genblk1[2].u_ce.Ain12b [7]),
    .B(_2528_),
    .Y(_2531_)
);

NOR2X1 _9012_ (
    .A(_2531_),
    .B(_2530_),
    .Y(_2532_)
);

INVX1 _9013_ (
    .A(_2532_),
    .Y(_2533_)
);

OR2X2 _9014_ (
    .A(_2525_),
    .B(_2533_),
    .Y(_2534_)
);

AOI21X1 _9015_ (
    .A(_2525_),
    .B(_2533_),
    .C(_1890__bF$buf2),
    .Y(_2535_)
);

AOI22X1 _9016_ (
    .A(_1843_),
    .B(_1890__bF$buf1),
    .C(_2534_),
    .D(_2535_),
    .Y(_1765_)
);

NAND2X1 _9017_ (
    .A(\genblk1[2].u_ce.Acalc [8]),
    .B(_1890__bF$buf0),
    .Y(_2536_)
);

OAI21X1 _9018_ (
    .A(_2531_),
    .B(_2519_),
    .C(_2529_),
    .Y(_2537_)
);

NAND2X1 _9019_ (
    .A(_2532_),
    .B(_2521_),
    .Y(_2538_)
);

INVX1 _9020_ (
    .A(_2538_),
    .Y(_2539_)
);

AOI21X1 _9021_ (
    .A(_2539_),
    .B(_2512_),
    .C(_2537_),
    .Y(_2540_)
);

NAND2X1 _9022_ (
    .A(_2511_),
    .B(_2539_),
    .Y(_2541_)
);

OAI21X1 _9023_ (
    .A(_2541_),
    .B(_2491_),
    .C(_2540_),
    .Y(_2542_)
);

INVX1 _9024_ (
    .A(\genblk1[2].u_ce.Ain12b [8]),
    .Y(_2543_)
);

NAND2X1 _9025_ (
    .A(_1985__bF$buf0),
    .B(_1893_),
    .Y(_2544_)
);

NAND2X1 _9026_ (
    .A(_2473_),
    .B(_2544_),
    .Y(_2545_)
);

OR2X2 _9027_ (
    .A(_2545_),
    .B(_2543_),
    .Y(_2546_)
);

NAND2X1 _9028_ (
    .A(_2543_),
    .B(_2545_),
    .Y(_2547_)
);

AND2X2 _9029_ (
    .A(_2546_),
    .B(_2547_),
    .Y(_2548_)
);

NOR2X1 _9030_ (
    .A(_2548_),
    .B(_2542_),
    .Y(_2549_)
);

NAND2X1 _9031_ (
    .A(_2548_),
    .B(_2542_),
    .Y(_2550_)
);

NAND2X1 _9032_ (
    .A(\genblk1[2].u_ce.Vld_bF$buf3 ),
    .B(_2550_),
    .Y(_2551_)
);

OAI21X1 _9033_ (
    .A(_2549_),
    .B(_2551_),
    .C(_2536_),
    .Y(_1766_)
);

NAND2X1 _9034_ (
    .A(\genblk1[2].u_ce.Acalc [9]),
    .B(_1890__bF$buf4),
    .Y(_2552_)
);

OAI21X1 _9035_ (
    .A(_2543_),
    .B(_2545_),
    .C(_2550_),
    .Y(_2553_)
);

INVX1 _9036_ (
    .A(\genblk1[2].u_ce.Ain12b [9]),
    .Y(_2554_)
);

NAND2X1 _9037_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf4 ),
    .B(_2554_),
    .Y(_2555_)
);

NOR2X1 _9038_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2554_),
    .Y(_2556_)
);

INVX1 _9039_ (
    .A(_2556_),
    .Y(_2557_)
);

NAND2X1 _9040_ (
    .A(_2555_),
    .B(_2557_),
    .Y(_2558_)
);

INVX1 _9041_ (
    .A(_2558_),
    .Y(_2559_)
);

NOR2X1 _9042_ (
    .A(_2559_),
    .B(_2553_),
    .Y(_2560_)
);

NAND2X1 _9043_ (
    .A(_2559_),
    .B(_2553_),
    .Y(_2561_)
);

NAND2X1 _9044_ (
    .A(\genblk1[2].u_ce.Vld_bF$buf2 ),
    .B(_2561_),
    .Y(_2562_)
);

OAI21X1 _9045_ (
    .A(_2560_),
    .B(_2562_),
    .C(_2552_),
    .Y(_1767_)
);

AOI21X1 _9046_ (
    .A(_2553_),
    .B(_2555_),
    .C(_2556_),
    .Y(_2563_)
);

INVX1 _9047_ (
    .A(\genblk1[2].u_ce.Ain12b [10]),
    .Y(_2564_)
);

NAND2X1 _9048_ (
    .A(\genblk1[2].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2564_),
    .Y(_2565_)
);

NAND2X1 _9049_ (
    .A(\genblk1[2].u_ce.Ain12b [10]),
    .B(_1985__bF$buf5),
    .Y(_2566_)
);

NAND2X1 _9050_ (
    .A(_2565_),
    .B(_2566_),
    .Y(_2567_)
);

AND2X2 _9051_ (
    .A(_2563_),
    .B(_2567_),
    .Y(_2568_)
);

OAI21X1 _9052_ (
    .A(_2567_),
    .B(_2563_),
    .C(\genblk1[2].u_ce.Vld_bF$buf1 ),
    .Y(_2569_)
);

OAI22X1 _9053_ (
    .A(_1825_),
    .B(\genblk1[2].u_ce.Vld_bF$buf0 ),
    .C(_2569_),
    .D(_2568_),
    .Y(_1768_)
);

NAND2X1 _9054_ (
    .A(\genblk1[2].u_ce.Acalc [11]),
    .B(_1890__bF$buf3),
    .Y(_2570_)
);

OAI21X1 _9055_ (
    .A(_2567_),
    .B(_2563_),
    .C(_2566_),
    .Y(_2571_)
);

OAI21X1 _9056_ (
    .A(_1890__bF$buf2),
    .B(_2571_),
    .C(_2570_),
    .Y(_1769_)
);

INVX1 _9057_ (
    .A(_1824_),
    .Y(_2572_)
);

NAND3X1 _9058_ (
    .A(_1877_),
    .B(\genblk1[2].u_ce.LoadCtl [5]),
    .C(_1835_),
    .Y(_2573_)
);

NOR2X1 _9059_ (
    .A(_2572_),
    .B(_2573_),
    .Y(_2574_)
);

NAND2X1 _9060_ (
    .A(\genblk1[1].u_ce.X_ [0]),
    .B(_2574_),
    .Y(_2575_)
);

OAI21X1 _9061_ (
    .A(_2019_),
    .B(_2574_),
    .C(_2575_),
    .Y(_1770_)
);

NAND2X1 _9062_ (
    .A(\genblk1[1].u_ce.X_ [1]),
    .B(_2574_),
    .Y(_2576_)
);

OAI21X1 _9063_ (
    .A(_2044_),
    .B(_2574_),
    .C(_2576_),
    .Y(_1771_)
);

INVX1 _9064_ (
    .A(\genblk1[1].u_ce.X_ [0]),
    .Y(_2577_)
);

NAND3X1 _9065_ (
    .A(\genblk1[2].u_ce.LoadCtl [4]),
    .B(_1824_),
    .C(_1835_),
    .Y(_2578_)
);

NAND2X1 _9066_ (
    .A(\genblk1[2].u_ce.Xin12b [8]),
    .B(_2578_),
    .Y(_2579_)
);

OAI21X1 _9067_ (
    .A(_2577_),
    .B(_2578_),
    .C(_2579_),
    .Y(_1772_)
);

INVX1 _9068_ (
    .A(\genblk1[1].u_ce.X_ [1]),
    .Y(_2580_)
);

NAND2X1 _9069_ (
    .A(\genblk1[2].u_ce.Xin12b [9]),
    .B(_2578_),
    .Y(_2581_)
);

OAI21X1 _9070_ (
    .A(_2580_),
    .B(_2578_),
    .C(_2581_),
    .Y(_1773_)
);

NAND2X1 _9071_ (
    .A(_1835_),
    .B(_1831_),
    .Y(_2582_)
);

OAI21X1 _9072_ (
    .A(_1836_),
    .B(_1844_),
    .C(\genblk1[2].u_ce.Xin12b [6]),
    .Y(_2583_)
);

OAI21X1 _9073_ (
    .A(_2577_),
    .B(_2582_),
    .C(_2583_),
    .Y(_1774_)
);

OAI21X1 _9074_ (
    .A(_1836_),
    .B(_1844_),
    .C(\genblk1[2].u_ce.Xin12b [7]),
    .Y(_2584_)
);

OAI21X1 _9075_ (
    .A(_2580_),
    .B(_2582_),
    .C(_2584_),
    .Y(_1775_)
);

NOR2X1 _9076_ (
    .A(_1828_),
    .B(_1836_),
    .Y(_2585_)
);

NAND2X1 _9077_ (
    .A(\genblk1[1].u_ce.X_ [0]),
    .B(_2585_),
    .Y(_2586_)
);

OAI21X1 _9078_ (
    .A(_1929_),
    .B(_2585_),
    .C(_2586_),
    .Y(_1776_)
);

NAND2X1 _9079_ (
    .A(\genblk1[1].u_ce.X_ [1]),
    .B(_2585_),
    .Y(_2587_)
);

OAI21X1 _9080_ (
    .A(_1937_),
    .B(_2585_),
    .C(_2587_),
    .Y(_1777_)
);

OAI21X1 _9081_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_1837_),
    .C(\genblk1[2].u_ce.Xin1 [0]),
    .Y(_2588_)
);

OAI21X1 _9082_ (
    .A(_2577_),
    .B(_1866_),
    .C(_2588_),
    .Y(_1778_)
);

OAI21X1 _9083_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_1837_),
    .C(\genblk1[2].u_ce.Xin1 [1]),
    .Y(_2589_)
);

OAI21X1 _9084_ (
    .A(_2580_),
    .B(_1866_),
    .C(_2589_),
    .Y(_1779_)
);

NAND2X1 _9085_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[1].u_ce.X_ [0]),
    .Y(_2590_)
);

OAI21X1 _9086_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_1952_),
    .C(_2590_),
    .Y(_1780_)
);

NAND2X1 _9087_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[1].u_ce.X_ [1]),
    .Y(_2591_)
);

OAI21X1 _9088_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 ),
    .B(_1932_),
    .C(_2591_),
    .Y(_1781_)
);

NAND2X1 _9089_ (
    .A(\genblk1[1].u_ce.Y_ [0]),
    .B(_2574_),
    .Y(_2592_)
);

OAI21X1 _9090_ (
    .A(_2152_),
    .B(_2574_),
    .C(_2592_),
    .Y(_1782_)
);

NAND2X1 _9091_ (
    .A(\genblk1[1].u_ce.Y_ [1]),
    .B(_2574_),
    .Y(_2593_)
);

OAI21X1 _9092_ (
    .A(_2176_),
    .B(_2574_),
    .C(_2593_),
    .Y(_1783_)
);

INVX1 _9093_ (
    .A(\genblk1[1].u_ce.Y_ [0]),
    .Y(_2594_)
);

NAND2X1 _9094_ (
    .A(\genblk1[2].u_ce.Yin12b [8]),
    .B(_2578_),
    .Y(_2595_)
);

OAI21X1 _9095_ (
    .A(_2594_),
    .B(_2578_),
    .C(_2595_),
    .Y(_1784_)
);

INVX1 _9096_ (
    .A(\genblk1[1].u_ce.Y_ [1]),
    .Y(_2596_)
);

NAND2X1 _9097_ (
    .A(\genblk1[2].u_ce.Yin12b [9]),
    .B(_2578_),
    .Y(_2597_)
);

OAI21X1 _9098_ (
    .A(_2596_),
    .B(_2578_),
    .C(_2597_),
    .Y(_1785_)
);

OAI21X1 _9099_ (
    .A(_1836_),
    .B(_1844_),
    .C(\genblk1[2].u_ce.Yin12b [6]),
    .Y(_1804_)
);

OAI21X1 _9100_ (
    .A(_2594_),
    .B(_2582_),
    .C(_1804_),
    .Y(_1786_)
);

OAI21X1 _9101_ (
    .A(_1836_),
    .B(_1844_),
    .C(\genblk1[2].u_ce.Yin12b [7]),
    .Y(_1805_)
);

OAI21X1 _9102_ (
    .A(_2596_),
    .B(_2582_),
    .C(_1805_),
    .Y(_1787_)
);

NAND2X1 _9103_ (
    .A(\genblk1[1].u_ce.Y_ [0]),
    .B(_2585_),
    .Y(_1806_)
);

OAI21X1 _9104_ (
    .A(_2017_),
    .B(_2585_),
    .C(_1806_),
    .Y(_1788_)
);

NAND2X1 _9105_ (
    .A(\genblk1[1].u_ce.Y_ [1]),
    .B(_2585_),
    .Y(_1807_)
);

OAI21X1 _9106_ (
    .A(_2042_),
    .B(_2585_),
    .C(_1807_),
    .Y(_1789_)
);

OAI21X1 _9107_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_1837_),
    .C(\genblk1[2].u_ce.Yin1 [0]),
    .Y(_1808_)
);

OAI21X1 _9108_ (
    .A(_2594_),
    .B(_1866_),
    .C(_1808_),
    .Y(_1790_)
);

OAI21X1 _9109_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_1837_),
    .C(\genblk1[2].u_ce.Yin1 [1]),
    .Y(_1809_)
);

OAI21X1 _9110_ (
    .A(_2596_),
    .B(_1866_),
    .C(_1809_),
    .Y(_1791_)
);

NAND2X1 _9111_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[1].u_ce.Y_ [0]),
    .Y(_1810_)
);

OAI21X1 _9112_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_2189_),
    .C(_1810_),
    .Y(_1792_)
);

NAND2X1 _9113_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[1].u_ce.Y_ [1]),
    .Y(_1811_)
);

OAI21X1 _9114_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf1 ),
    .B(_1974_),
    .C(_1811_),
    .Y(_1793_)
);

NAND2X1 _9115_ (
    .A(\a[2] [0]),
    .B(_2574_),
    .Y(_1812_)
);

OAI21X1 _9116_ (
    .A(_2564_),
    .B(_2574_),
    .C(_1812_),
    .Y(_1794_)
);

NAND2X1 _9117_ (
    .A(\a[2] [1]),
    .B(_2574_),
    .Y(_1813_)
);

OAI21X1 _9118_ (
    .A(_1985__bF$buf4),
    .B(_2574_),
    .C(_1813_),
    .Y(_1795_)
);

INVX1 _9119_ (
    .A(\a[2] [0]),
    .Y(_1814_)
);

NAND2X1 _9120_ (
    .A(\genblk1[2].u_ce.Ain12b [8]),
    .B(_2578_),
    .Y(_1815_)
);

OAI21X1 _9121_ (
    .A(_1814_),
    .B(_2578_),
    .C(_1815_),
    .Y(_1796_)
);

INVX1 _9122_ (
    .A(\a[2] [1]),
    .Y(_1816_)
);

NAND2X1 _9123_ (
    .A(\genblk1[2].u_ce.Ain12b [9]),
    .B(_2578_),
    .Y(_1817_)
);

OAI21X1 _9124_ (
    .A(_1816_),
    .B(_2578_),
    .C(_1817_),
    .Y(_1797_)
);

OAI21X1 _9125_ (
    .A(_1836_),
    .B(_1844_),
    .C(\genblk1[2].u_ce.Ain12b [6]),
    .Y(_1818_)
);

OAI21X1 _9126_ (
    .A(_1814_),
    .B(_2582_),
    .C(_1818_),
    .Y(_1798_)
);

OAI21X1 _9127_ (
    .A(_1836_),
    .B(_1844_),
    .C(\genblk1[2].u_ce.Ain12b [7]),
    .Y(_1819_)
);

OAI21X1 _9128_ (
    .A(_1816_),
    .B(_2582_),
    .C(_1819_),
    .Y(_1799_)
);

NAND2X1 _9129_ (
    .A(\a[2] [0]),
    .B(_2585_),
    .Y(_1820_)
);

OAI21X1 _9130_ (
    .A(_2488_),
    .B(_2585_),
    .C(_1820_),
    .Y(_1800_)
);

NAND2X1 _9131_ (
    .A(\a[2] [1]),
    .B(_2585_),
    .Y(_1821_)
);

OAI21X1 _9132_ (
    .A(_2502_),
    .B(_2585_),
    .C(_1821_),
    .Y(_1801_)
);

OAI21X1 _9133_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_1837_),
    .C(\genblk1[2].u_ce.Ain1 [0]),
    .Y(_1822_)
);

OAI21X1 _9134_ (
    .A(_1814_),
    .B(_1866_),
    .C(_1822_),
    .Y(_1802_)
);

OAI21X1 _9135_ (
    .A(\genblk1[2].u_ce.LoadCtl_0_bF$buf4 ),
    .B(_1837_),
    .C(\genblk1[2].u_ce.Ain1 [1]),
    .Y(_1823_)
);

OAI21X1 _9136_ (
    .A(_1816_),
    .B(_1866_),
    .C(_1823_),
    .Y(_1803_)
);

DFFPOSX1 _9137_ (
    .CLK(clk_bF$buf19),
    .D(_1732_),
    .Q(\genblk1[2].u_ce.Ain0 [0])
);

DFFPOSX1 _9138_ (
    .CLK(clk_bF$buf18),
    .D(_1733_),
    .Q(\genblk1[2].u_ce.Ain0 [1])
);

DFFPOSX1 _9139_ (
    .CLK(clk_bF$buf17),
    .D(_1734_),
    .Q(\genblk1[2].u_ce.Ycalc [2])
);

DFFPOSX1 _9140_ (
    .CLK(clk_bF$buf16),
    .D(_1735_),
    .Q(\genblk1[2].u_ce.Ycalc [3])
);

DFFPOSX1 _9141_ (
    .CLK(clk_bF$buf15),
    .D(_1736_),
    .Q(\genblk1[2].u_ce.Ycalc [4])
);

DFFPOSX1 _9142_ (
    .CLK(clk_bF$buf14),
    .D(_1737_),
    .Q(\genblk1[2].u_ce.Ycalc [5])
);

DFFPOSX1 _9143_ (
    .CLK(clk_bF$buf13),
    .D(_1738_),
    .Q(\genblk1[2].u_ce.Ycalc [6])
);

DFFPOSX1 _9144_ (
    .CLK(clk_bF$buf12),
    .D(_1739_),
    .Q(\genblk1[2].u_ce.Ycalc [7])
);

DFFPOSX1 _9145_ (
    .CLK(clk_bF$buf11),
    .D(_1740_),
    .Q(\genblk1[2].u_ce.Ycalc [8])
);

DFFPOSX1 _9146_ (
    .CLK(clk_bF$buf10),
    .D(_1741_),
    .Q(\genblk1[2].u_ce.Ycalc [9])
);

DFFPOSX1 _9147_ (
    .CLK(clk_bF$buf9),
    .D(_1742_),
    .Q(\genblk1[2].u_ce.Ycalc [10])
);

DFFPOSX1 _9148_ (
    .CLK(clk_bF$buf8),
    .D(_1743_),
    .Q(\genblk1[2].u_ce.Ycalc [11])
);

DFFPOSX1 _9149_ (
    .CLK(clk_bF$buf7),
    .D(_1744_),
    .Q(\genblk1[2].u_ce.Ycalc [0])
);

DFFPOSX1 _9150_ (
    .CLK(clk_bF$buf6),
    .D(_1745_),
    .Q(\genblk1[2].u_ce.Ycalc [1])
);

DFFPOSX1 _9151_ (
    .CLK(clk_bF$buf5),
    .D(_1746_),
    .Q(\genblk1[2].u_ce.Xcalc [0])
);

DFFPOSX1 _9152_ (
    .CLK(clk_bF$buf4),
    .D(_1747_),
    .Q(\genblk1[2].u_ce.Xcalc [1])
);

DFFPOSX1 _9153_ (
    .CLK(clk_bF$buf3),
    .D(_1748_),
    .Q(\genblk1[2].u_ce.Xcalc [2])
);

DFFPOSX1 _9154_ (
    .CLK(clk_bF$buf2),
    .D(_1749_),
    .Q(\genblk1[2].u_ce.Xcalc [3])
);

DFFPOSX1 _9155_ (
    .CLK(clk_bF$buf1),
    .D(_1750_),
    .Q(\genblk1[2].u_ce.Xcalc [4])
);

DFFPOSX1 _9156_ (
    .CLK(clk_bF$buf0),
    .D(_1751_),
    .Q(\genblk1[2].u_ce.Xcalc [5])
);

DFFPOSX1 _9157_ (
    .CLK(clk_bF$buf75),
    .D(_1752_),
    .Q(\genblk1[2].u_ce.Xcalc [6])
);

DFFPOSX1 _9158_ (
    .CLK(clk_bF$buf74),
    .D(_1753_),
    .Q(\genblk1[2].u_ce.Xcalc [7])
);

DFFPOSX1 _9159_ (
    .CLK(clk_bF$buf73),
    .D(_1754_),
    .Q(\genblk1[2].u_ce.Xcalc [8])
);

DFFPOSX1 _9160_ (
    .CLK(clk_bF$buf72),
    .D(_1755_),
    .Q(\genblk1[2].u_ce.Xcalc [9])
);

DFFPOSX1 _9161_ (
    .CLK(clk_bF$buf71),
    .D(_1756_),
    .Q(\genblk1[2].u_ce.Xcalc [10])
);

DFFPOSX1 _9162_ (
    .CLK(clk_bF$buf70),
    .D(_1757_),
    .Q(\genblk1[2].u_ce.Xcalc [11])
);

DFFPOSX1 _9163_ (
    .CLK(clk_bF$buf69),
    .D(_1758_),
    .Q(\genblk1[2].u_ce.Acalc [0])
);

DFFPOSX1 _9164_ (
    .CLK(clk_bF$buf68),
    .D(_1759_),
    .Q(\genblk1[2].u_ce.Acalc [1])
);

DFFPOSX1 _9165_ (
    .CLK(clk_bF$buf67),
    .D(_1760_),
    .Q(\genblk1[2].u_ce.Acalc [2])
);

DFFPOSX1 _9166_ (
    .CLK(clk_bF$buf66),
    .D(_1761_),
    .Q(\genblk1[2].u_ce.Acalc [3])
);

DFFPOSX1 _9167_ (
    .CLK(clk_bF$buf65),
    .D(_1762_),
    .Q(\genblk1[2].u_ce.Acalc [4])
);

DFFPOSX1 _9168_ (
    .CLK(clk_bF$buf64),
    .D(_1763_),
    .Q(\genblk1[2].u_ce.Acalc [5])
);

DFFPOSX1 _9169_ (
    .CLK(clk_bF$buf63),
    .D(_1764_),
    .Q(\genblk1[2].u_ce.Acalc [6])
);

DFFPOSX1 _9170_ (
    .CLK(clk_bF$buf62),
    .D(_1765_),
    .Q(\genblk1[2].u_ce.Acalc [7])
);

DFFPOSX1 _9171_ (
    .CLK(clk_bF$buf61),
    .D(_1766_),
    .Q(\genblk1[2].u_ce.Acalc [8])
);

DFFPOSX1 _9172_ (
    .CLK(clk_bF$buf60),
    .D(_1767_),
    .Q(\genblk1[2].u_ce.Acalc [9])
);

DFFPOSX1 _9173_ (
    .CLK(clk_bF$buf59),
    .D(_1768_),
    .Q(\genblk1[2].u_ce.Acalc [10])
);

DFFPOSX1 _9174_ (
    .CLK(clk_bF$buf58),
    .D(_1769_),
    .Q(\genblk1[2].u_ce.Acalc [11])
);

DFFPOSX1 _9175_ (
    .CLK(clk_bF$buf57),
    .D(_1770_),
    .Q(\genblk1[2].u_ce.Xin12b [10])
);

DFFPOSX1 _9176_ (
    .CLK(clk_bF$buf56),
    .D(_1771_),
    .Q(\genblk1[2].u_ce.Xin12b [11])
);

DFFPOSX1 _9177_ (
    .CLK(clk_bF$buf55),
    .D(_1772_),
    .Q(\genblk1[2].u_ce.Xin12b [8])
);

DFFPOSX1 _9178_ (
    .CLK(clk_bF$buf54),
    .D(_1773_),
    .Q(\genblk1[2].u_ce.Xin12b [9])
);

DFFPOSX1 _9179_ (
    .CLK(clk_bF$buf53),
    .D(_1774_),
    .Q(\genblk1[2].u_ce.Xin12b [6])
);

DFFPOSX1 _9180_ (
    .CLK(clk_bF$buf52),
    .D(_1775_),
    .Q(\genblk1[2].u_ce.Xin12b [7])
);

DFFPOSX1 _9181_ (
    .CLK(clk_bF$buf51),
    .D(_1776_),
    .Q(\genblk1[2].u_ce.Xin12b [4])
);

DFFPOSX1 _9182_ (
    .CLK(clk_bF$buf50),
    .D(_1777_),
    .Q(\genblk1[2].u_ce.Xin12b [5])
);

DFFPOSX1 _9183_ (
    .CLK(clk_bF$buf49),
    .D(_1778_),
    .Q(\genblk1[2].u_ce.Xin1 [0])
);

DFFPOSX1 _9184_ (
    .CLK(clk_bF$buf48),
    .D(_1779_),
    .Q(\genblk1[2].u_ce.Xin1 [1])
);

DFFPOSX1 _9185_ (
    .CLK(clk_bF$buf47),
    .D(_1780_),
    .Q(\genblk1[2].u_ce.Xin0 [0])
);

DFFPOSX1 _9186_ (
    .CLK(clk_bF$buf46),
    .D(_1781_),
    .Q(\genblk1[2].u_ce.Xin0 [1])
);

DFFPOSX1 _9187_ (
    .CLK(clk_bF$buf45),
    .D(_1782_),
    .Q(\genblk1[2].u_ce.Yin12b [10])
);

DFFPOSX1 _9188_ (
    .CLK(clk_bF$buf44),
    .D(_1783_),
    .Q(\genblk1[2].u_ce.Yin12b [11])
);

DFFPOSX1 _9189_ (
    .CLK(clk_bF$buf43),
    .D(_1784_),
    .Q(\genblk1[2].u_ce.Yin12b [8])
);

DFFPOSX1 _9190_ (
    .CLK(clk_bF$buf42),
    .D(_1785_),
    .Q(\genblk1[2].u_ce.Yin12b [9])
);

DFFPOSX1 _9191_ (
    .CLK(clk_bF$buf41),
    .D(_1786_),
    .Q(\genblk1[2].u_ce.Yin12b [6])
);

DFFPOSX1 _9192_ (
    .CLK(clk_bF$buf40),
    .D(_1787_),
    .Q(\genblk1[2].u_ce.Yin12b [7])
);

DFFPOSX1 _9193_ (
    .CLK(clk_bF$buf39),
    .D(_1788_),
    .Q(\genblk1[2].u_ce.Yin12b [4])
);

DFFPOSX1 _9194_ (
    .CLK(clk_bF$buf38),
    .D(_1789_),
    .Q(\genblk1[2].u_ce.Yin12b [5])
);

DFFPOSX1 _9195_ (
    .CLK(clk_bF$buf37),
    .D(_1790_),
    .Q(\genblk1[2].u_ce.Yin1 [0])
);

DFFPOSX1 _9196_ (
    .CLK(clk_bF$buf36),
    .D(_1791_),
    .Q(\genblk1[2].u_ce.Yin1 [1])
);

DFFPOSX1 _9197_ (
    .CLK(clk_bF$buf35),
    .D(_1792_),
    .Q(\genblk1[2].u_ce.Yin0 [0])
);

DFFPOSX1 _9198_ (
    .CLK(clk_bF$buf34),
    .D(_1793_),
    .Q(\genblk1[2].u_ce.Yin0 [1])
);

DFFPOSX1 _9199_ (
    .CLK(clk_bF$buf33),
    .D(_1794_),
    .Q(\genblk1[2].u_ce.Ain12b [10])
);

DFFPOSX1 _9200_ (
    .CLK(clk_bF$buf32),
    .D(_1795_),
    .Q(\genblk1[2].u_ce.Ain12b [11])
);

DFFPOSX1 _9201_ (
    .CLK(clk_bF$buf31),
    .D(_1796_),
    .Q(\genblk1[2].u_ce.Ain12b [8])
);

DFFPOSX1 _9202_ (
    .CLK(clk_bF$buf30),
    .D(_1797_),
    .Q(\genblk1[2].u_ce.Ain12b [9])
);

DFFPOSX1 _9203_ (
    .CLK(clk_bF$buf29),
    .D(_1798_),
    .Q(\genblk1[2].u_ce.Ain12b [6])
);

DFFPOSX1 _9204_ (
    .CLK(clk_bF$buf28),
    .D(_1799_),
    .Q(\genblk1[2].u_ce.Ain12b [7])
);

DFFPOSX1 _9205_ (
    .CLK(clk_bF$buf27),
    .D(_1800_),
    .Q(\genblk1[2].u_ce.Ain12b [4])
);

DFFPOSX1 _9206_ (
    .CLK(clk_bF$buf26),
    .D(_1801_),
    .Q(\genblk1[2].u_ce.Ain12b [5])
);

DFFPOSX1 _9207_ (
    .CLK(clk_bF$buf25),
    .D(_1802_),
    .Q(\genblk1[2].u_ce.Ain1 [0])
);

DFFPOSX1 _9208_ (
    .CLK(clk_bF$buf24),
    .D(_1803_),
    .Q(\genblk1[2].u_ce.Ain1 [1])
);

DFFPOSX1 _9209_ (
    .CLK(clk_bF$buf23),
    .D(\genblk1[1].u_ce.ISout ),
    .Q(\genblk1[2].u_ce.ISpipe [0])
);

DFFPOSX1 _9210_ (
    .CLK(clk_bF$buf22),
    .D(\genblk1[2].u_ce.ISpipe [0]),
    .Q(\genblk1[2].u_ce.ISpipe [1])
);

DFFPOSX1 _9211_ (
    .CLK(clk_bF$buf21),
    .D(\genblk1[2].u_ce.ISpipe [1]),
    .Q(\genblk1[2].u_ce.ISpipe [2])
);

DFFPOSX1 _9212_ (
    .CLK(clk_bF$buf20),
    .D(\genblk1[2].u_ce.ISpipe [2]),
    .Q(\genblk1[2].u_ce.ISpipe [3])
);

DFFPOSX1 _9213_ (
    .CLK(clk_bF$buf19),
    .D(\genblk1[2].u_ce.ISpipe [3]),
    .Q(\genblk1[2].u_ce.ISpipe [4])
);

DFFPOSX1 _9214_ (
    .CLK(clk_bF$buf18),
    .D(\genblk1[2].u_ce.ISpipe [4]),
    .Q(\genblk1[2].u_ce.ISpipe [5])
);

DFFPOSX1 _9215_ (
    .CLK(clk_bF$buf17),
    .D(\genblk1[2].u_ce.ISpipe [5]),
    .Q(\genblk1[2].u_ce.ISout )
);

DFFPOSX1 _9216_ (
    .CLK(clk_bF$buf16),
    .D(\genblk1[1].u_ce.Vld_bF$buf0 ),
    .Q(\genblk1[2].u_ce.LoadCtl [0])
);

DFFPOSX1 _9217_ (
    .CLK(clk_bF$buf15),
    .D(\genblk1[2].u_ce.LoadCtl_0_bF$buf3 ),
    .Q(\genblk1[2].u_ce.LoadCtl [1])
);

DFFPOSX1 _9218_ (
    .CLK(clk_bF$buf14),
    .D(\genblk1[2].u_ce.LoadCtl [1]),
    .Q(\genblk1[2].u_ce.LoadCtl [2])
);

DFFPOSX1 _9219_ (
    .CLK(clk_bF$buf13),
    .D(\genblk1[2].u_ce.LoadCtl [2]),
    .Q(\genblk1[2].u_ce.LoadCtl [3])
);

DFFPOSX1 _9220_ (
    .CLK(clk_bF$buf12),
    .D(\genblk1[2].u_ce.LoadCtl [3]),
    .Q(\genblk1[2].u_ce.LoadCtl [4])
);

DFFPOSX1 _9221_ (
    .CLK(clk_bF$buf11),
    .D(\genblk1[2].u_ce.LoadCtl [4]),
    .Q(\genblk1[2].u_ce.LoadCtl [5])
);

DFFPOSX1 _9222_ (
    .CLK(clk_bF$buf10),
    .D(\genblk1[2].u_ce.LoadCtl [5]),
    .Q(\genblk1[2].u_ce.Vld )
);

NOR2X1 _9223_ (
    .A(\genblk1[3].u_ce.LoadCtl [3]),
    .B(\genblk1[3].u_ce.LoadCtl [2]),
    .Y(_2690_)
);

INVX1 _9224_ (
    .A(\genblk1[3].u_ce.Acalc [10]),
    .Y(_2691_)
);

NAND2X1 _9225_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(\genblk1[3].u_ce.Acalc [8]),
    .Y(_2692_)
);

OAI21X1 _9226_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(_2691_),
    .C(_2692_),
    .Y(_2693_)
);

INVX2 _9227_ (
    .A(\genblk1[3].u_ce.LoadCtl [2]),
    .Y(_2694_)
);

INVX1 _9228_ (
    .A(\genblk1[3].u_ce.Acalc [4]),
    .Y(_2695_)
);

INVX1 _9229_ (
    .A(\genblk1[3].u_ce.LoadCtl [3]),
    .Y(_2696_)
);

NOR2X1 _9230_ (
    .A(\genblk1[3].u_ce.LoadCtl [2]),
    .B(_2696_),
    .Y(_2697_)
);

NAND2X1 _9231_ (
    .A(\genblk1[3].u_ce.Acalc [6]),
    .B(_2697_),
    .Y(_2698_)
);

OAI21X1 _9232_ (
    .A(_2694_),
    .B(_2695_),
    .C(_2698_),
    .Y(_2699_)
);

AOI21X1 _9233_ (
    .A(_2690_),
    .B(_2693_),
    .C(_2699_),
    .Y(_2700_)
);

NOR2X1 _9234_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[3].u_ce.LoadCtl [1]),
    .Y(_2701_)
);

INVX4 _9235_ (
    .A(_2701_),
    .Y(_2702_)
);

INVX2 _9236_ (
    .A(\genblk1[3].u_ce.LoadCtl [1]),
    .Y(_2703_)
);

NOR2X1 _9237_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_2703_),
    .Y(_2704_)
);

AOI22X1 _9238_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[3].u_ce.Acalc [0]),
    .C(_2704_),
    .D(\genblk1[3].u_ce.Acalc [2]),
    .Y(_2705_)
);

OAI21X1 _9239_ (
    .A(_2702_),
    .B(_2700_),
    .C(_2705_),
    .Y(\a[4] [0])
);

INVX1 _9240_ (
    .A(\genblk1[3].u_ce.Acalc [11]),
    .Y(_2706_)
);

NAND2X1 _9241_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(\genblk1[3].u_ce.Acalc [9]),
    .Y(_2707_)
);

OAI21X1 _9242_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(_2706_),
    .C(_2707_),
    .Y(_2708_)
);

INVX1 _9243_ (
    .A(\genblk1[3].u_ce.Acalc [7]),
    .Y(_2709_)
);

INVX4 _9244_ (
    .A(_2697_),
    .Y(_2710_)
);

NAND2X1 _9245_ (
    .A(\genblk1[3].u_ce.LoadCtl [2]),
    .B(\genblk1[3].u_ce.Acalc [5]),
    .Y(_2711_)
);

OAI21X1 _9246_ (
    .A(_2709_),
    .B(_2710_),
    .C(_2711_),
    .Y(_2712_)
);

AOI21X1 _9247_ (
    .A(_2690_),
    .B(_2708_),
    .C(_2712_),
    .Y(_2713_)
);

AOI22X1 _9248_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\genblk1[3].u_ce.Acalc [1]),
    .C(_2704_),
    .D(\genblk1[3].u_ce.Acalc [3]),
    .Y(_2714_)
);

OAI21X1 _9249_ (
    .A(_2702_),
    .B(_2713_),
    .C(_2714_),
    .Y(\a[4] [1])
);

INVX1 _9250_ (
    .A(\genblk1[3].u_ce.Ycalc [10]),
    .Y(_2715_)
);

NAND2X1 _9251_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(\genblk1[3].u_ce.Ycalc [8]),
    .Y(_2716_)
);

OAI21X1 _9252_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(_2715_),
    .C(_2716_),
    .Y(_2717_)
);

INVX1 _9253_ (
    .A(\genblk1[3].u_ce.Ycalc [6]),
    .Y(_2718_)
);

INVX1 _9254_ (
    .A(\genblk1[3].u_ce.Ycalc [4]),
    .Y(_2719_)
);

OAI22X1 _9255_ (
    .A(_2694_),
    .B(_2719_),
    .C(_2718_),
    .D(_2710_),
    .Y(_2720_)
);

AOI21X1 _9256_ (
    .A(_2690_),
    .B(_2717_),
    .C(_2720_),
    .Y(_2721_)
);

AOI22X1 _9257_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 ),
    .B(\genblk1[3].u_ce.Ycalc [0]),
    .C(_2704_),
    .D(\genblk1[3].u_ce.Ycalc [2]),
    .Y(_2722_)
);

OAI21X1 _9258_ (
    .A(_2702_),
    .B(_2721_),
    .C(_2722_),
    .Y(\genblk1[3].u_ce.Y_ [0])
);

INVX1 _9259_ (
    .A(\genblk1[3].u_ce.Ycalc [11]),
    .Y(_2723_)
);

NAND2X1 _9260_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(\genblk1[3].u_ce.Ycalc [9]),
    .Y(_2724_)
);

OAI21X1 _9261_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(_2723_),
    .C(_2724_),
    .Y(_2725_)
);

INVX1 _9262_ (
    .A(\genblk1[3].u_ce.Ycalc [7]),
    .Y(_2726_)
);

INVX1 _9263_ (
    .A(\genblk1[3].u_ce.Ycalc [5]),
    .Y(_2727_)
);

OAI22X1 _9264_ (
    .A(_2694_),
    .B(_2727_),
    .C(_2726_),
    .D(_2710_),
    .Y(_2728_)
);

AOI21X1 _9265_ (
    .A(_2690_),
    .B(_2725_),
    .C(_2728_),
    .Y(_2729_)
);

AOI22X1 _9266_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\genblk1[3].u_ce.Ycalc [1]),
    .C(_2704_),
    .D(\genblk1[3].u_ce.Ycalc [3]),
    .Y(_2730_)
);

OAI21X1 _9267_ (
    .A(_2702_),
    .B(_2729_),
    .C(_2730_),
    .Y(\genblk1[3].u_ce.Y_ [1])
);

INVX1 _9268_ (
    .A(\genblk1[3].u_ce.Xcalc [2]),
    .Y(_2731_)
);

INVX2 _9269_ (
    .A(_2704_),
    .Y(_2732_)
);

INVX1 _9270_ (
    .A(\genblk1[3].u_ce.Xcalc [4]),
    .Y(_2733_)
);

INVX1 _9271_ (
    .A(\genblk1[3].u_ce.Xcalc [6]),
    .Y(_2734_)
);

NOR2X1 _9272_ (
    .A(_2696_),
    .B(_2734_),
    .Y(_2735_)
);

INVX1 _9273_ (
    .A(\genblk1[3].u_ce.Xcalc [8]),
    .Y(_2736_)
);

NAND2X1 _9274_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(_2736_),
    .Y(_2737_)
);

OAI21X1 _9275_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .B(\genblk1[3].u_ce.Xcalc [10]),
    .C(_2737_),
    .Y(_2738_)
);

NOR2X1 _9276_ (
    .A(\genblk1[3].u_ce.LoadCtl [3]),
    .B(_2738_),
    .Y(_2739_)
);

OAI21X1 _9277_ (
    .A(_2735_),
    .B(_2739_),
    .C(_2694_),
    .Y(_2740_)
);

OAI21X1 _9278_ (
    .A(_2694_),
    .B(_2733_),
    .C(_2740_),
    .Y(_2741_)
);

AOI22X1 _9279_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(\genblk1[3].u_ce.Xcalc [0]),
    .C(_2741_),
    .D(_2701_),
    .Y(_2742_)
);

OAI21X1 _9280_ (
    .A(_2731_),
    .B(_2732_),
    .C(_2742_),
    .Y(\genblk1[3].u_ce.X_ [0])
);

INVX1 _9281_ (
    .A(\genblk1[3].u_ce.LoadCtl [4]),
    .Y(_2743_)
);

INVX1 _9282_ (
    .A(\genblk1[3].u_ce.Xcalc [9]),
    .Y(_2744_)
);

NAND2X1 _9283_ (
    .A(\genblk1[3].u_ce.Xcalc [11]),
    .B(_2743_),
    .Y(_2745_)
);

OAI21X1 _9284_ (
    .A(_2743_),
    .B(_2744_),
    .C(_2745_),
    .Y(_2746_)
);

INVX1 _9285_ (
    .A(\genblk1[3].u_ce.Xcalc [7]),
    .Y(_2747_)
);

INVX1 _9286_ (
    .A(\genblk1[3].u_ce.Xcalc [5]),
    .Y(_2748_)
);

OAI22X1 _9287_ (
    .A(_2694_),
    .B(_2748_),
    .C(_2747_),
    .D(_2710_),
    .Y(_2749_)
);

AOI21X1 _9288_ (
    .A(_2690_),
    .B(_2746_),
    .C(_2749_),
    .Y(_2750_)
);

AOI22X1 _9289_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf2 ),
    .B(\genblk1[3].u_ce.Xcalc [1]),
    .C(_2704_),
    .D(\genblk1[3].u_ce.Xcalc [3]),
    .Y(_2751_)
);

OAI21X1 _9290_ (
    .A(_2702_),
    .B(_2750_),
    .C(_2751_),
    .Y(\genblk1[3].u_ce.X_ [1])
);

INVX1 _9291_ (
    .A(\genblk1[3].u_ce.Ain0 [0]),
    .Y(_2752_)
);

NAND2X1 _9292_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf1 ),
    .B(\a[3] [0]),
    .Y(_2753_)
);

OAI21X1 _9293_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf0 ),
    .B(_2752_),
    .C(_2753_),
    .Y(_2598_)
);

INVX1 _9294_ (
    .A(\genblk1[3].u_ce.Ain0 [1]),
    .Y(_2754_)
);

NAND2X1 _9295_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf4 ),
    .B(\a[3] [1]),
    .Y(_2755_)
);

OAI21X1 _9296_ (
    .A(\genblk1[3].u_ce.LoadCtl_0_bF$buf3 ),
    .B(_2754_),
    .C(_2755_),
    .Y(_2599_)
);

INVX8 _9297_ (
    .A(\genblk1[3].u_ce.Vld_bF$buf0 ),
    .Y(_2756_)
);

NAND2X1 _9298_ (
    .A(\genblk1[3].u_ce.Ycalc [2]),
    .B(_2756__bF$buf2),
    .Y(_2757_)
);

INVX2 _9299_ (
    .A(1'h1),
    .Y(_2758_)
);

NOR2X1 _9300_ (
    .A(1'h0),
    .B(1'h1),
    .Y(_2759_)
);

NAND2X1 _9301_ (
    .A(_2758_),
    .B(_2759_),
    .Y(_2760_)
);

INVX2 _9302_ (
    .A(_2760_),
    .Y(_2761_)
);

INVX8 _9303_ (
    .A(1'h1),
    .Y(_2762_)
);

MUX2X1 _9304_ (
    .A(\genblk1[3].u_ce.Xin12b [4]),
    .B(\genblk1[3].u_ce.Xin1 [1]),
    .S(1'h1),
    .Y(_2763_)
);

MUX2X1 _9305_ (
    .A(\genblk1[3].u_ce.Xin1 [0]),
    .B(\genblk1[3].u_ce.Xin0 [1]),
    .S(1'h1),
    .Y(_2764_)
);

MUX2X1 _9306_ (
    .A(_2764_),
    .B(_2763_),
    .S(_2762__bF$buf4),
    .Y(_2765_)
);

MUX2X1 _9307_ (
    .A(\genblk1[3].u_ce.Xin12b [8]),
    .B(\genblk1[3].u_ce.Xin12b [7]),
    .S(1'h1),
    .Y(_2766_)
);

MUX2X1 _9308_ (
    .A(\genblk1[3].u_ce.Xin12b [6]),
    .B(\genblk1[3].u_ce.Xin12b [5]),
    .S(1'h1),
    .Y(_2767_)
);

MUX2X1 _9309_ (
    .A(_2767_),
    .B(_2766_),
    .S(_2762__bF$buf3),
    .Y(_2768_)
);

MUX2X1 _9310_ (
    .A(_2768_),
    .B(_2765_),
    .S(1'h0),
    .Y(_2769_)
);

INVX1 _9311_ (
    .A(_2769_),
    .Y(_2770_)
);

MUX2X1 _9312_ (
    .A(\genblk1[3].u_ce.Xin1 [1]),
    .B(\genblk1[3].u_ce.Xin1 [0]),
    .S(1'h1),
    .Y(_2771_)
);

MUX2X1 _9313_ (
    .A(\genblk1[3].u_ce.Xin0 [1]),
    .B(\genblk1[3].u_ce.Xin0 [0]),
    .S(1'h1),
    .Y(_2772_)
);

MUX2X1 _9314_ (
    .A(_2772_),
    .B(_2771_),
    .S(_2762__bF$buf2),
    .Y(_2773_)
);

MUX2X1 _9315_ (
    .A(\genblk1[3].u_ce.Xin12b [7]),
    .B(\genblk1[3].u_ce.Xin12b [6]),
    .S(1'h1),
    .Y(_2774_)
);

MUX2X1 _9316_ (
    .A(\genblk1[3].u_ce.Xin12b [5]),
    .B(\genblk1[3].u_ce.Xin12b [4]),
    .S(1'h1),
    .Y(_2775_)
);

MUX2X1 _9317_ (
    .A(_2775_),
    .B(_2774_),
    .S(_2762__bF$buf1),
    .Y(_2776_)
);

MUX2X1 _9318_ (
    .A(_2776_),
    .B(_2773_),
    .S(1'h0),
    .Y(_2777_)
);

OAI21X1 _9319_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2777_),
    .C(_2770_),
    .Y(_2778_)
);

NOR2X1 _9320_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2777_),
    .Y(_2779_)
);

NAND2X1 _9321_ (
    .A(_2769_),
    .B(_2779_),
    .Y(_2780_)
);

NAND3X1 _9322_ (
    .A(\genblk1[3].u_ce.Yin0 [1]),
    .B(_2778_),
    .C(_2780_),
    .Y(_2781_)
);

NOR2X1 _9323_ (
    .A(\genblk1[3].u_ce.Yin0 [0]),
    .B(_2777_),
    .Y(_2782_)
);

AOI21X1 _9324_ (
    .A(_2780_),
    .B(_2778_),
    .C(\genblk1[3].u_ce.Yin0 [1]),
    .Y(_2783_)
);

OAI21X1 _9325_ (
    .A(_2782_),
    .B(_2783_),
    .C(_2781_),
    .Y(_2784_)
);

INVX1 _9326_ (
    .A(\genblk1[3].u_ce.Yin1 [0]),
    .Y(_2785_)
);

MUX2X1 _9327_ (
    .A(\genblk1[3].u_ce.Xin12b [9]),
    .B(\genblk1[3].u_ce.Xin12b [8]),
    .S(1'h1),
    .Y(_2786_)
);

MUX2X1 _9328_ (
    .A(_2786_),
    .B(_2774_),
    .S(1'h1),
    .Y(_2787_)
);

AND2X2 _9329_ (
    .A(_2787_),
    .B(1'h0),
    .Y(_2788_)
);

INVX4 _9330_ (
    .A(1'h0),
    .Y(_2789_)
);

NAND2X1 _9331_ (
    .A(_2789__bF$buf3),
    .B(_2762__bF$buf0),
    .Y(_2790_)
);

NAND2X1 _9332_ (
    .A(1'h1),
    .B(_2789__bF$buf2),
    .Y(_2791_)
);

OAI22X1 _9333_ (
    .A(_2790_),
    .B(_2771_),
    .C(_2775_),
    .D(_2791_),
    .Y(_2792_)
);

INVX1 _9334_ (
    .A(\genblk1[3].u_ce.Xin1 [1]),
    .Y(_2793_)
);

NAND2X1 _9335_ (
    .A(_2758_),
    .B(_2793_),
    .Y(_2794_)
);

INVX1 _9336_ (
    .A(\genblk1[3].u_ce.Xin12b [4]),
    .Y(_2795_)
);

NAND2X1 _9337_ (
    .A(1'h1),
    .B(_2795_),
    .Y(_2796_)
);

NAND3X1 _9338_ (
    .A(1'h1),
    .B(_2796_),
    .C(_2794_),
    .Y(_2797_)
);

INVX1 _9339_ (
    .A(\genblk1[3].u_ce.Xin0 [1]),
    .Y(_2798_)
);

NAND2X1 _9340_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Xin1 [0]),
    .Y(_2799_)
);

OAI21X1 _9341_ (
    .A(1'h1),
    .B(_2798_),
    .C(_2799_),
    .Y(_2800_)
);

NAND2X1 _9342_ (
    .A(_2762__bF$buf4),
    .B(_2800_),
    .Y(_2801_)
);

NAND3X1 _9343_ (
    .A(_2789__bF$buf1),
    .B(_2797_),
    .C(_2801_),
    .Y(_2802_)
);

INVX1 _9344_ (
    .A(\genblk1[3].u_ce.Xin12b [5]),
    .Y(_2803_)
);

NAND2X1 _9345_ (
    .A(_2758_),
    .B(_2803_),
    .Y(_2804_)
);

INVX1 _9346_ (
    .A(\genblk1[3].u_ce.Xin12b [6]),
    .Y(_2805_)
);

NAND2X1 _9347_ (
    .A(1'h1),
    .B(_2805_),
    .Y(_2806_)
);

NAND3X1 _9348_ (
    .A(_2762__bF$buf3),
    .B(_2806_),
    .C(_2804_),
    .Y(_2807_)
);

INVX1 _9349_ (
    .A(\genblk1[3].u_ce.Xin12b [7]),
    .Y(_2808_)
);

NAND2X1 _9350_ (
    .A(_2758_),
    .B(_2808_),
    .Y(_2809_)
);

INVX1 _9351_ (
    .A(\genblk1[3].u_ce.Xin12b [8]),
    .Y(_2810_)
);

NAND2X1 _9352_ (
    .A(1'h1),
    .B(_2810_),
    .Y(_2811_)
);

NAND3X1 _9353_ (
    .A(1'h1),
    .B(_2811_),
    .C(_2809_),
    .Y(_2812_)
);

NAND3X1 _9354_ (
    .A(1'h0),
    .B(_2807_),
    .C(_2812_),
    .Y(_2813_)
);

INVX1 _9355_ (
    .A(\genblk1[3].u_ce.Xin1 [0]),
    .Y(_2814_)
);

NAND2X1 _9356_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Xin1 [1]),
    .Y(_2815_)
);

OAI21X1 _9357_ (
    .A(1'h1),
    .B(_2814_),
    .C(_2815_),
    .Y(_2816_)
);

NAND2X1 _9358_ (
    .A(1'h1),
    .B(_2816_),
    .Y(_2817_)
);

INVX1 _9359_ (
    .A(\genblk1[3].u_ce.Xin0 [0]),
    .Y(_2818_)
);

NAND2X1 _9360_ (
    .A(\genblk1[3].u_ce.Xin0 [1]),
    .B(1'h1),
    .Y(_2819_)
);

OAI21X1 _9361_ (
    .A(1'h1),
    .B(_2818_),
    .C(_2819_),
    .Y(_2820_)
);

NAND2X1 _9362_ (
    .A(_2762__bF$buf2),
    .B(_2820_),
    .Y(_2821_)
);

NAND3X1 _9363_ (
    .A(_2789__bF$buf0),
    .B(_2817_),
    .C(_2821_),
    .Y(_2822_)
);

NAND2X1 _9364_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Xin12b [5]),
    .Y(_2823_)
);

OAI21X1 _9365_ (
    .A(1'h1),
    .B(_2795_),
    .C(_2823_),
    .Y(_2824_)
);

NAND2X1 _9366_ (
    .A(_2762__bF$buf1),
    .B(_2824_),
    .Y(_2825_)
);

NAND2X1 _9367_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Xin12b [7]),
    .Y(_2826_)
);

OAI21X1 _9368_ (
    .A(1'h1),
    .B(_2805_),
    .C(_2826_),
    .Y(_2827_)
);

NAND2X1 _9369_ (
    .A(1'h1),
    .B(_2827_),
    .Y(_2828_)
);

NAND3X1 _9370_ (
    .A(1'h0),
    .B(_2825_),
    .C(_2828_),
    .Y(_2829_)
);

AOI22X1 _9371_ (
    .A(_2802_),
    .B(_2813_),
    .C(_2822_),
    .D(_2829_),
    .Y(_2830_)
);

NOR2X1 _9372_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .B(_2830_),
    .Y(_2831_)
);

OAI21X1 _9373_ (
    .A(_2788_),
    .B(_2792_),
    .C(_2831_),
    .Y(_2832_)
);

AOI21X1 _9374_ (
    .A(1'h0),
    .B(_2787_),
    .C(_2792_),
    .Y(_2833_)
);

OAI21X1 _9375_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2830_),
    .C(_2833_),
    .Y(_2834_)
);

NAND3X1 _9376_ (
    .A(_2785_),
    .B(_2834_),
    .C(_2832_),
    .Y(_2835_)
);

NAND2X1 _9377_ (
    .A(_2833_),
    .B(_2831_),
    .Y(_2836_)
);

OAI22X1 _9378_ (
    .A(_2788_),
    .B(_2792_),
    .C(\genblk1[3].u_ce.Ain12b_11_bF$buf4 ),
    .D(_2830_),
    .Y(_2837_)
);

NAND3X1 _9379_ (
    .A(\genblk1[3].u_ce.Yin1 [0]),
    .B(_2837_),
    .C(_2836_),
    .Y(_2838_)
);

NAND3X1 _9380_ (
    .A(_2835_),
    .B(_2838_),
    .C(_2784_),
    .Y(_2839_)
);

INVX1 _9381_ (
    .A(\genblk1[3].u_ce.Yin0 [1]),
    .Y(_2840_)
);

NAND2X1 _9382_ (
    .A(_2770_),
    .B(_2779_),
    .Y(_2841_)
);

OAI21X1 _9383_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2777_),
    .C(_2769_),
    .Y(_2842_)
);

AOI21X1 _9384_ (
    .A(_2841_),
    .B(_2842_),
    .C(_2840_),
    .Y(_2843_)
);

INVX1 _9385_ (
    .A(_2782_),
    .Y(_2844_)
);

NAND3X1 _9386_ (
    .A(_2840_),
    .B(_2842_),
    .C(_2841_),
    .Y(_2845_)
);

AOI21X1 _9387_ (
    .A(_2844_),
    .B(_2845_),
    .C(_2843_),
    .Y(_2846_)
);

AOI21X1 _9388_ (
    .A(_2836_),
    .B(_2837_),
    .C(\genblk1[3].u_ce.Yin1 [0]),
    .Y(_2847_)
);

AOI21X1 _9389_ (
    .A(_2832_),
    .B(_2834_),
    .C(_2785_),
    .Y(_2848_)
);

OAI21X1 _9390_ (
    .A(_2847_),
    .B(_2848_),
    .C(_2846_),
    .Y(_2849_)
);

AOI21X1 _9391_ (
    .A(_2839_),
    .B(_2849_),
    .C(_2761_),
    .Y(_2850_)
);

INVX8 _9392_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .Y(_2851_)
);

NAND3X1 _9393_ (
    .A(_2789__bF$buf3),
    .B(_2758_),
    .C(_2851__bF$buf3),
    .Y(_2852_)
);

OAI21X1 _9394_ (
    .A(1'h1),
    .B(_2852_),
    .C(\genblk1[3].u_ce.Vld_bF$buf4 ),
    .Y(_2853_)
);

OAI21X1 _9395_ (
    .A(_2853_),
    .B(_2850_),
    .C(_2757_),
    .Y(_2600_)
);

INVX1 _9396_ (
    .A(\genblk1[3].u_ce.Ycalc [3]),
    .Y(_2854_)
);

INVX1 _9397_ (
    .A(\genblk1[3].u_ce.Xin12b [9]),
    .Y(_2855_)
);

NAND2X1 _9398_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Xin12b [10]),
    .Y(_2856_)
);

OAI21X1 _9399_ (
    .A(1'h1),
    .B(_2855_),
    .C(_2856_),
    .Y(_2857_)
);

NAND2X1 _9400_ (
    .A(1'h1),
    .B(_2857_),
    .Y(_2858_)
);

OAI21X1 _9401_ (
    .A(1'h1),
    .B(_2766_),
    .C(_2858_),
    .Y(_2859_)
);

OAI22X1 _9402_ (
    .A(_2790_),
    .B(_2763_),
    .C(_2767_),
    .D(_2791_),
    .Y(_2860_)
);

AOI21X1 _9403_ (
    .A(_2859_),
    .B(1'h0),
    .C(_2860_),
    .Y(_2861_)
);

NAND3X1 _9404_ (
    .A(_2833_),
    .B(_2769_),
    .C(_2777_),
    .Y(_2862_)
);

INVX1 _9405_ (
    .A(_2862_),
    .Y(_2863_)
);

NOR2X1 _9406_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .B(_2863_),
    .Y(_2864_)
);

NAND2X1 _9407_ (
    .A(_2861_),
    .B(_2864_),
    .Y(_2865_)
);

INVX1 _9408_ (
    .A(_2861_),
    .Y(_2866_)
);

OAI21X1 _9409_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2863_),
    .C(_2866_),
    .Y(_2867_)
);

AOI21X1 _9410_ (
    .A(_2865_),
    .B(_2867_),
    .C(\genblk1[3].u_ce.Yin1 [1]),
    .Y(_2868_)
);

AOI21X1 _9411_ (
    .A(_2784_),
    .B(_2835_),
    .C(_2848_),
    .Y(_2869_)
);

NAND3X1 _9412_ (
    .A(\genblk1[3].u_ce.Yin1 [1]),
    .B(_2867_),
    .C(_2865_),
    .Y(_2870_)
);

NAND2X1 _9413_ (
    .A(_2870_),
    .B(_2869_),
    .Y(_2871_)
);

OAI21X1 _9414_ (
    .A(_2847_),
    .B(_2846_),
    .C(_2838_),
    .Y(_2872_)
);

INVX1 _9415_ (
    .A(\genblk1[3].u_ce.Yin1 [1]),
    .Y(_2873_)
);

NAND2X1 _9416_ (
    .A(_2866_),
    .B(_2864_),
    .Y(_2874_)
);

OAI21X1 _9417_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf4 ),
    .B(_2863_),
    .C(_2861_),
    .Y(_2875_)
);

AOI21X1 _9418_ (
    .A(_2874_),
    .B(_2875_),
    .C(_2873_),
    .Y(_2876_)
);

OAI21X1 _9419_ (
    .A(_2868_),
    .B(_2876_),
    .C(_2872_),
    .Y(_2877_)
);

OAI21X1 _9420_ (
    .A(_2868_),
    .B(_2871_),
    .C(_2877_),
    .Y(_2878_)
);

OAI21X1 _9421_ (
    .A(_2851__bF$buf2),
    .B(_2760_),
    .C(\genblk1[3].u_ce.Vld_bF$buf3 ),
    .Y(_2879_)
);

INVX1 _9422_ (
    .A(_2879_),
    .Y(_2880_)
);

OAI21X1 _9423_ (
    .A(_2761_),
    .B(_2878_),
    .C(_2880_),
    .Y(_2881_)
);

OAI21X1 _9424_ (
    .A(_2854_),
    .B(\genblk1[3].u_ce.Vld_bF$buf2 ),
    .C(_2881_),
    .Y(_2601_)
);

INVX1 _9425_ (
    .A(_2853_),
    .Y(_2882_)
);

INVX1 _9426_ (
    .A(\genblk1[3].u_ce.Yin12b [4]),
    .Y(_2883_)
);

NAND3X1 _9427_ (
    .A(_2833_),
    .B(_2861_),
    .C(_2830_),
    .Y(_2884_)
);

INVX1 _9428_ (
    .A(\genblk1[3].u_ce.Xin12b [10]),
    .Y(_2885_)
);

NAND2X1 _9429_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Xin12b [11]),
    .Y(_2886_)
);

OAI21X1 _9430_ (
    .A(1'h1),
    .B(_2885_),
    .C(_2886_),
    .Y(_2887_)
);

NAND2X1 _9431_ (
    .A(_2762__bF$buf0),
    .B(_2786_),
    .Y(_2888_)
);

OAI21X1 _9432_ (
    .A(_2762__bF$buf4),
    .B(_2887_),
    .C(_2888_),
    .Y(_2889_)
);

NAND2X1 _9433_ (
    .A(_2789__bF$buf2),
    .B(_2776_),
    .Y(_2890_)
);

OAI21X1 _9434_ (
    .A(_2789__bF$buf1),
    .B(_2889_),
    .C(_2890_),
    .Y(_2891_)
);

INVX1 _9435_ (
    .A(_2891_),
    .Y(_2892_)
);

NAND3X1 _9436_ (
    .A(_2851__bF$buf1),
    .B(_2892_),
    .C(_2884_),
    .Y(_2893_)
);

INVX1 _9437_ (
    .A(_2893_),
    .Y(_2894_)
);

AOI21X1 _9438_ (
    .A(_2884_),
    .B(_2851__bF$buf0),
    .C(_2892_),
    .Y(_2895_)
);

OAI21X1 _9439_ (
    .A(_2895_),
    .B(_2894_),
    .C(_2883_),
    .Y(_2896_)
);

OAI21X1 _9440_ (
    .A(_2862_),
    .B(_2866_),
    .C(_2851__bF$buf5),
    .Y(_2897_)
);

NAND2X1 _9441_ (
    .A(_2891_),
    .B(_2897_),
    .Y(_2898_)
);

NAND3X1 _9442_ (
    .A(\genblk1[3].u_ce.Yin12b [4]),
    .B(_2893_),
    .C(_2898_),
    .Y(_2899_)
);

NAND2X1 _9443_ (
    .A(_2899_),
    .B(_2896_),
    .Y(_2900_)
);

INVX1 _9444_ (
    .A(_2868_),
    .Y(_2901_)
);

OAI21X1 _9445_ (
    .A(_2876_),
    .B(_2872_),
    .C(_2901_),
    .Y(_2902_)
);

AOI21X1 _9446_ (
    .A(_2902_),
    .B(_2900_),
    .C(_2761_),
    .Y(_2903_)
);

OAI21X1 _9447_ (
    .A(_2900_),
    .B(_2902_),
    .C(_2903_),
    .Y(_2904_)
);

AOI22X1 _9448_ (
    .A(_2719_),
    .B(_2756__bF$buf1),
    .C(_2904_),
    .D(_2882_),
    .Y(_2602_)
);

INVX1 _9449_ (
    .A(_2899_),
    .Y(_2905_)
);

AOI21X1 _9450_ (
    .A(_2869_),
    .B(_2870_),
    .C(_2868_),
    .Y(_2906_)
);

AOI21X1 _9451_ (
    .A(_2906_),
    .B(_2896_),
    .C(_2905_),
    .Y(_2907_)
);

INVX1 _9452_ (
    .A(\genblk1[3].u_ce.Yin12b [5]),
    .Y(_2908_)
);

NAND3X1 _9453_ (
    .A(_2861_),
    .B(_2892_),
    .C(_2863_),
    .Y(_2909_)
);

INVX1 _9454_ (
    .A(\genblk1[3].u_ce.Xin12b [11]),
    .Y(_2910_)
);

NOR2X1 _9455_ (
    .A(_2762__bF$buf3),
    .B(_2910_),
    .Y(_2911_)
);

AOI21X1 _9456_ (
    .A(_2762__bF$buf2),
    .B(_2857_),
    .C(_2911_),
    .Y(_2912_)
);

NAND2X1 _9457_ (
    .A(_2789__bF$buf0),
    .B(_2768_),
    .Y(_2913_)
);

OAI21X1 _9458_ (
    .A(_2789__bF$buf3),
    .B(_2912_),
    .C(_2913_),
    .Y(_2914_)
);

NAND3X1 _9459_ (
    .A(_2851__bF$buf4),
    .B(_2914_),
    .C(_2909_),
    .Y(_2915_)
);

INVX1 _9460_ (
    .A(_2914_),
    .Y(_2916_)
);

OAI21X1 _9461_ (
    .A(_2891_),
    .B(_2884_),
    .C(_2851__bF$buf3),
    .Y(_2917_)
);

NAND2X1 _9462_ (
    .A(_2916_),
    .B(_2917_),
    .Y(_2918_)
);

NAND3X1 _9463_ (
    .A(_2908_),
    .B(_2918_),
    .C(_2915_),
    .Y(_2919_)
);

NAND3X1 _9464_ (
    .A(_2851__bF$buf2),
    .B(_2916_),
    .C(_2909_),
    .Y(_2920_)
);

NAND2X1 _9465_ (
    .A(_2914_),
    .B(_2917_),
    .Y(_2921_)
);

NAND3X1 _9466_ (
    .A(\genblk1[3].u_ce.Yin12b [5]),
    .B(_2921_),
    .C(_2920_),
    .Y(_2922_)
);

NAND2X1 _9467_ (
    .A(_2919_),
    .B(_2922_),
    .Y(_2923_)
);

INVX1 _9468_ (
    .A(_2923_),
    .Y(_2924_)
);

NOR2X1 _9469_ (
    .A(_2924_),
    .B(_2907_),
    .Y(_2925_)
);

OAI21X1 _9470_ (
    .A(_2900_),
    .B(_2902_),
    .C(_2899_),
    .Y(_2926_)
);

OAI21X1 _9471_ (
    .A(_2923_),
    .B(_2926_),
    .C(_2760_),
    .Y(_2927_)
);

OAI21X1 _9472_ (
    .A(_2927_),
    .B(_2925_),
    .C(_2882_),
    .Y(_2928_)
);

OAI21X1 _9473_ (
    .A(_2727_),
    .B(\genblk1[3].u_ce.Vld_bF$buf1 ),
    .C(_2928_),
    .Y(_2603_)
);

NOR2X1 _9474_ (
    .A(_2900_),
    .B(_2923_),
    .Y(_2929_)
);

OAI21X1 _9475_ (
    .A(_2899_),
    .B(_2923_),
    .C(_2922_),
    .Y(_2930_)
);

AOI21X1 _9476_ (
    .A(_2929_),
    .B(_2906_),
    .C(_2930_),
    .Y(_2931_)
);

INVX1 _9477_ (
    .A(\genblk1[3].u_ce.Yin12b [6]),
    .Y(_2932_)
);

NOR2X1 _9478_ (
    .A(_2891_),
    .B(_2884_),
    .Y(_2933_)
);

NAND2X1 _9479_ (
    .A(_2916_),
    .B(_2933_),
    .Y(_2934_)
);

AOI21X1 _9480_ (
    .A(_2762__bF$buf1),
    .B(_2887_),
    .C(_2911_),
    .Y(_2935_)
);

NAND2X1 _9481_ (
    .A(_2789__bF$buf2),
    .B(_2787_),
    .Y(_2936_)
);

OAI21X1 _9482_ (
    .A(_2789__bF$buf1),
    .B(_2935_),
    .C(_2936_),
    .Y(_2937_)
);

NAND3X1 _9483_ (
    .A(_2851__bF$buf1),
    .B(_2937_),
    .C(_2934_),
    .Y(_2938_)
);

NOR3X1 _9484_ (
    .A(_2891_),
    .B(_2914_),
    .C(_2884_),
    .Y(_2939_)
);

INVX1 _9485_ (
    .A(_2937_),
    .Y(_2940_)
);

OAI21X1 _9486_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .B(_2939_),
    .C(_2940_),
    .Y(_2941_)
);

NAND3X1 _9487_ (
    .A(_2932_),
    .B(_2941_),
    .C(_2938_),
    .Y(_2942_)
);

NAND3X1 _9488_ (
    .A(_2851__bF$buf0),
    .B(_2940_),
    .C(_2934_),
    .Y(_2943_)
);

OAI21X1 _9489_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .B(_2939_),
    .C(_2937_),
    .Y(_2944_)
);

NAND3X1 _9490_ (
    .A(\genblk1[3].u_ce.Yin12b [6]),
    .B(_2944_),
    .C(_2943_),
    .Y(_2945_)
);

AND2X2 _9491_ (
    .A(_2942_),
    .B(_2945_),
    .Y(_2946_)
);

INVX1 _9492_ (
    .A(_2946_),
    .Y(_2947_)
);

AOI21X1 _9493_ (
    .A(_2931_),
    .B(_2947_),
    .C(_2761_),
    .Y(_2948_)
);

OAI21X1 _9494_ (
    .A(_2931_),
    .B(_2947_),
    .C(_2948_),
    .Y(_2949_)
);

AOI22X1 _9495_ (
    .A(_2718_),
    .B(_2756__bF$buf0),
    .C(_2949_),
    .D(_2882_),
    .Y(_2604_)
);

AND2X2 _9496_ (
    .A(_2896_),
    .B(_2899_),
    .Y(_2950_)
);

NAND3X1 _9497_ (
    .A(_2919_),
    .B(_2922_),
    .C(_2950_),
    .Y(_2951_)
);

INVX1 _9498_ (
    .A(_2922_),
    .Y(_2952_)
);

AOI21X1 _9499_ (
    .A(_2905_),
    .B(_2919_),
    .C(_2952_),
    .Y(_2953_)
);

OAI21X1 _9500_ (
    .A(_2902_),
    .B(_2951_),
    .C(_2953_),
    .Y(_2954_)
);

INVX1 _9501_ (
    .A(_2945_),
    .Y(_2955_)
);

AOI21X1 _9502_ (
    .A(_2954_),
    .B(_2942_),
    .C(_2955_),
    .Y(_2956_)
);

INVX1 _9503_ (
    .A(\genblk1[3].u_ce.Yin12b [7]),
    .Y(_2957_)
);

NAND2X1 _9504_ (
    .A(_2940_),
    .B(_2939_),
    .Y(_2958_)
);

NOR2X1 _9505_ (
    .A(_2789__bF$buf0),
    .B(_2910_),
    .Y(_2959_)
);

AOI21X1 _9506_ (
    .A(_2859_),
    .B(_2789__bF$buf3),
    .C(_2959_),
    .Y(_2960_)
);

INVX1 _9507_ (
    .A(_2960_),
    .Y(_2961_)
);

NAND3X1 _9508_ (
    .A(_2851__bF$buf5),
    .B(_2961_),
    .C(_2958_),
    .Y(_2962_)
);

AND2X2 _9509_ (
    .A(_2939_),
    .B(_2940_),
    .Y(_2963_)
);

OAI21X1 _9510_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .B(_2963_),
    .C(_2960_),
    .Y(_2964_)
);

NAND3X1 _9511_ (
    .A(_2957_),
    .B(_2962_),
    .C(_2964_),
    .Y(_2965_)
);

NAND3X1 _9512_ (
    .A(_2851__bF$buf4),
    .B(_2960_),
    .C(_2958_),
    .Y(_2966_)
);

OAI21X1 _9513_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .B(_2963_),
    .C(_2961_),
    .Y(_2967_)
);

NAND3X1 _9514_ (
    .A(\genblk1[3].u_ce.Yin12b [7]),
    .B(_2966_),
    .C(_2967_),
    .Y(_2968_)
);

AND2X2 _9515_ (
    .A(_2965_),
    .B(_2968_),
    .Y(_2969_)
);

NOR2X1 _9516_ (
    .A(_2969_),
    .B(_2956_),
    .Y(_2970_)
);

NAND2X1 _9517_ (
    .A(_2758_),
    .B(_2762__bF$buf0),
    .Y(_2971_)
);

NAND2X1 _9518_ (
    .A(_2969_),
    .B(_2956_),
    .Y(_2972_)
);

OAI21X1 _9519_ (
    .A(1'h0),
    .B(_2971_),
    .C(_2972_),
    .Y(_2973_)
);

OAI21X1 _9520_ (
    .A(_2970_),
    .B(_2973_),
    .C(_2880_),
    .Y(_2974_)
);

OAI21X1 _9521_ (
    .A(_2726_),
    .B(\genblk1[3].u_ce.Vld_bF$buf0 ),
    .C(_2974_),
    .Y(_2605_)
);

INVX1 _9522_ (
    .A(\genblk1[3].u_ce.Ycalc [8]),
    .Y(_2975_)
);

AOI21X1 _9523_ (
    .A(_2964_),
    .B(_2962_),
    .C(_2957_),
    .Y(_2976_)
);

OAI21X1 _9524_ (
    .A(_2955_),
    .B(_2976_),
    .C(_2965_),
    .Y(_2977_)
);

NAND3X1 _9525_ (
    .A(_2946_),
    .B(_2969_),
    .C(_2954_),
    .Y(_2978_)
);

INVX1 _9526_ (
    .A(\genblk1[3].u_ce.Yin12b [8]),
    .Y(_2979_)
);

NAND3X1 _9527_ (
    .A(_2940_),
    .B(_2960_),
    .C(_2939_),
    .Y(_2980_)
);

INVX1 _9528_ (
    .A(_2959_),
    .Y(_2981_)
);

OAI21X1 _9529_ (
    .A(1'h0),
    .B(_2889_),
    .C(_2981_),
    .Y(_2982_)
);

NAND3X1 _9530_ (
    .A(_2851__bF$buf3),
    .B(_2982_),
    .C(_2980_),
    .Y(_2983_)
);

INVX1 _9531_ (
    .A(_2982_),
    .Y(_2984_)
);

NAND2X1 _9532_ (
    .A(_2851__bF$buf2),
    .B(_2980_),
    .Y(_2985_)
);

NAND2X1 _9533_ (
    .A(_2984_),
    .B(_2985_),
    .Y(_2986_)
);

NAND3X1 _9534_ (
    .A(_2979_),
    .B(_2983_),
    .C(_2986_),
    .Y(_2987_)
);

NAND3X1 _9535_ (
    .A(_2851__bF$buf1),
    .B(_2984_),
    .C(_2980_),
    .Y(_2988_)
);

NAND2X1 _9536_ (
    .A(_2982_),
    .B(_2985_),
    .Y(_2989_)
);

NAND3X1 _9537_ (
    .A(\genblk1[3].u_ce.Yin12b [8]),
    .B(_2988_),
    .C(_2989_),
    .Y(_2990_)
);

AND2X2 _9538_ (
    .A(_2987_),
    .B(_2990_),
    .Y(_2991_)
);

INVX1 _9539_ (
    .A(_2991_),
    .Y(_2992_)
);

AOI21X1 _9540_ (
    .A(_2978_),
    .B(_2977_),
    .C(_2992_),
    .Y(_2993_)
);

NAND3X1 _9541_ (
    .A(_2965_),
    .B(_2968_),
    .C(_2946_),
    .Y(_2994_)
);

OAI21X1 _9542_ (
    .A(_2994_),
    .B(_2931_),
    .C(_2977_),
    .Y(_2995_)
);

OAI21X1 _9543_ (
    .A(_2991_),
    .B(_2995_),
    .C(_2760_),
    .Y(_2996_)
);

OR2X2 _9544_ (
    .A(_2996_),
    .B(_2993_),
    .Y(_2997_)
);

AOI22X1 _9545_ (
    .A(_2975_),
    .B(_2756__bF$buf4),
    .C(_2997_),
    .D(_2880_),
    .Y(_2606_)
);

INVX1 _9546_ (
    .A(\genblk1[3].u_ce.Ycalc [9]),
    .Y(_2998_)
);

INVX1 _9547_ (
    .A(_2990_),
    .Y(_2999_)
);

NOR2X1 _9548_ (
    .A(_2999_),
    .B(_2993_),
    .Y(_3000_)
);

INVX1 _9549_ (
    .A(\genblk1[3].u_ce.Yin12b [9]),
    .Y(_3001_)
);

OAI21X1 _9550_ (
    .A(1'h0),
    .B(_2912_),
    .C(_2981_),
    .Y(_3002_)
);

INVX1 _9551_ (
    .A(_3002_),
    .Y(_3003_)
);

OAI21X1 _9552_ (
    .A(_2982_),
    .B(_2980_),
    .C(_2851__bF$buf0),
    .Y(_3004_)
);

NAND2X1 _9553_ (
    .A(_3003_),
    .B(_3004_),
    .Y(_3005_)
);

NAND3X1 _9554_ (
    .A(_2960_),
    .B(_2984_),
    .C(_2963_),
    .Y(_3006_)
);

NAND3X1 _9555_ (
    .A(_2851__bF$buf5),
    .B(_3002_),
    .C(_3006_),
    .Y(_3007_)
);

NAND3X1 _9556_ (
    .A(_3001_),
    .B(_3005_),
    .C(_3007_),
    .Y(_3008_)
);

AND2X2 _9557_ (
    .A(_3004_),
    .B(_3003_),
    .Y(_3009_)
);

NOR2X1 _9558_ (
    .A(_3003_),
    .B(_3004_),
    .Y(_3010_)
);

OAI21X1 _9559_ (
    .A(_3010_),
    .B(_3009_),
    .C(\genblk1[3].u_ce.Yin12b [9]),
    .Y(_3011_)
);

NAND2X1 _9560_ (
    .A(_3008_),
    .B(_3011_),
    .Y(_3012_)
);

AOI21X1 _9561_ (
    .A(_3000_),
    .B(_3012_),
    .C(_2761_),
    .Y(_3013_)
);

OAI21X1 _9562_ (
    .A(_3000_),
    .B(_3012_),
    .C(_3013_),
    .Y(_3014_)
);

AOI22X1 _9563_ (
    .A(_2998_),
    .B(_2756__bF$buf3),
    .C(_3014_),
    .D(_2880_),
    .Y(_2607_)
);

OAI21X1 _9564_ (
    .A(_2990_),
    .B(_3012_),
    .C(_3011_),
    .Y(_3015_)
);

NAND3X1 _9565_ (
    .A(_3008_),
    .B(_3011_),
    .C(_2991_),
    .Y(_3016_)
);

AOI21X1 _9566_ (
    .A(_2977_),
    .B(_2978_),
    .C(_3016_),
    .Y(_3017_)
);

INVX1 _9567_ (
    .A(\genblk1[3].u_ce.Yin12b [10]),
    .Y(_3018_)
);

OAI21X1 _9568_ (
    .A(1'h0),
    .B(_2935_),
    .C(_2981_),
    .Y(_3019_)
);

INVX1 _9569_ (
    .A(_3019_),
    .Y(_3020_)
);

OAI21X1 _9570_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf4 ),
    .B(_3003_),
    .C(_3004_),
    .Y(_3021_)
);

NAND2X1 _9571_ (
    .A(_3020_),
    .B(_3021_),
    .Y(_3022_)
);

OAI21X1 _9572_ (
    .A(_3002_),
    .B(_3006_),
    .C(_2851__bF$buf4),
    .Y(_3023_)
);

NAND2X1 _9573_ (
    .A(_3019_),
    .B(_3023_),
    .Y(_3024_)
);

NAND2X1 _9574_ (
    .A(_3022_),
    .B(_3024_),
    .Y(_3025_)
);

NAND2X1 _9575_ (
    .A(_3018_),
    .B(_3025_),
    .Y(_3026_)
);

NAND3X1 _9576_ (
    .A(\genblk1[3].u_ce.Yin12b [10]),
    .B(_3022_),
    .C(_3024_),
    .Y(_3027_)
);

AND2X2 _9577_ (
    .A(_3026_),
    .B(_3027_),
    .Y(_3028_)
);

OAI21X1 _9578_ (
    .A(_3015_),
    .B(_3017_),
    .C(_3028_),
    .Y(_3029_)
);

INVX1 _9579_ (
    .A(_3011_),
    .Y(_3030_)
);

AOI21X1 _9580_ (
    .A(_2999_),
    .B(_3008_),
    .C(_3030_),
    .Y(_3031_)
);

AND2X2 _9581_ (
    .A(_3011_),
    .B(_3008_),
    .Y(_3032_)
);

NAND3X1 _9582_ (
    .A(_2991_),
    .B(_3032_),
    .C(_2995_),
    .Y(_3033_)
);

NAND2X1 _9583_ (
    .A(_3027_),
    .B(_3026_),
    .Y(_3034_)
);

NAND3X1 _9584_ (
    .A(_3031_),
    .B(_3034_),
    .C(_3033_),
    .Y(_3035_)
);

NAND3X1 _9585_ (
    .A(_2760_),
    .B(_3035_),
    .C(_3029_),
    .Y(_3036_)
);

AOI22X1 _9586_ (
    .A(_2715_),
    .B(_2756__bF$buf2),
    .C(_3036_),
    .D(_2882_),
    .Y(_2608_)
);

INVX1 _9587_ (
    .A(_3027_),
    .Y(_3037_)
);

AOI21X1 _9588_ (
    .A(_3033_),
    .B(_3031_),
    .C(_3034_),
    .Y(_3038_)
);

OAI21X1 _9589_ (
    .A(_3019_),
    .B(_3021_),
    .C(_2851__bF$buf3),
    .Y(_3039_)
);

INVX1 _9590_ (
    .A(_3039_),
    .Y(_3040_)
);

NAND2X1 _9591_ (
    .A(\genblk1[3].u_ce.Yin12b [11]),
    .B(_2910_),
    .Y(_3041_)
);

INVX1 _9592_ (
    .A(\genblk1[3].u_ce.Yin12b [11]),
    .Y(_3042_)
);

NAND2X1 _9593_ (
    .A(\genblk1[3].u_ce.Xin12b [11]),
    .B(_3042_),
    .Y(_3043_)
);

NAND2X1 _9594_ (
    .A(_3041_),
    .B(_3043_),
    .Y(_3044_)
);

OR2X2 _9595_ (
    .A(_3040_),
    .B(_3044_),
    .Y(_3045_)
);

NAND2X1 _9596_ (
    .A(_3044_),
    .B(_3040_),
    .Y(_3046_)
);

NAND2X1 _9597_ (
    .A(_3046_),
    .B(_3045_),
    .Y(_3047_)
);

OAI21X1 _9598_ (
    .A(_3037_),
    .B(_3038_),
    .C(_3047_),
    .Y(_3048_)
);

INVX1 _9599_ (
    .A(_3047_),
    .Y(_3049_)
);

NAND3X1 _9600_ (
    .A(_3027_),
    .B(_3049_),
    .C(_3029_),
    .Y(_3050_)
);

NAND3X1 _9601_ (
    .A(_2760_),
    .B(_3050_),
    .C(_3048_),
    .Y(_3051_)
);

AOI22X1 _9602_ (
    .A(_2723_),
    .B(_2756__bF$buf1),
    .C(_3051_),
    .D(_2880_),
    .Y(_2609_)
);

INVX1 _9603_ (
    .A(\genblk1[3].u_ce.Ycalc [0]),
    .Y(_3052_)
);

OAI21X1 _9604_ (
    .A(1'h0),
    .B(_2971_),
    .C(\genblk1[3].u_ce.Vld_bF$buf4 ),
    .Y(_3053_)
);

INVX2 _9605_ (
    .A(_3053_),
    .Y(_3054_)
);

INVX1 _9606_ (
    .A(\genblk1[3].u_ce.Yin0 [0]),
    .Y(_3055_)
);

AOI21X1 _9607_ (
    .A(_2822_),
    .B(_2829_),
    .C(_3055_),
    .Y(_3056_)
);

OAI21X1 _9608_ (
    .A(_3056_),
    .B(_2782_),
    .C(_3054_),
    .Y(_3057_)
);

OAI21X1 _9609_ (
    .A(_3052_),
    .B(\genblk1[3].u_ce.Vld_bF$buf3 ),
    .C(_3057_),
    .Y(_2610_)
);

NAND2X1 _9610_ (
    .A(\genblk1[3].u_ce.Ycalc [1]),
    .B(_2756__bF$buf0),
    .Y(_3058_)
);

NAND3X1 _9611_ (
    .A(_2844_),
    .B(_2781_),
    .C(_2845_),
    .Y(_3059_)
);

OAI21X1 _9612_ (
    .A(_2843_),
    .B(_2783_),
    .C(_2782_),
    .Y(_3060_)
);

AOI21X1 _9613_ (
    .A(_3060_),
    .B(_3059_),
    .C(_2761_),
    .Y(_3061_)
);

OAI21X1 _9614_ (
    .A(_2756__bF$buf4),
    .B(_3061_),
    .C(_3058_),
    .Y(_2611_)
);

NAND2X1 _9615_ (
    .A(\genblk1[3].u_ce.Xcalc [0]),
    .B(_2756__bF$buf3),
    .Y(_3062_)
);

MUX2X1 _9616_ (
    .A(\genblk1[3].u_ce.Yin12b [7]),
    .B(\genblk1[3].u_ce.Yin12b [6]),
    .S(1'h1),
    .Y(_3063_)
);

NAND2X1 _9617_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin12b [5]),
    .Y(_3064_)
);

OAI21X1 _9618_ (
    .A(1'h1),
    .B(_2883_),
    .C(_3064_),
    .Y(_3065_)
);

NAND2X1 _9619_ (
    .A(_2762__bF$buf4),
    .B(_3065_),
    .Y(_3066_)
);

OAI21X1 _9620_ (
    .A(_2762__bF$buf3),
    .B(_3063_),
    .C(_3066_),
    .Y(_3067_)
);

NAND2X1 _9621_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin1 [1]),
    .Y(_3068_)
);

OAI21X1 _9622_ (
    .A(1'h1),
    .B(_2785_),
    .C(_3068_),
    .Y(_3069_)
);

NAND2X1 _9623_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin0 [1]),
    .Y(_3070_)
);

OAI21X1 _9624_ (
    .A(1'h1),
    .B(_3055_),
    .C(_3070_),
    .Y(_3071_)
);

MUX2X1 _9625_ (
    .A(_3071_),
    .B(_3069_),
    .S(_2762__bF$buf2),
    .Y(_3072_)
);

NAND2X1 _9626_ (
    .A(_2789__bF$buf2),
    .B(_3072_),
    .Y(_3073_)
);

OAI21X1 _9627_ (
    .A(_2789__bF$buf1),
    .B(_3067_),
    .C(_3073_),
    .Y(_3074_)
);

INVX1 _9628_ (
    .A(_3074_),
    .Y(_3075_)
);

NOR2X1 _9629_ (
    .A(\genblk1[3].u_ce.Xin0 [0]),
    .B(_3075_),
    .Y(_3076_)
);

OAI21X1 _9630_ (
    .A(_2818_),
    .B(_3074_),
    .C(_3054_),
    .Y(_3077_)
);

OAI21X1 _9631_ (
    .A(_3077_),
    .B(_3076_),
    .C(_3062_),
    .Y(_2612_)
);

NAND2X1 _9632_ (
    .A(\genblk1[3].u_ce.Xcalc [1]),
    .B(_2756__bF$buf2),
    .Y(_3078_)
);

NOR2X1 _9633_ (
    .A(_2818_),
    .B(_3074_),
    .Y(_3079_)
);

NAND2X1 _9634_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin12b [4]),
    .Y(_3080_)
);

OAI21X1 _9635_ (
    .A(1'h1),
    .B(_2873_),
    .C(_3080_),
    .Y(_3081_)
);

NAND2X1 _9636_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin1 [0]),
    .Y(_3082_)
);

OAI21X1 _9637_ (
    .A(1'h1),
    .B(_2840_),
    .C(_3082_),
    .Y(_3083_)
);

MUX2X1 _9638_ (
    .A(_3083_),
    .B(_3081_),
    .S(_2762__bF$buf1),
    .Y(_3084_)
);

NAND2X1 _9639_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin12b [8]),
    .Y(_3085_)
);

OAI21X1 _9640_ (
    .A(1'h1),
    .B(_2957_),
    .C(_3085_),
    .Y(_3086_)
);

NAND2X1 _9641_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin12b [6]),
    .Y(_3087_)
);

OAI21X1 _9642_ (
    .A(1'h1),
    .B(_2908_),
    .C(_3087_),
    .Y(_3088_)
);

MUX2X1 _9643_ (
    .A(_3088_),
    .B(_3086_),
    .S(_2762__bF$buf0),
    .Y(_3089_)
);

MUX2X1 _9644_ (
    .A(_3089_),
    .B(_3084_),
    .S(1'h0),
    .Y(_3090_)
);

NOR2X1 _9645_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3074_),
    .Y(_3091_)
);

NAND2X1 _9646_ (
    .A(_3090_),
    .B(_3091_),
    .Y(_3092_)
);

NAND2X1 _9647_ (
    .A(_2789__bF$buf0),
    .B(_3084_),
    .Y(_3093_)
);

NAND2X1 _9648_ (
    .A(1'h0),
    .B(_3089_),
    .Y(_3094_)
);

NAND2X1 _9649_ (
    .A(_3093_),
    .B(_3094_),
    .Y(_3095_)
);

OAI21X1 _9650_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3074_),
    .C(_3095_),
    .Y(_3096_)
);

NAND3X1 _9651_ (
    .A(\genblk1[3].u_ce.Xin0 [1]),
    .B(_3096_),
    .C(_3092_),
    .Y(_3097_)
);

OAI21X1 _9652_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .B(_3074_),
    .C(_3090_),
    .Y(_3098_)
);

NAND2X1 _9653_ (
    .A(_3095_),
    .B(_3091_),
    .Y(_3099_)
);

NAND3X1 _9654_ (
    .A(_2798_),
    .B(_3098_),
    .C(_3099_),
    .Y(_3100_)
);

NAND3X1 _9655_ (
    .A(_3079_),
    .B(_3097_),
    .C(_3100_),
    .Y(_3101_)
);

INVX1 _9656_ (
    .A(_3079_),
    .Y(_3102_)
);

AOI21X1 _9657_ (
    .A(_3099_),
    .B(_3098_),
    .C(_2798_),
    .Y(_3103_)
);

AOI21X1 _9658_ (
    .A(_3092_),
    .B(_3096_),
    .C(\genblk1[3].u_ce.Xin0 [1]),
    .Y(_3104_)
);

OAI21X1 _9659_ (
    .A(_3103_),
    .B(_3104_),
    .C(_3102_),
    .Y(_3105_)
);

AOI21X1 _9660_ (
    .A(_3105_),
    .B(_3101_),
    .C(_2761_),
    .Y(_3106_)
);

OAI21X1 _9661_ (
    .A(_2756__bF$buf1),
    .B(_3106_),
    .C(_3078_),
    .Y(_2613_)
);

OAI21X1 _9662_ (
    .A(_3102_),
    .B(_3104_),
    .C(_3097_),
    .Y(_3107_)
);

MUX2X1 _9663_ (
    .A(\genblk1[3].u_ce.Yin12b [9]),
    .B(\genblk1[3].u_ce.Yin12b [8]),
    .S(1'h1),
    .Y(_3108_)
);

MUX2X1 _9664_ (
    .A(_3108_),
    .B(_3063_),
    .S(1'h1),
    .Y(_3109_)
);

NOR2X1 _9665_ (
    .A(1'h0),
    .B(_2762__bF$buf4),
    .Y(_3110_)
);

NAND2X1 _9666_ (
    .A(_3065_),
    .B(_3110_),
    .Y(_3111_)
);

NAND2X1 _9667_ (
    .A(_2759_),
    .B(_3069_),
    .Y(_3112_)
);

NAND2X1 _9668_ (
    .A(_3112_),
    .B(_3111_),
    .Y(_3113_)
);

AOI21X1 _9669_ (
    .A(1'h0),
    .B(_3109_),
    .C(_3113_),
    .Y(_3114_)
);

NAND2X1 _9670_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin12b [7]),
    .Y(_3115_)
);

OAI21X1 _9671_ (
    .A(1'h1),
    .B(_2932_),
    .C(_3115_),
    .Y(_3116_)
);

MUX2X1 _9672_ (
    .A(_3065_),
    .B(_3116_),
    .S(_2762__bF$buf3),
    .Y(_3117_)
);

NAND2X1 _9673_ (
    .A(1'h0),
    .B(_3117_),
    .Y(_3118_)
);

AOI21X1 _9674_ (
    .A(_3073_),
    .B(_3118_),
    .C(_3090_),
    .Y(_3119_)
);

NOR2X1 _9675_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .B(_3119_),
    .Y(_3120_)
);

NAND2X1 _9676_ (
    .A(_3114_),
    .B(_3120_),
    .Y(_3121_)
);

INVX1 _9677_ (
    .A(_3114_),
    .Y(_3122_)
);

OAI21X1 _9678_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf4 ),
    .B(_3119_),
    .C(_3122_),
    .Y(_3123_)
);

AOI21X1 _9679_ (
    .A(_3121_),
    .B(_3123_),
    .C(_2814_),
    .Y(_3124_)
);

NAND3X1 _9680_ (
    .A(_2814_),
    .B(_3123_),
    .C(_3121_),
    .Y(_3125_)
);

INVX1 _9681_ (
    .A(_3125_),
    .Y(_3126_)
);

NOR2X1 _9682_ (
    .A(_3124_),
    .B(_3126_),
    .Y(_3127_)
);

NOR2X1 _9683_ (
    .A(_3107_),
    .B(_3127_),
    .Y(_3128_)
);

AOI21X1 _9684_ (
    .A(_3079_),
    .B(_3100_),
    .C(_3103_),
    .Y(_3129_)
);

INVX1 _9685_ (
    .A(_3127_),
    .Y(_3130_)
);

OAI21X1 _9686_ (
    .A(_3129_),
    .B(_3130_),
    .C(_3054_),
    .Y(_3131_)
);

OAI22X1 _9687_ (
    .A(_2731_),
    .B(\genblk1[3].u_ce.Vld_bF$buf2 ),
    .C(_3128_),
    .D(_3131_),
    .Y(_2614_)
);

NAND2X1 _9688_ (
    .A(\genblk1[3].u_ce.Xcalc [3]),
    .B(_2756__bF$buf0),
    .Y(_3132_)
);

AOI21X1 _9689_ (
    .A(_3107_),
    .B(_3125_),
    .C(_3124_),
    .Y(_3133_)
);

NAND2X1 _9690_ (
    .A(1'h1),
    .B(_3018_),
    .Y(_3134_)
);

OAI21X1 _9691_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin12b [9]),
    .C(_3134_),
    .Y(_3135_)
);

NAND2X1 _9692_ (
    .A(_2762__bF$buf2),
    .B(_3086_),
    .Y(_3136_)
);

OAI21X1 _9693_ (
    .A(_2762__bF$buf1),
    .B(_3135_),
    .C(_3136_),
    .Y(_3137_)
);

NAND2X1 _9694_ (
    .A(_3088_),
    .B(_3110_),
    .Y(_3138_)
);

NAND2X1 _9695_ (
    .A(_2759_),
    .B(_3081_),
    .Y(_3139_)
);

NAND2X1 _9696_ (
    .A(_3139_),
    .B(_3138_),
    .Y(_3140_)
);

AOI21X1 _9697_ (
    .A(_3137_),
    .B(1'h0),
    .C(_3140_),
    .Y(_3141_)
);

NAND3X1 _9698_ (
    .A(_3114_),
    .B(_3095_),
    .C(_3074_),
    .Y(_3142_)
);

NAND2X1 _9699_ (
    .A(_2851__bF$buf2),
    .B(_3142_),
    .Y(_3143_)
);

OR2X2 _9700_ (
    .A(_3143_),
    .B(_3141_),
    .Y(_3144_)
);

INVX1 _9701_ (
    .A(_3142_),
    .Y(_3145_)
);

OAI21X1 _9702_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3145_),
    .C(_3141_),
    .Y(_3146_)
);

NAND3X1 _9703_ (
    .A(\genblk1[3].u_ce.Xin1 [1]),
    .B(_3146_),
    .C(_3144_),
    .Y(_3147_)
);

INVX1 _9704_ (
    .A(_3141_),
    .Y(_3148_)
);

OR2X2 _9705_ (
    .A(_3143_),
    .B(_3148_),
    .Y(_3149_)
);

OAI21X1 _9706_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3145_),
    .C(_3148_),
    .Y(_3150_)
);

NAND3X1 _9707_ (
    .A(_2793_),
    .B(_3150_),
    .C(_3149_),
    .Y(_3151_)
);

NAND2X1 _9708_ (
    .A(_3147_),
    .B(_3151_),
    .Y(_3152_)
);

OR2X2 _9709_ (
    .A(_3133_),
    .B(_3152_),
    .Y(_3153_)
);

NAND2X1 _9710_ (
    .A(_3152_),
    .B(_3133_),
    .Y(_3154_)
);

AOI21X1 _9711_ (
    .A(_3153_),
    .B(_3154_),
    .C(_2761_),
    .Y(_3155_)
);

OAI21X1 _9712_ (
    .A(_2756__bF$buf4),
    .B(_3155_),
    .C(_3132_),
    .Y(_2615_)
);

OAI21X1 _9713_ (
    .A(_3152_),
    .B(_3133_),
    .C(_3147_),
    .Y(_3156_)
);

NAND2X1 _9714_ (
    .A(1'h1),
    .B(\genblk1[3].u_ce.Yin12b [11]),
    .Y(_3157_)
);

OAI21X1 _9715_ (
    .A(1'h1),
    .B(_3018_),
    .C(_3157_),
    .Y(_3158_)
);

NAND2X1 _9716_ (
    .A(1'h1),
    .B(_3158_),
    .Y(_3159_)
);

OAI21X1 _9717_ (
    .A(1'h1),
    .B(_3108_),
    .C(_3159_),
    .Y(_3160_)
);

NAND2X1 _9718_ (
    .A(1'h0),
    .B(_3160_),
    .Y(_3161_)
);

OAI21X1 _9719_ (
    .A(1'h0),
    .B(_3117_),
    .C(_3161_),
    .Y(_3162_)
);

INVX1 _9720_ (
    .A(_3162_),
    .Y(_3163_)
);

OAI21X1 _9721_ (
    .A(_3148_),
    .B(_3142_),
    .C(_2851__bF$buf1),
    .Y(_3164_)
);

OR2X2 _9722_ (
    .A(_3164_),
    .B(_3163_),
    .Y(_3165_)
);

NAND2X1 _9723_ (
    .A(_3163_),
    .B(_3164_),
    .Y(_3166_)
);

NAND3X1 _9724_ (
    .A(\genblk1[3].u_ce.Xin12b [4]),
    .B(_3166_),
    .C(_3165_),
    .Y(_3167_)
);

OR2X2 _9725_ (
    .A(_3164_),
    .B(_3162_),
    .Y(_3168_)
);

NAND2X1 _9726_ (
    .A(_3162_),
    .B(_3164_),
    .Y(_3169_)
);

NAND3X1 _9727_ (
    .A(_2795_),
    .B(_3169_),
    .C(_3168_),
    .Y(_3170_)
);

AND2X2 _9728_ (
    .A(_3167_),
    .B(_3170_),
    .Y(_3171_)
);

NAND2X1 _9729_ (
    .A(_3171_),
    .B(_3156_),
    .Y(_3172_)
);

INVX1 _9730_ (
    .A(_3124_),
    .Y(_3173_)
);

OAI21X1 _9731_ (
    .A(_3126_),
    .B(_3129_),
    .C(_3173_),
    .Y(_3174_)
);

INVX1 _9732_ (
    .A(_3147_),
    .Y(_3175_)
);

AOI21X1 _9733_ (
    .A(_3174_),
    .B(_3151_),
    .C(_3175_),
    .Y(_3176_)
);

NAND2X1 _9734_ (
    .A(_3170_),
    .B(_3167_),
    .Y(_3177_)
);

NAND2X1 _9735_ (
    .A(_3177_),
    .B(_3176_),
    .Y(_3178_)
);

NAND2X1 _9736_ (
    .A(_3172_),
    .B(_3178_),
    .Y(_3179_)
);

AOI22X1 _9737_ (
    .A(_2733_),
    .B(_2756__bF$buf3),
    .C(_3179_),
    .D(_3054_),
    .Y(_2616_)
);

NAND3X1 _9738_ (
    .A(_3141_),
    .B(_3163_),
    .C(_3145_),
    .Y(_3180_)
);

NOR2X1 _9739_ (
    .A(1'h1),
    .B(_3135_),
    .Y(_3181_)
);

NOR2X1 _9740_ (
    .A(_2762__bF$buf0),
    .B(_3042_),
    .Y(_3182_)
);

OAI21X1 _9741_ (
    .A(_3182_),
    .B(_3181_),
    .C(1'h0),
    .Y(_3183_)
);

OAI21X1 _9742_ (
    .A(1'h0),
    .B(_3089_),
    .C(_3183_),
    .Y(_3184_)
);

NAND3X1 _9743_ (
    .A(_2851__bF$buf0),
    .B(_3184_),
    .C(_3180_),
    .Y(_3185_)
);

INVX1 _9744_ (
    .A(_3184_),
    .Y(_3186_)
);

NAND3X1 _9745_ (
    .A(_3114_),
    .B(_3141_),
    .C(_3119_),
    .Y(_3187_)
);

OAI21X1 _9746_ (
    .A(_3162_),
    .B(_3187_),
    .C(_2851__bF$buf5),
    .Y(_3188_)
);

NAND2X1 _9747_ (
    .A(_3186_),
    .B(_3188_),
    .Y(_3189_)
);

NAND3X1 _9748_ (
    .A(\genblk1[3].u_ce.Xin12b [5]),
    .B(_3189_),
    .C(_3185_),
    .Y(_3190_)
);

NAND3X1 _9749_ (
    .A(_2851__bF$buf4),
    .B(_3186_),
    .C(_3180_),
    .Y(_3191_)
);

NAND2X1 _9750_ (
    .A(_3184_),
    .B(_3188_),
    .Y(_3192_)
);

NAND3X1 _9751_ (
    .A(_2803_),
    .B(_3192_),
    .C(_3191_),
    .Y(_3193_)
);

NAND2X1 _9752_ (
    .A(_3190_),
    .B(_3193_),
    .Y(_3194_)
);

AOI21X1 _9753_ (
    .A(_3172_),
    .B(_3167_),
    .C(_3194_),
    .Y(_3195_)
);

OAI21X1 _9754_ (
    .A(_3177_),
    .B(_3176_),
    .C(_3167_),
    .Y(_3196_)
);

AND2X2 _9755_ (
    .A(_3190_),
    .B(_3193_),
    .Y(_3197_)
);

OAI21X1 _9756_ (
    .A(_3197_),
    .B(_3196_),
    .C(_3054_),
    .Y(_3198_)
);

OAI22X1 _9757_ (
    .A(_2748_),
    .B(\genblk1[3].u_ce.Vld_bF$buf1 ),
    .C(_3195_),
    .D(_3198_),
    .Y(_2617_)
);

NOR2X1 _9758_ (
    .A(_3162_),
    .B(_3187_),
    .Y(_3199_)
);

NAND2X1 _9759_ (
    .A(_3186_),
    .B(_3199_),
    .Y(_3200_)
);

AOI21X1 _9760_ (
    .A(_2762__bF$buf4),
    .B(_3158_),
    .C(_3182_),
    .Y(_3201_)
);

NAND2X1 _9761_ (
    .A(_2789__bF$buf3),
    .B(_3109_),
    .Y(_3202_)
);

OAI21X1 _9762_ (
    .A(_2789__bF$buf2),
    .B(_3201_),
    .C(_3202_),
    .Y(_3203_)
);

NAND3X1 _9763_ (
    .A(_2851__bF$buf3),
    .B(_3203_),
    .C(_3200_),
    .Y(_3204_)
);

NOR3X1 _9764_ (
    .A(_3162_),
    .B(_3184_),
    .C(_3187_),
    .Y(_3205_)
);

INVX1 _9765_ (
    .A(_3203_),
    .Y(_3206_)
);

OAI21X1 _9766_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .B(_3205_),
    .C(_3206_),
    .Y(_3207_)
);

NAND3X1 _9767_ (
    .A(\genblk1[3].u_ce.Xin12b [6]),
    .B(_3207_),
    .C(_3204_),
    .Y(_3208_)
);

NAND3X1 _9768_ (
    .A(_2851__bF$buf2),
    .B(_3206_),
    .C(_3200_),
    .Y(_3209_)
);

OAI21X1 _9769_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .B(_3205_),
    .C(_3203_),
    .Y(_3210_)
);

NAND3X1 _9770_ (
    .A(_2805_),
    .B(_3210_),
    .C(_3209_),
    .Y(_3211_)
);

AND2X2 _9771_ (
    .A(_3208_),
    .B(_3211_),
    .Y(_3212_)
);

NAND2X1 _9772_ (
    .A(_3171_),
    .B(_3197_),
    .Y(_3213_)
);

INVX1 _9773_ (
    .A(_3167_),
    .Y(_3214_)
);

INVX1 _9774_ (
    .A(_3190_),
    .Y(_3215_)
);

AOI21X1 _9775_ (
    .A(_3214_),
    .B(_3193_),
    .C(_3215_),
    .Y(_3216_)
);

OAI21X1 _9776_ (
    .A(_3176_),
    .B(_3213_),
    .C(_3216_),
    .Y(_3217_)
);

AND2X2 _9777_ (
    .A(_3217_),
    .B(_3212_),
    .Y(_3218_)
);

NOR2X1 _9778_ (
    .A(_3212_),
    .B(_3217_),
    .Y(_3219_)
);

OAI21X1 _9779_ (
    .A(_3219_),
    .B(_3218_),
    .C(_2760_),
    .Y(_3220_)
);

NAND2X1 _9780_ (
    .A(\genblk1[3].u_ce.Vld_bF$buf0 ),
    .B(_3220_),
    .Y(_3221_)
);

OAI21X1 _9781_ (
    .A(_2734_),
    .B(\genblk1[3].u_ce.Vld_bF$buf4 ),
    .C(_3221_),
    .Y(_2618_)
);

INVX1 _9782_ (
    .A(_3208_),
    .Y(_3222_)
);

NOR2X1 _9783_ (
    .A(_3222_),
    .B(_3218_),
    .Y(_3223_)
);

NAND2X1 _9784_ (
    .A(_3206_),
    .B(_3205_),
    .Y(_3224_)
);

NOR2X1 _9785_ (
    .A(_2789__bF$buf1),
    .B(_3042_),
    .Y(_3225_)
);

AOI21X1 _9786_ (
    .A(_3137_),
    .B(_2789__bF$buf0),
    .C(_3225_),
    .Y(_3226_)
);

NAND3X1 _9787_ (
    .A(_2851__bF$buf1),
    .B(_3226_),
    .C(_3224_),
    .Y(_3227_)
);

INVX1 _9788_ (
    .A(_3227_),
    .Y(_3228_)
);

AOI21X1 _9789_ (
    .A(_3224_),
    .B(_2851__bF$buf0),
    .C(_3226_),
    .Y(_3229_)
);

OAI21X1 _9790_ (
    .A(_3229_),
    .B(_3228_),
    .C(\genblk1[3].u_ce.Xin12b [7]),
    .Y(_3230_)
);

INVX1 _9791_ (
    .A(_3229_),
    .Y(_3231_)
);

NAND3X1 _9792_ (
    .A(_2808_),
    .B(_3227_),
    .C(_3231_),
    .Y(_3232_)
);

AND2X2 _9793_ (
    .A(_3232_),
    .B(_3230_),
    .Y(_3233_)
);

OR2X2 _9794_ (
    .A(_3223_),
    .B(_3233_),
    .Y(_3234_)
);

AOI21X1 _9795_ (
    .A(_3223_),
    .B(_3233_),
    .C(_3053_),
    .Y(_3235_)
);

AOI22X1 _9796_ (
    .A(_2747_),
    .B(_2756__bF$buf2),
    .C(_3234_),
    .D(_3235_),
    .Y(_2619_)
);

NOR2X1 _9797_ (
    .A(_3177_),
    .B(_3194_),
    .Y(_3236_)
);

OAI21X1 _9798_ (
    .A(_3167_),
    .B(_3194_),
    .C(_3190_),
    .Y(_3237_)
);

AOI21X1 _9799_ (
    .A(_3236_),
    .B(_3156_),
    .C(_3237_),
    .Y(_3238_)
);

AOI21X1 _9800_ (
    .A(_3231_),
    .B(_3227_),
    .C(_2808_),
    .Y(_3239_)
);

AOI21X1 _9801_ (
    .A(_3222_),
    .B(_3232_),
    .C(_3239_),
    .Y(_3240_)
);

NAND3X1 _9802_ (
    .A(_3212_),
    .B(_3230_),
    .C(_3232_),
    .Y(_3241_)
);

OAI21X1 _9803_ (
    .A(_3241_),
    .B(_3238_),
    .C(_3240_),
    .Y(_3242_)
);

NAND3X1 _9804_ (
    .A(_3206_),
    .B(_3226_),
    .C(_3205_),
    .Y(_3243_)
);

INVX1 _9805_ (
    .A(_3160_),
    .Y(_3244_)
);

INVX1 _9806_ (
    .A(_3225_),
    .Y(_3245_)
);

OAI21X1 _9807_ (
    .A(1'h0),
    .B(_3244_),
    .C(_3245_),
    .Y(_3246_)
);

INVX1 _9808_ (
    .A(_3246_),
    .Y(_3247_)
);

NAND3X1 _9809_ (
    .A(_2851__bF$buf5),
    .B(_3247_),
    .C(_3243_),
    .Y(_3248_)
);

INVX1 _9810_ (
    .A(_3248_),
    .Y(_3249_)
);

AOI21X1 _9811_ (
    .A(_3243_),
    .B(_2851__bF$buf4),
    .C(_3247_),
    .Y(_3250_)
);

OAI21X1 _9812_ (
    .A(_3250_),
    .B(_3249_),
    .C(\genblk1[3].u_ce.Xin12b [8]),
    .Y(_3251_)
);

INVX1 _9813_ (
    .A(_3250_),
    .Y(_3252_)
);

NAND3X1 _9814_ (
    .A(_2810_),
    .B(_3248_),
    .C(_3252_),
    .Y(_3253_)
);

AND2X2 _9815_ (
    .A(_3253_),
    .B(_3251_),
    .Y(_3254_)
);

OR2X2 _9816_ (
    .A(_3242_),
    .B(_3254_),
    .Y(_3255_)
);

INVX1 _9817_ (
    .A(_3255_),
    .Y(_3256_)
);

NAND2X1 _9818_ (
    .A(_3254_),
    .B(_3242_),
    .Y(_3257_)
);

NAND2X1 _9819_ (
    .A(_3054_),
    .B(_3257_),
    .Y(_3258_)
);

OAI22X1 _9820_ (
    .A(_2736_),
    .B(\genblk1[3].u_ce.Vld_bF$buf3 ),
    .C(_3258_),
    .D(_3256_),
    .Y(_2620_)
);

NOR3X1 _9821_ (
    .A(_3184_),
    .B(_3203_),
    .C(_3180_),
    .Y(_3259_)
);

NAND3X1 _9822_ (
    .A(_3226_),
    .B(_3247_),
    .C(_3259_),
    .Y(_3260_)
);

OR2X2 _9823_ (
    .A(_3181_),
    .B(_3182_),
    .Y(_3261_)
);

AOI21X1 _9824_ (
    .A(_3261_),
    .B(_2789__bF$buf3),
    .C(_3225_),
    .Y(_3262_)
);

INVX1 _9825_ (
    .A(_3262_),
    .Y(_3263_)
);

NAND3X1 _9826_ (
    .A(_2851__bF$buf3),
    .B(_3263_),
    .C(_3260_),
    .Y(_3264_)
);

OAI21X1 _9827_ (
    .A(_3246_),
    .B(_3243_),
    .C(_2851__bF$buf2),
    .Y(_3265_)
);

NAND2X1 _9828_ (
    .A(_3262_),
    .B(_3265_),
    .Y(_3266_)
);

NAND3X1 _9829_ (
    .A(\genblk1[3].u_ce.Xin12b [9]),
    .B(_3266_),
    .C(_3264_),
    .Y(_3267_)
);

NAND3X1 _9830_ (
    .A(_2851__bF$buf1),
    .B(_3262_),
    .C(_3260_),
    .Y(_3268_)
);

NAND2X1 _9831_ (
    .A(_3263_),
    .B(_3265_),
    .Y(_3269_)
);

NAND3X1 _9832_ (
    .A(_2855_),
    .B(_3269_),
    .C(_3268_),
    .Y(_3270_)
);

NAND2X1 _9833_ (
    .A(_3267_),
    .B(_3270_),
    .Y(_3271_)
);

AOI21X1 _9834_ (
    .A(_3257_),
    .B(_3251_),
    .C(_3271_),
    .Y(_3272_)
);

NAND3X1 _9835_ (
    .A(_3251_),
    .B(_3271_),
    .C(_3257_),
    .Y(_3273_)
);

NAND2X1 _9836_ (
    .A(_3054_),
    .B(_3273_),
    .Y(_3274_)
);

OAI22X1 _9837_ (
    .A(_2744_),
    .B(\genblk1[3].u_ce.Vld_bF$buf2 ),
    .C(_3272_),
    .D(_3274_),
    .Y(_2621_)
);

NAND2X1 _9838_ (
    .A(\genblk1[3].u_ce.Xcalc [10]),
    .B(_2756__bF$buf1),
    .Y(_3275_)
);

OAI21X1 _9839_ (
    .A(1'h0),
    .B(_3201_),
    .C(_3245_),
    .Y(_3276_)
);

OAI21X1 _9840_ (
    .A(_3263_),
    .B(_3260_),
    .C(_2851__bF$buf0),
    .Y(_3277_)
);

NOR2X1 _9841_ (
    .A(_3276_),
    .B(_3277_),
    .Y(_3278_)
);

NAND2X1 _9842_ (
    .A(_3276_),
    .B(_3277_),
    .Y(_3279_)
);

INVX1 _9843_ (
    .A(_3279_),
    .Y(_3280_)
);

OAI21X1 _9844_ (
    .A(_3278_),
    .B(_3280_),
    .C(\genblk1[3].u_ce.Xin12b [10]),
    .Y(_3281_)
);

INVX1 _9845_ (
    .A(_3278_),
    .Y(_3282_)
);

NAND3X1 _9846_ (
    .A(_2885_),
    .B(_3279_),
    .C(_3282_),
    .Y(_3283_)
);

AND2X2 _9847_ (
    .A(_3283_),
    .B(_3281_),
    .Y(_3284_)
);

OAI21X1 _9848_ (
    .A(_3251_),
    .B(_3271_),
    .C(_3267_),
    .Y(_3285_)
);

NAND3X1 _9849_ (
    .A(_3212_),
    .B(_3217_),
    .C(_3233_),
    .Y(_3286_)
);

NAND3X1 _9850_ (
    .A(_3267_),
    .B(_3270_),
    .C(_3254_),
    .Y(_3287_)
);

AOI21X1 _9851_ (
    .A(_3286_),
    .B(_3240_),
    .C(_3287_),
    .Y(_3288_)
);

OAI21X1 _9852_ (
    .A(_3285_),
    .B(_3288_),
    .C(_3284_),
    .Y(_3289_)
);

NAND2X1 _9853_ (
    .A(_3281_),
    .B(_3283_),
    .Y(_3290_)
);

NAND2X1 _9854_ (
    .A(_3251_),
    .B(_3253_),
    .Y(_3291_)
);

NOR2X1 _9855_ (
    .A(_3291_),
    .B(_3271_),
    .Y(_3292_)
);

AOI21X1 _9856_ (
    .A(_3242_),
    .B(_3292_),
    .C(_3285_),
    .Y(_3293_)
);

NAND2X1 _9857_ (
    .A(_3290_),
    .B(_3293_),
    .Y(_3294_)
);

AOI21X1 _9858_ (
    .A(_3289_),
    .B(_3294_),
    .C(_2761_),
    .Y(_3295_)
);

OAI21X1 _9859_ (
    .A(_2756__bF$buf0),
    .B(_3295_),
    .C(_3275_),
    .Y(_2622_)
);

NAND2X1 _9860_ (
    .A(\genblk1[3].u_ce.Xcalc [11]),
    .B(_2756__bF$buf4),
    .Y(_3296_)
);

OR2X2 _9861_ (
    .A(_3260_),
    .B(_3263_),
    .Y(_3297_)
);

OAI21X1 _9862_ (
    .A(_3276_),
    .B(_3297_),
    .C(_2851__bF$buf5),
    .Y(_3298_)
);

OR2X2 _9863_ (
    .A(_3298_),
    .B(_3044_),
    .Y(_3299_)
);

NAND2X1 _9864_ (
    .A(_3044_),
    .B(_3298_),
    .Y(_3300_)
);

AOI22X1 _9865_ (
    .A(_3299_),
    .B(_3300_),
    .C(_3289_),
    .D(_3281_),
    .Y(_3301_)
);

OAI21X1 _9866_ (
    .A(_3290_),
    .B(_3293_),
    .C(_3281_),
    .Y(_3302_)
);

NAND2X1 _9867_ (
    .A(_3300_),
    .B(_3299_),
    .Y(_3303_)
);

OAI21X1 _9868_ (
    .A(_3303_),
    .B(_3302_),
    .C(_3054_),
    .Y(_3304_)
);

OAI21X1 _9869_ (
    .A(_3301_),
    .B(_3304_),
    .C(_3296_),
    .Y(_2623_)
);

NAND2X1 _9870_ (
    .A(1'h1),
    .B(1'h1),
    .Y(_3305_)
);

OAI21X1 _9871_ (
    .A(_2789__bF$buf2),
    .B(_2971_),
    .C(_3305_),
    .Y(_3306_)
);

NOR2X1 _9872_ (
    .A(_2752_),
    .B(_3306_),
    .Y(_3307_)
);

AND2X2 _9873_ (
    .A(_3306_),
    .B(_2752_),
    .Y(_3308_)
);

OR2X2 _9874_ (
    .A(_3308_),
    .B(_3307_),
    .Y(_3309_)
);

NAND2X1 _9875_ (
    .A(\genblk1[3].u_ce.Acalc [0]),
    .B(_2756__bF$buf3),
    .Y(_3310_)
);

OAI21X1 _9876_ (
    .A(_2756__bF$buf2),
    .B(_3309_),
    .C(_3310_),
    .Y(_2624_)
);

NAND2X1 _9877_ (
    .A(\genblk1[3].u_ce.Acalc [1]),
    .B(_2756__bF$buf1),
    .Y(_3311_)
);

OAI21X1 _9878_ (
    .A(1'h1),
    .B(_2758_),
    .C(1'h0),
    .Y(_3312_)
);

OAI21X1 _9879_ (
    .A(1'h0),
    .B(_2758_),
    .C(_3312_),
    .Y(_3313_)
);

OAI21X1 _9880_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf4 ),
    .B(_3306_),
    .C(_3313_),
    .Y(_3314_)
);

OAI21X1 _9881_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3313_),
    .C(_3314_),
    .Y(_3315_)
);

OR2X2 _9882_ (
    .A(_3315_),
    .B(\genblk1[3].u_ce.Ain0 [1]),
    .Y(_3316_)
);

NAND2X1 _9883_ (
    .A(\genblk1[3].u_ce.Ain0 [1]),
    .B(_3315_),
    .Y(_3317_)
);

NAND2X1 _9884_ (
    .A(_3317_),
    .B(_3316_),
    .Y(_3318_)
);

NOR2X1 _9885_ (
    .A(_3307_),
    .B(_3318_),
    .Y(_3319_)
);

NAND2X1 _9886_ (
    .A(_3307_),
    .B(_3318_),
    .Y(_3320_)
);

NAND2X1 _9887_ (
    .A(\genblk1[3].u_ce.Vld_bF$buf1 ),
    .B(_3320_),
    .Y(_3321_)
);

OAI21X1 _9888_ (
    .A(_3319_),
    .B(_3321_),
    .C(_3311_),
    .Y(_2625_)
);

NAND2X1 _9889_ (
    .A(\genblk1[3].u_ce.Acalc [2]),
    .B(_2756__bF$buf0),
    .Y(_3322_)
);

OAI21X1 _9890_ (
    .A(_2754_),
    .B(_3315_),
    .C(_3320_),
    .Y(_3323_)
);

OAI21X1 _9891_ (
    .A(_2758_),
    .B(_2762__bF$buf3),
    .C(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .Y(_3324_)
);

NAND3X1 _9892_ (
    .A(1'h0),
    .B(_2971_),
    .C(_3324_),
    .Y(_3325_)
);

OAI21X1 _9893_ (
    .A(1'h0),
    .B(_3324_),
    .C(_3325_),
    .Y(_3326_)
);

NAND2X1 _9894_ (
    .A(\genblk1[3].u_ce.Ain1 [0]),
    .B(_3326_),
    .Y(_3327_)
);

OR2X2 _9895_ (
    .A(_3326_),
    .B(\genblk1[3].u_ce.Ain1 [0]),
    .Y(_3328_)
);

NAND2X1 _9896_ (
    .A(_3327_),
    .B(_3328_),
    .Y(_3329_)
);

INVX1 _9897_ (
    .A(_3329_),
    .Y(_3330_)
);

NOR2X1 _9898_ (
    .A(_3330_),
    .B(_3323_),
    .Y(_3331_)
);

NAND2X1 _9899_ (
    .A(_3330_),
    .B(_3323_),
    .Y(_3332_)
);

NAND2X1 _9900_ (
    .A(\genblk1[3].u_ce.Vld_bF$buf0 ),
    .B(_3332_),
    .Y(_3333_)
);

OAI21X1 _9901_ (
    .A(_3331_),
    .B(_3333_),
    .C(_3322_),
    .Y(_2626_)
);

NAND2X1 _9902_ (
    .A(_3327_),
    .B(_3332_),
    .Y(_3334_)
);

INVX1 _9903_ (
    .A(_3334_),
    .Y(_3335_)
);

INVX1 _9904_ (
    .A(\genblk1[3].u_ce.Ain1 [1]),
    .Y(_3336_)
);

OAI21X1 _9905_ (
    .A(1'h1),
    .B(_2762__bF$buf2),
    .C(1'h0),
    .Y(_3337_)
);

NAND2X1 _9906_ (
    .A(_2851__bF$buf4),
    .B(_3337_),
    .Y(_3338_)
);

OAI21X1 _9907_ (
    .A(1'h0),
    .B(1'h1),
    .C(\genblk1[3].u_ce.Ain12b_11_bF$buf1 ),
    .Y(_3339_)
);

OAI21X1 _9908_ (
    .A(_2758_),
    .B(_3339_),
    .C(_3338_),
    .Y(_3340_)
);

NOR2X1 _9909_ (
    .A(_3336_),
    .B(_3340_),
    .Y(_3341_)
);

NAND2X1 _9910_ (
    .A(_3336_),
    .B(_3340_),
    .Y(_3342_)
);

INVX1 _9911_ (
    .A(_3342_),
    .Y(_3343_)
);

OAI21X1 _9912_ (
    .A(_3341_),
    .B(_3343_),
    .C(_3335_),
    .Y(_3344_)
);

INVX1 _9913_ (
    .A(_3341_),
    .Y(_3345_)
);

NAND3X1 _9914_ (
    .A(_3345_),
    .B(_3342_),
    .C(_3334_),
    .Y(_3346_)
);

NAND2X1 _9915_ (
    .A(_3346_),
    .B(_3344_),
    .Y(_3347_)
);

NAND2X1 _9916_ (
    .A(\genblk1[3].u_ce.Acalc [3]),
    .B(_2756__bF$buf4),
    .Y(_3348_)
);

OAI21X1 _9917_ (
    .A(_2756__bF$buf3),
    .B(_3347_),
    .C(_3348_),
    .Y(_2627_)
);

NOR2X1 _9918_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf0 ),
    .B(_3313_),
    .Y(_3349_)
);

NAND3X1 _9919_ (
    .A(1'h1),
    .B(_2789__bF$buf1),
    .C(_2762__bF$buf1),
    .Y(_3350_)
);

AOI21X1 _9920_ (
    .A(_3312_),
    .B(_3350_),
    .C(_2851__bF$buf3),
    .Y(_3351_)
);

NOR2X1 _9921_ (
    .A(_3351_),
    .B(_3349_),
    .Y(_3352_)
);

NAND2X1 _9922_ (
    .A(\genblk1[3].u_ce.Ain12b [4]),
    .B(_3352_),
    .Y(_3353_)
);

INVX1 _9923_ (
    .A(\genblk1[3].u_ce.Ain12b [4]),
    .Y(_3354_)
);

OAI21X1 _9924_ (
    .A(_3351_),
    .B(_3349_),
    .C(_3354_),
    .Y(_3355_)
);

NAND2X1 _9925_ (
    .A(_3355_),
    .B(_3353_),
    .Y(_3356_)
);

AOI21X1 _9926_ (
    .A(_3334_),
    .B(_3342_),
    .C(_3341_),
    .Y(_3357_)
);

AND2X2 _9927_ (
    .A(_3357_),
    .B(_3356_),
    .Y(_3358_)
);

OAI21X1 _9928_ (
    .A(_3356_),
    .B(_3357_),
    .C(\genblk1[3].u_ce.Vld_bF$buf4 ),
    .Y(_3359_)
);

OAI22X1 _9929_ (
    .A(_2695_),
    .B(\genblk1[3].u_ce.Vld_bF$buf3 ),
    .C(_3359_),
    .D(_3358_),
    .Y(_2628_)
);

NAND2X1 _9930_ (
    .A(\genblk1[3].u_ce.Acalc [5]),
    .B(_2756__bF$buf2),
    .Y(_3360_)
);

OAI21X1 _9931_ (
    .A(_3356_),
    .B(_3357_),
    .C(_3353_),
    .Y(_3361_)
);

OAI21X1 _9932_ (
    .A(1'h1),
    .B(1'h1),
    .C(_2790_),
    .Y(_3362_)
);

NAND2X1 _9933_ (
    .A(_2851__bF$buf2),
    .B(_3362_),
    .Y(_3363_)
);

INVX1 _9934_ (
    .A(_3363_),
    .Y(_3364_)
);

NOR2X1 _9935_ (
    .A(_2851__bF$buf1),
    .B(_3362_),
    .Y(_3365_)
);

NOR2X1 _9936_ (
    .A(_3365_),
    .B(_3364_),
    .Y(_3366_)
);

NAND2X1 _9937_ (
    .A(\genblk1[3].u_ce.Ain12b [5]),
    .B(_3366_),
    .Y(_3367_)
);

INVX1 _9938_ (
    .A(\genblk1[3].u_ce.Ain12b [5]),
    .Y(_3368_)
);

OAI21X1 _9939_ (
    .A(_3365_),
    .B(_3364_),
    .C(_3368_),
    .Y(_3369_)
);

NAND2X1 _9940_ (
    .A(_3369_),
    .B(_3367_),
    .Y(_3370_)
);

INVX1 _9941_ (
    .A(_3370_),
    .Y(_3371_)
);

NOR2X1 _9942_ (
    .A(_3371_),
    .B(_3361_),
    .Y(_3372_)
);

NAND2X1 _9943_ (
    .A(_3371_),
    .B(_3361_),
    .Y(_3373_)
);

NAND2X1 _9944_ (
    .A(\genblk1[3].u_ce.Vld_bF$buf2 ),
    .B(_3373_),
    .Y(_3374_)
);

OAI21X1 _9945_ (
    .A(_3372_),
    .B(_3374_),
    .C(_3360_),
    .Y(_2629_)
);

NAND2X1 _9946_ (
    .A(\genblk1[3].u_ce.Acalc [6]),
    .B(_2756__bF$buf1),
    .Y(_3375_)
);

INVX1 _9947_ (
    .A(_3357_),
    .Y(_3376_)
);

NOR2X1 _9948_ (
    .A(_3356_),
    .B(_3370_),
    .Y(_3377_)
);

OAI21X1 _9949_ (
    .A(_3353_),
    .B(_3370_),
    .C(_3367_),
    .Y(_3378_)
);

AOI21X1 _9950_ (
    .A(_3376_),
    .B(_3377_),
    .C(_3378_),
    .Y(_3379_)
);

OAI21X1 _9951_ (
    .A(1'h0),
    .B(_3305_),
    .C(_2760_),
    .Y(_3380_)
);

NOR2X1 _9952_ (
    .A(_2851__bF$buf0),
    .B(_3380_),
    .Y(_3381_)
);

NAND2X1 _9953_ (
    .A(_2851__bF$buf5),
    .B(_3380_),
    .Y(_3382_)
);

INVX1 _9954_ (
    .A(_3382_),
    .Y(_3383_)
);

NOR2X1 _9955_ (
    .A(_3381_),
    .B(_3383_),
    .Y(_3384_)
);

NAND2X1 _9956_ (
    .A(\genblk1[3].u_ce.Ain12b [6]),
    .B(_3384_),
    .Y(_3385_)
);

OR2X2 _9957_ (
    .A(_3384_),
    .B(\genblk1[3].u_ce.Ain12b [6]),
    .Y(_3386_)
);

AND2X2 _9958_ (
    .A(_3386_),
    .B(_3385_),
    .Y(_3387_)
);

INVX1 _9959_ (
    .A(_3387_),
    .Y(_3388_)
);

AND2X2 _9960_ (
    .A(_3379_),
    .B(_3388_),
    .Y(_3389_)
);

OAI21X1 _9961_ (
    .A(_3388_),
    .B(_3379_),
    .C(\genblk1[3].u_ce.Vld_bF$buf1 ),
    .Y(_3390_)
);

OAI21X1 _9962_ (
    .A(_3390_),
    .B(_3389_),
    .C(_3375_),
    .Y(_2630_)
);

OAI21X1 _9963_ (
    .A(_3388_),
    .B(_3379_),
    .C(_3385_),
    .Y(_3391_)
);

OAI21X1 _9964_ (
    .A(1'h0),
    .B(1'h1),
    .C(\genblk1[3].u_ce.Ain12b_11_bF$buf4 ),
    .Y(_3392_)
);

NAND2X1 _9965_ (
    .A(_3392_),
    .B(_2852_),
    .Y(_3393_)
);

INVX1 _9966_ (
    .A(_3393_),
    .Y(_3394_)
);

NAND2X1 _9967_ (
    .A(\genblk1[3].u_ce.Ain12b [7]),
    .B(_3394_),
    .Y(_3395_)
);

INVX1 _9968_ (
    .A(_3395_),
    .Y(_3396_)
);

NOR2X1 _9969_ (
    .A(\genblk1[3].u_ce.Ain12b [7]),
    .B(_3394_),
    .Y(_3397_)
);

NOR2X1 _9970_ (
    .A(_3397_),
    .B(_3396_),
    .Y(_3398_)
);

INVX1 _9971_ (
    .A(_3398_),
    .Y(_3399_)
);

OR2X2 _9972_ (
    .A(_3391_),
    .B(_3399_),
    .Y(_3400_)
);

AOI21X1 _9973_ (
    .A(_3391_),
    .B(_3399_),
    .C(_2756__bF$buf0),
    .Y(_3401_)
);

AOI22X1 _9974_ (
    .A(_2709_),
    .B(_2756__bF$buf4),
    .C(_3400_),
    .D(_3401_),
    .Y(_2631_)
);

NAND2X1 _9975_ (
    .A(\genblk1[3].u_ce.Acalc [8]),
    .B(_2756__bF$buf3),
    .Y(_3402_)
);

OAI21X1 _9976_ (
    .A(_3397_),
    .B(_3385_),
    .C(_3395_),
    .Y(_3403_)
);

NAND2X1 _9977_ (
    .A(_3398_),
    .B(_3387_),
    .Y(_3404_)
);

INVX1 _9978_ (
    .A(_3404_),
    .Y(_3405_)
);

AOI21X1 _9979_ (
    .A(_3405_),
    .B(_3378_),
    .C(_3403_),
    .Y(_3406_)
);

NAND2X1 _9980_ (
    .A(_3377_),
    .B(_3405_),
    .Y(_3407_)
);

OAI21X1 _9981_ (
    .A(_3407_),
    .B(_3357_),
    .C(_3406_),
    .Y(_3408_)
);

INVX1 _9982_ (
    .A(\genblk1[3].u_ce.Ain12b [8]),
    .Y(_3409_)
);

NAND2X1 _9983_ (
    .A(_2851__bF$buf4),
    .B(_2759_),
    .Y(_3410_)
);

NAND2X1 _9984_ (
    .A(_3339_),
    .B(_3410_),
    .Y(_3411_)
);

OR2X2 _9985_ (
    .A(_3411_),
    .B(_3409_),
    .Y(_3412_)
);

NAND2X1 _9986_ (
    .A(_3409_),
    .B(_3411_),
    .Y(_3413_)
);

AND2X2 _9987_ (
    .A(_3412_),
    .B(_3413_),
    .Y(_3414_)
);

NOR2X1 _9988_ (
    .A(_3414_),
    .B(_3408_),
    .Y(_3415_)
);

NAND2X1 _9989_ (
    .A(_3414_),
    .B(_3408_),
    .Y(_3416_)
);

NAND2X1 _9990_ (
    .A(\genblk1[3].u_ce.Vld_bF$buf0 ),
    .B(_3416_),
    .Y(_3417_)
);

OAI21X1 _9991_ (
    .A(_3415_),
    .B(_3417_),
    .C(_3402_),
    .Y(_2632_)
);

NAND2X1 _9992_ (
    .A(\genblk1[3].u_ce.Acalc [9]),
    .B(_2756__bF$buf2),
    .Y(_3418_)
);

OAI21X1 _9993_ (
    .A(_3409_),
    .B(_3411_),
    .C(_3416_),
    .Y(_3419_)
);

INVX1 _9994_ (
    .A(\genblk1[3].u_ce.Ain12b [9]),
    .Y(_3420_)
);

NAND2X1 _9995_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf3 ),
    .B(_3420_),
    .Y(_3421_)
);

NOR2X1 _9996_ (
    .A(\genblk1[3].u_ce.Ain12b_11_bF$buf2 ),
    .B(_3420_),
    .Y(_3422_)
);

INVX1 _9997_ (
    .A(_3422_),
    .Y(_3423_)
);

NAND2X1 _9998_ (
    .A(_3421_),
    .B(_3423_),
    .Y(_3424_)
);

INVX1 _9999_ (
    .A(_3424_),
    .Y(_3425_)
);

endmodule
