magic
tech scmos
magscale 1 6
timestamp 1569533753
<< checkpaint >>
rect -140 -1950 2540 5180
<< metal2 >>
rect 2260 5032 2324 5060
use CMD_TR$1  CMD_TR$1_0
timestamp 1569533753
transform 1 0 1524 0 1 4798
box 10 -35 254 178
use DOUBLE_GUARD$1  DOUBLE_GUARD$1_0
timestamp 1569533753
transform 1 0 0 0 1 1660
box -20 -20 2419 500
use GUARD$1  GUARD$1_0
timestamp 1569533753
transform 1 0 0 0 1 4220
box -20 -20 2419 792
use INV$1  INV$1_0
timestamp 1569533753
transform 1 0 1738 0 1 4314
box -2 -42 186 614
use INV2$1  INV2$1_0
timestamp 1569533753
transform 1 0 1914 0 1 4314
box -2 -42 426 646
use METAL_RING$1  METAL_RING$1_0
timestamp 1569533753
transform 1 0 0 0 1 0
box 0 0 2400 5012
use NDRV$1  NDRV$1_0
timestamp 1569533753
transform 1 0 0 0 1 0
box 0 0 2400 1560
use PAD_80$1  PAD_80$1_0
timestamp 1569533753
transform 1 0 1200 0 1 -980
box -850 -850 850 980
use PAD_METAL_PIC$1  PAD_METAL_PIC$1_0
timestamp 1569533753
transform 1 0 0 0 1 0
box 0 0 2400 5060
use PDRV$1  PDRV$1_0
timestamp 1569533753
transform 1 0 0 0 1 2260
box -20 -20 2420 1580
use SINGLE_GUARD$1  SINGLE_GUARD$1_0
timestamp 1569533753
transform 1 0 0 0 1 3920
box 0 0 2400 200
<< labels >>
flabel m2p s 2292 5060 2292 5060 0 FreeSans 400 0 0 0 Y
flabel space 1200 -980 1200 -980 0 FreeSans 1000 0 0 0 PAD
flabel m3p s 0 3018 0 3018 0 FreeSans 1000 0 0 0 VDD
flabel m3p s 0 4339 0 4339 0 FreeSans 1000 0 0 0 VDD
flabel m3p s 0 4788 0 4788 0 FreeSans 1000 0 0 0 VSS
flabel m3p s 0 752 0 752 0 FreeSans 1000 0 0 0 VSS
<< end >>
